module FIR_Lowpass_Filter (clk,
    data_in,
    data_out);
 input clk;
 input [15:0] data_in;
 output [40:0] data_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire _19089_;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire _19096_;
 wire _19097_;
 wire _19098_;
 wire _19099_;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire _19106_;
 wire _19107_;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire _19112_;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire _19135_;
 wire _19136_;
 wire _19137_;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire _19141_;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire _19168_;
 wire _19169_;
 wire _19170_;
 wire _19171_;
 wire _19172_;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire _19179_;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire _19194_;
 wire _19195_;
 wire _19196_;
 wire _19197_;
 wire _19198_;
 wire _19199_;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire _19216_;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire _19228_;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire _19235_;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire _19241_;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire _19260_;
 wire _19261_;
 wire _19262_;
 wire _19263_;
 wire _19264_;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire _19268_;
 wire _19269_;
 wire _19270_;
 wire _19271_;
 wire _19272_;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire _19395_;
 wire _19396_;
 wire _19397_;
 wire _19398_;
 wire _19399_;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire _19407_;
 wire _19408_;
 wire _19409_;
 wire _19410_;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire _19424_;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire _19461_;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire _19472_;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire _19506_;
 wire _19507_;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire _19512_;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire _19519_;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire _19524_;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire _19530_;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire _19534_;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire _19545_;
 wire _19546_;
 wire _19547_;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire _19557_;
 wire _19558_;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire _19583_;
 wire _19584_;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire _19590_;
 wire _19591_;
 wire _19592_;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire _19605_;
 wire _19606_;
 wire _19607_;
 wire _19608_;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire _19624_;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire _19631_;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire _19635_;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire _19642_;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire _19648_;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire _19653_;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire _19671_;
 wire _19672_;
 wire _19673_;
 wire _19674_;
 wire _19675_;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire _19683_;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire _19692_;
 wire _19693_;
 wire _19694_;
 wire _19695_;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire _19719_;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire _19797_;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire _19839_;
 wire _19840_;
 wire _19841_;
 wire _19842_;
 wire _19843_;
 wire _19844_;
 wire _19845_;
 wire _19846_;
 wire _19847_;
 wire _19848_;
 wire _19849_;
 wire _19850_;
 wire _19851_;
 wire _19852_;
 wire _19853_;
 wire _19854_;
 wire _19855_;
 wire _19856_;
 wire _19857_;
 wire _19858_;
 wire _19859_;
 wire _19860_;
 wire _19861_;
 wire _19862_;
 wire _19863_;
 wire _19864_;
 wire _19865_;
 wire _19866_;
 wire _19867_;
 wire _19868_;
 wire _19869_;
 wire _19870_;
 wire _19871_;
 wire _19872_;
 wire _19873_;
 wire _19874_;
 wire _19875_;
 wire _19876_;
 wire _19877_;
 wire _19878_;
 wire _19879_;
 wire _19880_;
 wire _19881_;
 wire _19882_;
 wire _19883_;
 wire _19884_;
 wire _19885_;
 wire _19886_;
 wire _19887_;
 wire _19888_;
 wire _19889_;
 wire _19890_;
 wire _19891_;
 wire _19892_;
 wire _19893_;
 wire _19894_;
 wire _19895_;
 wire _19896_;
 wire _19897_;
 wire _19898_;
 wire _19899_;
 wire _19900_;
 wire _19901_;
 wire _19902_;
 wire _19903_;
 wire _19904_;
 wire _19905_;
 wire _19906_;
 wire _19907_;
 wire _19908_;
 wire _19909_;
 wire _19910_;
 wire _19911_;
 wire _19912_;
 wire _19913_;
 wire _19914_;
 wire _19915_;
 wire _19916_;
 wire _19917_;
 wire _19918_;
 wire _19919_;
 wire _19920_;
 wire _19921_;
 wire _19922_;
 wire _19923_;
 wire _19924_;
 wire _19925_;
 wire _19926_;
 wire _19927_;
 wire _19928_;
 wire _19929_;
 wire _19930_;
 wire _19931_;
 wire _19932_;
 wire _19933_;
 wire _19934_;
 wire _19935_;
 wire _19936_;
 wire _19937_;
 wire _19938_;
 wire _19939_;
 wire _19940_;
 wire _19941_;
 wire _19942_;
 wire _19943_;
 wire _19944_;
 wire _19945_;
 wire _19946_;
 wire _19947_;
 wire _19948_;
 wire _19949_;
 wire _19950_;
 wire _19951_;
 wire _19952_;
 wire _19953_;
 wire _19954_;
 wire _19955_;
 wire _19956_;
 wire _19957_;
 wire _19958_;
 wire _19959_;
 wire _19960_;
 wire _19961_;
 wire _19962_;
 wire _19963_;
 wire _19964_;
 wire _19965_;
 wire _19966_;
 wire _19967_;
 wire _19968_;
 wire _19969_;
 wire _19970_;
 wire _19971_;
 wire _19972_;
 wire _19973_;
 wire _19974_;
 wire _19975_;
 wire _19976_;
 wire _19977_;
 wire _19978_;
 wire _19979_;
 wire _19980_;
 wire _19981_;
 wire _19982_;
 wire _19983_;
 wire _19984_;
 wire _19985_;
 wire _19986_;
 wire _19987_;
 wire _19988_;
 wire _19989_;
 wire _19990_;
 wire _19991_;
 wire _19992_;
 wire _19993_;
 wire _19994_;
 wire _19995_;
 wire _19996_;
 wire _19997_;
 wire _19998_;
 wire _19999_;
 wire _20000_;
 wire _20001_;
 wire _20002_;
 wire _20003_;
 wire _20004_;
 wire _20005_;
 wire _20006_;
 wire _20007_;
 wire _20008_;
 wire _20009_;
 wire _20010_;
 wire _20011_;
 wire _20012_;
 wire _20013_;
 wire _20014_;
 wire _20015_;
 wire _20016_;
 wire _20017_;
 wire _20018_;
 wire _20019_;
 wire _20020_;
 wire _20021_;
 wire _20022_;
 wire _20023_;
 wire _20024_;
 wire _20025_;
 wire _20026_;
 wire _20027_;
 wire _20028_;
 wire _20029_;
 wire _20030_;
 wire _20031_;
 wire _20032_;
 wire _20033_;
 wire _20034_;
 wire _20035_;
 wire _20036_;
 wire _20037_;
 wire _20038_;
 wire _20039_;
 wire _20040_;
 wire _20041_;
 wire _20042_;
 wire _20043_;
 wire _20044_;
 wire _20045_;
 wire _20046_;
 wire _20047_;
 wire _20048_;
 wire _20049_;
 wire _20050_;
 wire _20051_;
 wire _20052_;
 wire _20053_;
 wire _20054_;
 wire _20055_;
 wire _20056_;
 wire _20057_;
 wire _20058_;
 wire _20059_;
 wire _20060_;
 wire _20061_;
 wire _20062_;
 wire _20063_;
 wire _20064_;
 wire _20065_;
 wire _20066_;
 wire _20067_;
 wire _20068_;
 wire _20069_;
 wire _20070_;
 wire _20071_;
 wire _20072_;
 wire _20073_;
 wire _20074_;
 wire _20075_;
 wire _20076_;
 wire _20077_;
 wire _20078_;
 wire _20079_;
 wire _20080_;
 wire _20081_;
 wire _20082_;
 wire _20083_;
 wire _20084_;
 wire _20085_;
 wire _20086_;
 wire _20087_;
 wire _20088_;
 wire _20089_;
 wire _20090_;
 wire _20091_;
 wire _20092_;
 wire _20093_;
 wire _20094_;
 wire _20095_;
 wire _20096_;
 wire _20097_;
 wire _20098_;
 wire _20099_;
 wire _20100_;
 wire _20101_;
 wire _20102_;
 wire _20103_;
 wire _20104_;
 wire _20105_;
 wire _20106_;
 wire _20107_;
 wire _20108_;
 wire _20109_;
 wire _20110_;
 wire _20111_;
 wire _20112_;
 wire _20113_;
 wire _20114_;
 wire _20115_;
 wire _20116_;
 wire _20117_;
 wire _20118_;
 wire _20119_;
 wire _20120_;
 wire _20121_;
 wire _20122_;
 wire _20123_;
 wire _20124_;
 wire _20125_;
 wire _20126_;
 wire _20127_;
 wire _20128_;
 wire _20129_;
 wire _20130_;
 wire _20131_;
 wire _20132_;
 wire _20133_;
 wire _20134_;
 wire _20135_;
 wire _20136_;
 wire _20137_;
 wire _20138_;
 wire _20139_;
 wire _20140_;
 wire _20141_;
 wire _20142_;
 wire _20143_;
 wire _20144_;
 wire _20145_;
 wire _20146_;
 wire _20147_;
 wire _20148_;
 wire _20149_;
 wire _20150_;
 wire _20151_;
 wire _20152_;
 wire _20153_;
 wire _20154_;
 wire _20155_;
 wire _20156_;
 wire _20157_;
 wire _20158_;
 wire _20159_;
 wire _20160_;
 wire _20161_;
 wire _20162_;
 wire _20163_;
 wire _20164_;
 wire _20165_;
 wire _20166_;
 wire _20167_;
 wire _20168_;
 wire _20169_;
 wire _20170_;
 wire _20171_;
 wire _20172_;
 wire _20173_;
 wire _20174_;
 wire _20175_;
 wire _20176_;
 wire _20177_;
 wire _20178_;
 wire _20179_;
 wire _20180_;
 wire _20181_;
 wire _20182_;
 wire _20183_;
 wire _20184_;
 wire _20185_;
 wire _20186_;
 wire _20187_;
 wire _20188_;
 wire _20189_;
 wire _20190_;
 wire _20191_;
 wire _20192_;
 wire _20193_;
 wire _20194_;
 wire _20195_;
 wire _20196_;
 wire _20197_;
 wire _20198_;
 wire _20199_;
 wire _20200_;
 wire _20201_;
 wire _20202_;
 wire _20203_;
 wire _20204_;
 wire _20205_;
 wire _20206_;
 wire _20207_;
 wire _20208_;
 wire _20209_;
 wire _20210_;
 wire _20211_;
 wire _20212_;
 wire _20213_;
 wire _20214_;
 wire _20215_;
 wire _20216_;
 wire _20217_;
 wire _20218_;
 wire _20219_;
 wire _20220_;
 wire _20221_;
 wire _20222_;
 wire _20223_;
 wire _20224_;
 wire _20225_;
 wire _20226_;
 wire _20227_;
 wire _20228_;
 wire _20229_;
 wire _20230_;
 wire _20231_;
 wire _20232_;
 wire _20233_;
 wire _20234_;
 wire _20235_;
 wire _20236_;
 wire _20237_;
 wire _20238_;
 wire _20239_;
 wire _20240_;
 wire _20241_;
 wire _20242_;
 wire _20243_;
 wire _20244_;
 wire _20245_;
 wire _20246_;
 wire _20247_;
 wire _20248_;
 wire _20249_;
 wire _20250_;
 wire _20251_;
 wire _20252_;
 wire _20253_;
 wire _20254_;
 wire _20255_;
 wire _20256_;
 wire _20257_;
 wire _20258_;
 wire _20259_;
 wire _20260_;
 wire _20261_;
 wire _20262_;
 wire _20263_;
 wire _20264_;
 wire _20265_;
 wire _20266_;
 wire _20267_;
 wire _20268_;
 wire _20269_;
 wire _20270_;
 wire _20271_;
 wire _20272_;
 wire _20273_;
 wire _20274_;
 wire _20275_;
 wire _20276_;
 wire _20277_;
 wire _20278_;
 wire _20279_;
 wire _20280_;
 wire _20281_;
 wire _20282_;
 wire _20283_;
 wire _20284_;
 wire _20285_;
 wire _20286_;
 wire _20287_;
 wire _20288_;
 wire _20289_;
 wire _20290_;
 wire _20291_;
 wire _20292_;
 wire _20293_;
 wire _20294_;
 wire _20295_;
 wire _20296_;
 wire _20297_;
 wire _20298_;
 wire _20299_;
 wire _20300_;
 wire _20301_;
 wire _20302_;
 wire _20303_;
 wire _20304_;
 wire _20305_;
 wire _20306_;
 wire _20307_;
 wire _20308_;
 wire _20309_;
 wire _20310_;
 wire _20311_;
 wire _20312_;
 wire _20313_;
 wire _20314_;
 wire _20315_;
 wire _20316_;
 wire _20317_;
 wire _20318_;
 wire _20319_;
 wire _20320_;
 wire _20321_;
 wire _20322_;
 wire _20323_;
 wire _20324_;
 wire _20325_;
 wire _20326_;
 wire _20327_;
 wire _20328_;
 wire _20329_;
 wire _20330_;
 wire _20331_;
 wire _20332_;
 wire _20333_;
 wire _20334_;
 wire _20335_;
 wire _20336_;
 wire _20337_;
 wire _20338_;
 wire _20339_;
 wire _20340_;
 wire _20341_;
 wire _20342_;
 wire _20343_;
 wire _20344_;
 wire _20345_;
 wire _20346_;
 wire _20347_;
 wire _20348_;
 wire _20349_;
 wire _20350_;
 wire _20351_;
 wire _20352_;
 wire _20353_;
 wire _20354_;
 wire _20355_;
 wire _20356_;
 wire _20357_;
 wire _20358_;
 wire _20359_;
 wire _20360_;
 wire _20361_;
 wire _20362_;
 wire _20363_;
 wire _20364_;
 wire _20365_;
 wire _20366_;
 wire _20367_;
 wire _20368_;
 wire _20369_;
 wire _20370_;
 wire _20371_;
 wire _20372_;
 wire _20373_;
 wire _20374_;
 wire _20375_;
 wire _20376_;
 wire _20377_;
 wire _20378_;
 wire _20379_;
 wire _20380_;
 wire _20381_;
 wire _20382_;
 wire _20383_;
 wire _20384_;
 wire _20385_;
 wire _20386_;
 wire _20387_;
 wire _20388_;
 wire _20389_;
 wire _20390_;
 wire _20391_;
 wire _20392_;
 wire _20393_;
 wire _20394_;
 wire _20395_;
 wire _20396_;
 wire _20397_;
 wire _20398_;
 wire _20399_;
 wire _20400_;
 wire _20401_;
 wire _20402_;
 wire _20403_;
 wire _20404_;
 wire _20405_;
 wire _20406_;
 wire _20407_;
 wire _20408_;
 wire _20409_;
 wire _20410_;
 wire _20411_;
 wire _20412_;
 wire _20413_;
 wire _20414_;
 wire _20415_;
 wire _20416_;
 wire _20417_;
 wire _20418_;
 wire _20419_;
 wire _20420_;
 wire _20421_;
 wire _20422_;
 wire _20423_;
 wire _20424_;
 wire _20425_;
 wire _20426_;
 wire _20427_;
 wire _20428_;
 wire _20429_;
 wire _20430_;
 wire _20431_;
 wire _20432_;
 wire _20433_;
 wire _20434_;
 wire _20435_;
 wire _20436_;
 wire _20437_;
 wire _20438_;
 wire _20439_;
 wire _20440_;
 wire _20441_;
 wire _20442_;
 wire _20443_;
 wire _20444_;
 wire _20445_;
 wire _20446_;
 wire _20447_;
 wire _20448_;
 wire _20449_;
 wire _20450_;
 wire _20451_;
 wire _20452_;
 wire _20453_;
 wire _20454_;
 wire _20455_;
 wire _20456_;
 wire _20457_;
 wire _20458_;
 wire _20459_;
 wire _20460_;
 wire _20461_;
 wire _20462_;
 wire _20463_;
 wire _20464_;
 wire _20465_;
 wire _20466_;
 wire _20467_;
 wire _20468_;
 wire _20469_;
 wire _20470_;
 wire _20471_;
 wire _20472_;
 wire _20473_;
 wire _20474_;
 wire _20475_;
 wire _20476_;
 wire _20477_;
 wire _20478_;
 wire _20479_;
 wire _20480_;
 wire _20481_;
 wire _20482_;
 wire _20483_;
 wire _20484_;
 wire _20485_;
 wire _20486_;
 wire _20487_;
 wire _20488_;
 wire _20489_;
 wire _20490_;
 wire _20491_;
 wire _20492_;
 wire _20493_;
 wire _20494_;
 wire _20495_;
 wire _20496_;
 wire _20497_;
 wire _20498_;
 wire _20499_;
 wire _20500_;
 wire _20501_;
 wire _20502_;
 wire _20503_;
 wire _20504_;
 wire _20505_;
 wire _20506_;
 wire _20507_;
 wire _20508_;
 wire _20509_;
 wire _20510_;
 wire _20511_;
 wire _20512_;
 wire _20513_;
 wire _20514_;
 wire _20515_;
 wire _20516_;
 wire _20517_;
 wire _20518_;
 wire _20519_;
 wire _20520_;
 wire _20521_;
 wire _20522_;
 wire _20523_;
 wire _20524_;
 wire _20525_;
 wire _20526_;
 wire _20527_;
 wire _20528_;
 wire _20529_;
 wire _20530_;
 wire _20531_;
 wire _20532_;
 wire _20533_;
 wire _20534_;
 wire _20535_;
 wire _20536_;
 wire _20537_;
 wire _20538_;
 wire _20539_;
 wire _20540_;
 wire _20541_;
 wire _20542_;
 wire _20543_;
 wire _20544_;
 wire _20545_;
 wire _20546_;
 wire _20547_;
 wire _20548_;
 wire _20549_;
 wire _20550_;
 wire _20551_;
 wire _20552_;
 wire _20553_;
 wire _20554_;
 wire _20555_;
 wire _20556_;
 wire _20557_;
 wire _20558_;
 wire _20559_;
 wire _20560_;
 wire _20561_;
 wire _20562_;
 wire _20563_;
 wire _20564_;
 wire _20565_;
 wire _20566_;
 wire _20567_;
 wire _20568_;
 wire _20569_;
 wire _20570_;
 wire _20571_;
 wire _20572_;
 wire _20573_;
 wire _20574_;
 wire _20575_;
 wire _20576_;
 wire _20577_;
 wire _20578_;
 wire _20579_;
 wire _20580_;
 wire _20581_;
 wire _20582_;
 wire _20583_;
 wire _20584_;
 wire _20585_;
 wire _20586_;
 wire _20587_;
 wire _20588_;
 wire _20589_;
 wire _20590_;
 wire _20591_;
 wire _20592_;
 wire _20593_;
 wire _20594_;
 wire _20595_;
 wire _20596_;
 wire _20597_;
 wire _20598_;
 wire _20599_;
 wire _20600_;
 wire _20601_;
 wire _20602_;
 wire _20603_;
 wire _20604_;
 wire _20605_;
 wire _20606_;
 wire _20607_;
 wire _20608_;
 wire _20609_;
 wire _20610_;
 wire _20611_;
 wire _20612_;
 wire _20613_;
 wire _20614_;
 wire _20615_;
 wire _20616_;
 wire _20617_;
 wire _20618_;
 wire _20619_;
 wire _20620_;
 wire _20621_;
 wire _20622_;
 wire _20623_;
 wire _20624_;
 wire _20625_;
 wire _20626_;
 wire _20627_;
 wire _20628_;
 wire _20629_;
 wire _20630_;
 wire _20631_;
 wire _20632_;
 wire _20633_;
 wire _20634_;
 wire _20635_;
 wire _20636_;
 wire _20637_;
 wire _20638_;
 wire _20639_;
 wire _20640_;
 wire _20641_;
 wire _20642_;
 wire _20643_;
 wire _20644_;
 wire _20645_;
 wire _20646_;
 wire _20647_;
 wire _20648_;
 wire _20649_;
 wire _20650_;
 wire _20651_;
 wire _20652_;
 wire _20653_;
 wire _20654_;
 wire _20655_;
 wire _20656_;
 wire _20657_;
 wire _20658_;
 wire _20659_;
 wire _20660_;
 wire _20661_;
 wire _20662_;
 wire _20663_;
 wire _20664_;
 wire _20665_;
 wire _20666_;
 wire _20667_;
 wire _20668_;
 wire _20669_;
 wire _20670_;
 wire _20671_;
 wire _20672_;
 wire _20673_;
 wire _20674_;
 wire _20675_;
 wire _20676_;
 wire _20677_;
 wire _20678_;
 wire _20679_;
 wire _20680_;
 wire _20681_;
 wire _20682_;
 wire _20683_;
 wire _20684_;
 wire _20685_;
 wire _20686_;
 wire _20687_;
 wire _20688_;
 wire _20689_;
 wire _20690_;
 wire _20691_;
 wire _20692_;
 wire _20693_;
 wire _20694_;
 wire _20695_;
 wire _20696_;
 wire _20697_;
 wire _20698_;
 wire _20699_;
 wire _20700_;
 wire _20701_;
 wire _20702_;
 wire _20703_;
 wire _20704_;
 wire _20705_;
 wire _20706_;
 wire _20707_;
 wire _20708_;
 wire _20709_;
 wire _20710_;
 wire _20711_;
 wire _20712_;
 wire _20713_;
 wire _20714_;
 wire _20715_;
 wire _20716_;
 wire _20717_;
 wire _20718_;
 wire _20719_;
 wire _20720_;
 wire _20721_;
 wire _20722_;
 wire _20723_;
 wire _20724_;
 wire _20725_;
 wire _20726_;
 wire _20727_;
 wire _20728_;
 wire _20729_;
 wire _20730_;
 wire _20731_;
 wire _20732_;
 wire _20733_;
 wire _20734_;
 wire _20735_;
 wire _20736_;
 wire _20737_;
 wire _20738_;
 wire _20739_;
 wire _20740_;
 wire _20741_;
 wire _20742_;
 wire _20743_;
 wire _20744_;
 wire _20745_;
 wire _20746_;
 wire _20747_;
 wire _20748_;
 wire _20749_;
 wire _20750_;
 wire _20751_;
 wire _20752_;
 wire _20753_;
 wire _20754_;
 wire _20755_;
 wire _20756_;
 wire _20757_;
 wire _20758_;
 wire _20759_;
 wire _20760_;
 wire _20761_;
 wire _20762_;
 wire _20763_;
 wire _20764_;
 wire _20765_;
 wire _20766_;
 wire _20767_;
 wire _20768_;
 wire _20769_;
 wire _20770_;
 wire _20771_;
 wire _20772_;
 wire _20773_;
 wire _20774_;
 wire _20775_;
 wire _20776_;
 wire _20777_;
 wire _20778_;
 wire _20779_;
 wire _20780_;
 wire _20781_;
 wire _20782_;
 wire _20783_;
 wire _20784_;
 wire _20785_;
 wire _20786_;
 wire _20787_;
 wire _20788_;
 wire _20789_;
 wire _20790_;
 wire _20791_;
 wire _20792_;
 wire _20793_;
 wire _20794_;
 wire _20795_;
 wire _20796_;
 wire _20797_;
 wire _20798_;
 wire _20799_;
 wire _20800_;
 wire _20801_;
 wire _20802_;
 wire _20803_;
 wire _20804_;
 wire _20805_;
 wire _20806_;
 wire _20807_;
 wire _20808_;
 wire _20809_;
 wire _20810_;
 wire _20811_;
 wire _20812_;
 wire _20813_;
 wire _20814_;
 wire _20815_;
 wire _20816_;
 wire _20817_;
 wire _20818_;
 wire _20819_;
 wire _20820_;
 wire _20821_;
 wire _20822_;
 wire _20823_;
 wire _20824_;
 wire _20825_;
 wire _20826_;
 wire _20827_;
 wire _20828_;
 wire _20829_;
 wire _20830_;
 wire _20831_;
 wire _20832_;
 wire _20833_;
 wire _20834_;
 wire _20835_;
 wire _20836_;
 wire _20837_;
 wire _20838_;
 wire _20839_;
 wire _20840_;
 wire _20841_;
 wire _20842_;
 wire _20843_;
 wire _20844_;
 wire _20845_;
 wire _20846_;
 wire _20847_;
 wire _20848_;
 wire _20849_;
 wire _20850_;
 wire _20851_;
 wire _20852_;
 wire _20853_;
 wire _20854_;
 wire _20855_;
 wire _20856_;
 wire _20857_;
 wire _20858_;
 wire _20859_;
 wire _20860_;
 wire _20861_;
 wire _20862_;
 wire _20863_;
 wire _20864_;
 wire _20865_;
 wire _20866_;
 wire _20867_;
 wire _20868_;
 wire _20869_;
 wire _20870_;
 wire _20871_;
 wire _20872_;
 wire _20873_;
 wire _20874_;
 wire _20875_;
 wire _20876_;
 wire _20877_;
 wire _20878_;
 wire _20879_;
 wire _20880_;
 wire _20881_;
 wire _20882_;
 wire _20883_;
 wire _20884_;
 wire _20885_;
 wire _20886_;
 wire _20887_;
 wire _20888_;
 wire _20889_;
 wire _20890_;
 wire _20891_;
 wire _20892_;
 wire _20893_;
 wire _20894_;
 wire _20895_;
 wire _20896_;
 wire _20897_;
 wire _20898_;
 wire _20899_;
 wire _20900_;
 wire _20901_;
 wire _20902_;
 wire _20903_;
 wire _20904_;
 wire _20905_;
 wire _20906_;
 wire _20907_;
 wire _20908_;
 wire _20909_;
 wire _20910_;
 wire _20911_;
 wire _20912_;
 wire _20913_;
 wire _20914_;
 wire _20915_;
 wire _20916_;
 wire _20917_;
 wire _20918_;
 wire _20919_;
 wire _20920_;
 wire _20921_;
 wire _20922_;
 wire _20923_;
 wire _20924_;
 wire _20925_;
 wire _20926_;
 wire _20927_;
 wire _20928_;
 wire _20929_;
 wire _20930_;
 wire _20931_;
 wire _20932_;
 wire _20933_;
 wire _20934_;
 wire _20935_;
 wire _20936_;
 wire _20937_;
 wire _20938_;
 wire _20939_;
 wire _20940_;
 wire _20941_;
 wire _20942_;
 wire _20943_;
 wire _20944_;
 wire _20945_;
 wire _20946_;
 wire _20947_;
 wire _20948_;
 wire _20949_;
 wire _20950_;
 wire _20951_;
 wire _20952_;
 wire _20953_;
 wire _20954_;
 wire _20955_;
 wire _20956_;
 wire _20957_;
 wire _20958_;
 wire _20959_;
 wire _20960_;
 wire _20961_;
 wire _20962_;
 wire _20963_;
 wire _20964_;
 wire _20965_;
 wire _20966_;
 wire _20967_;
 wire _20968_;
 wire _20969_;
 wire _20970_;
 wire _20971_;
 wire _20972_;
 wire _20973_;
 wire _20974_;
 wire _20975_;
 wire _20976_;
 wire _20977_;
 wire _20978_;
 wire _20979_;
 wire _20980_;
 wire _20981_;
 wire _20982_;
 wire _20983_;
 wire _20984_;
 wire _20985_;
 wire _20986_;
 wire _20987_;
 wire _20988_;
 wire _20989_;
 wire _20990_;
 wire _20991_;
 wire _20992_;
 wire _20993_;
 wire _20994_;
 wire _20995_;
 wire _20996_;
 wire _20997_;
 wire _20998_;
 wire _20999_;
 wire _21000_;
 wire _21001_;
 wire _21002_;
 wire _21003_;
 wire _21004_;
 wire _21005_;
 wire _21006_;
 wire _21007_;
 wire _21008_;
 wire _21009_;
 wire _21010_;
 wire _21011_;
 wire _21012_;
 wire _21013_;
 wire _21014_;
 wire _21015_;
 wire _21016_;
 wire _21017_;
 wire _21018_;
 wire _21019_;
 wire _21020_;
 wire _21021_;
 wire _21022_;
 wire _21023_;
 wire _21024_;
 wire _21025_;
 wire _21026_;
 wire _21027_;
 wire _21028_;
 wire _21029_;
 wire _21030_;
 wire _21031_;
 wire _21032_;
 wire _21033_;
 wire _21034_;
 wire _21035_;
 wire _21036_;
 wire _21037_;
 wire _21038_;
 wire _21039_;
 wire _21040_;
 wire _21041_;
 wire _21042_;
 wire _21043_;
 wire _21044_;
 wire _21045_;
 wire _21046_;
 wire _21047_;
 wire _21048_;
 wire _21049_;
 wire _21050_;
 wire _21051_;
 wire _21052_;
 wire _21053_;
 wire _21054_;
 wire _21055_;
 wire _21056_;
 wire _21057_;
 wire _21058_;
 wire _21059_;
 wire _21060_;
 wire _21061_;
 wire _21062_;
 wire _21063_;
 wire _21064_;
 wire _21065_;
 wire _21066_;
 wire _21067_;
 wire _21068_;
 wire _21069_;
 wire _21070_;
 wire _21071_;
 wire _21072_;
 wire _21073_;
 wire _21074_;
 wire _21075_;
 wire _21076_;
 wire _21077_;
 wire _21078_;
 wire _21079_;
 wire _21080_;
 wire _21081_;
 wire _21082_;
 wire _21083_;
 wire _21084_;
 wire _21085_;
 wire _21086_;
 wire _21087_;
 wire _21088_;
 wire _21089_;
 wire _21090_;
 wire _21091_;
 wire _21092_;
 wire _21093_;
 wire _21094_;
 wire _21095_;
 wire _21096_;
 wire _21097_;
 wire _21098_;
 wire _21099_;
 wire _21100_;
 wire _21101_;
 wire _21102_;
 wire _21103_;
 wire _21104_;
 wire _21105_;
 wire _21106_;
 wire _21107_;
 wire _21108_;
 wire _21109_;
 wire _21110_;
 wire _21111_;
 wire _21112_;
 wire _21113_;
 wire _21114_;
 wire _21115_;
 wire _21116_;
 wire _21117_;
 wire _21118_;
 wire _21119_;
 wire _21120_;
 wire _21121_;
 wire _21122_;
 wire _21123_;
 wire _21124_;
 wire _21125_;
 wire _21126_;
 wire _21127_;
 wire _21128_;
 wire _21129_;
 wire _21130_;
 wire _21131_;
 wire _21132_;
 wire _21133_;
 wire _21134_;
 wire _21135_;
 wire _21136_;
 wire _21137_;
 wire _21138_;
 wire _21139_;
 wire _21140_;
 wire _21141_;
 wire _21142_;
 wire _21143_;
 wire _21144_;
 wire _21145_;
 wire _21146_;
 wire _21147_;
 wire _21148_;
 wire _21149_;
 wire _21150_;
 wire _21151_;
 wire _21152_;
 wire _21153_;
 wire _21154_;
 wire _21155_;
 wire _21156_;
 wire _21157_;
 wire _21158_;
 wire _21159_;
 wire _21160_;
 wire _21161_;
 wire _21162_;
 wire _21163_;
 wire _21164_;
 wire _21165_;
 wire _21166_;
 wire _21167_;
 wire _21168_;
 wire _21169_;
 wire _21170_;
 wire _21171_;
 wire _21172_;
 wire _21173_;
 wire _21174_;
 wire _21175_;
 wire _21176_;
 wire _21177_;
 wire _21178_;
 wire _21179_;
 wire _21180_;
 wire _21181_;
 wire _21182_;
 wire _21183_;
 wire _21184_;
 wire _21185_;
 wire _21186_;
 wire _21187_;
 wire _21188_;
 wire _21189_;
 wire _21190_;
 wire _21191_;
 wire _21192_;
 wire _21193_;
 wire _21194_;
 wire _21195_;
 wire _21196_;
 wire _21197_;
 wire _21198_;
 wire _21199_;
 wire _21200_;
 wire _21201_;
 wire _21202_;
 wire _21203_;
 wire _21204_;
 wire _21205_;
 wire _21206_;
 wire _21207_;
 wire _21208_;
 wire _21209_;
 wire _21210_;
 wire _21211_;
 wire _21212_;
 wire _21213_;
 wire _21214_;
 wire _21215_;
 wire _21216_;
 wire _21217_;
 wire _21218_;
 wire _21219_;
 wire _21220_;
 wire _21221_;
 wire _21222_;
 wire _21223_;
 wire _21224_;
 wire _21225_;
 wire _21226_;
 wire _21227_;
 wire _21228_;
 wire _21229_;
 wire _21230_;
 wire _21231_;
 wire _21232_;
 wire _21233_;
 wire _21234_;
 wire _21235_;
 wire _21236_;
 wire _21237_;
 wire _21238_;
 wire _21239_;
 wire _21240_;
 wire _21241_;
 wire _21242_;
 wire _21243_;
 wire _21244_;
 wire _21245_;
 wire _21246_;
 wire _21247_;
 wire _21248_;
 wire _21249_;
 wire _21250_;
 wire _21251_;
 wire _21252_;
 wire _21253_;
 wire _21254_;
 wire _21255_;
 wire _21256_;
 wire _21257_;
 wire _21258_;
 wire _21259_;
 wire _21260_;
 wire _21261_;
 wire _21262_;
 wire _21263_;
 wire _21264_;
 wire _21265_;
 wire _21266_;
 wire _21267_;
 wire _21268_;
 wire _21269_;
 wire _21270_;
 wire _21271_;
 wire _21272_;
 wire _21273_;
 wire _21274_;
 wire _21275_;
 wire _21276_;
 wire _21277_;
 wire _21278_;
 wire _21279_;
 wire _21280_;
 wire _21281_;
 wire _21282_;
 wire _21283_;
 wire _21284_;
 wire _21285_;
 wire _21286_;
 wire _21287_;
 wire _21288_;
 wire _21289_;
 wire _21290_;
 wire _21291_;
 wire _21292_;
 wire _21293_;
 wire _21294_;
 wire _21295_;
 wire _21296_;
 wire _21297_;
 wire _21298_;
 wire _21299_;
 wire _21300_;
 wire _21301_;
 wire _21302_;
 wire _21303_;
 wire _21304_;
 wire _21305_;
 wire _21306_;
 wire _21307_;
 wire _21308_;
 wire _21309_;
 wire _21310_;
 wire _21311_;
 wire _21312_;
 wire _21313_;
 wire _21314_;
 wire _21315_;
 wire _21316_;
 wire _21317_;
 wire _21318_;
 wire _21319_;
 wire _21320_;
 wire _21321_;
 wire _21322_;
 wire _21323_;
 wire _21324_;
 wire _21325_;
 wire _21326_;
 wire _21327_;
 wire _21328_;
 wire _21329_;
 wire _21330_;
 wire _21331_;
 wire _21332_;
 wire _21333_;
 wire _21334_;
 wire _21335_;
 wire _21336_;
 wire _21337_;
 wire _21338_;
 wire _21339_;
 wire _21340_;
 wire _21341_;
 wire _21342_;
 wire _21343_;
 wire _21344_;
 wire _21345_;
 wire _21346_;
 wire _21347_;
 wire _21348_;
 wire _21349_;
 wire _21350_;
 wire _21351_;
 wire _21352_;
 wire _21353_;
 wire _21354_;
 wire _21355_;
 wire _21356_;
 wire _21357_;
 wire _21358_;
 wire _21359_;
 wire _21360_;
 wire _21361_;
 wire _21362_;
 wire _21363_;
 wire _21364_;
 wire _21365_;
 wire _21366_;
 wire _21367_;
 wire _21368_;
 wire _21369_;
 wire _21370_;
 wire _21371_;
 wire _21372_;
 wire _21373_;
 wire _21374_;
 wire _21375_;
 wire _21376_;
 wire _21377_;
 wire _21378_;
 wire _21379_;
 wire _21380_;
 wire _21381_;
 wire _21382_;
 wire _21383_;
 wire _21384_;
 wire _21385_;
 wire _21386_;
 wire _21387_;
 wire _21388_;
 wire _21389_;
 wire _21390_;
 wire _21391_;
 wire _21392_;
 wire _21393_;
 wire _21394_;
 wire _21395_;
 wire _21396_;
 wire _21397_;
 wire _21398_;
 wire _21399_;
 wire _21400_;
 wire _21401_;
 wire _21402_;
 wire _21403_;
 wire _21404_;
 wire _21405_;
 wire _21406_;
 wire _21407_;
 wire _21408_;
 wire _21409_;
 wire _21410_;
 wire _21411_;
 wire _21412_;
 wire _21413_;
 wire _21414_;
 wire _21415_;
 wire _21416_;
 wire _21417_;
 wire _21418_;
 wire _21419_;
 wire _21420_;
 wire _21421_;
 wire _21422_;
 wire _21423_;
 wire _21424_;
 wire _21425_;
 wire _21426_;
 wire _21427_;
 wire _21428_;
 wire _21429_;
 wire _21430_;
 wire _21431_;
 wire _21432_;
 wire _21433_;
 wire _21434_;
 wire _21435_;
 wire _21436_;
 wire _21437_;
 wire _21438_;
 wire _21439_;
 wire _21440_;
 wire _21441_;
 wire _21442_;
 wire _21443_;
 wire _21444_;
 wire _21445_;
 wire _21446_;
 wire _21447_;
 wire _21448_;
 wire _21449_;
 wire _21450_;
 wire _21451_;
 wire _21452_;
 wire _21453_;
 wire _21454_;
 wire _21455_;
 wire _21456_;
 wire _21457_;
 wire _21458_;
 wire _21459_;
 wire _21460_;
 wire _21461_;
 wire _21462_;
 wire _21463_;
 wire _21464_;
 wire _21465_;
 wire _21466_;
 wire _21467_;
 wire _21468_;
 wire _21469_;
 wire _21470_;
 wire _21471_;
 wire _21472_;
 wire _21473_;
 wire _21474_;
 wire _21475_;
 wire _21476_;
 wire _21477_;
 wire _21478_;
 wire _21479_;
 wire _21480_;
 wire _21481_;
 wire _21482_;
 wire _21483_;
 wire _21484_;
 wire _21485_;
 wire _21486_;
 wire _21487_;
 wire _21488_;
 wire _21489_;
 wire _21490_;
 wire _21491_;
 wire _21492_;
 wire _21493_;
 wire _21494_;
 wire _21495_;
 wire _21496_;
 wire _21497_;
 wire _21498_;
 wire _21499_;
 wire _21500_;
 wire _21501_;
 wire _21502_;
 wire _21503_;
 wire _21504_;
 wire _21505_;
 wire _21506_;
 wire _21507_;
 wire _21508_;
 wire _21509_;
 wire _21510_;
 wire _21511_;
 wire _21512_;
 wire _21513_;
 wire _21514_;
 wire _21515_;
 wire _21516_;
 wire _21517_;
 wire _21518_;
 wire _21519_;
 wire _21520_;
 wire _21521_;
 wire _21522_;
 wire _21523_;
 wire _21524_;
 wire _21525_;
 wire _21526_;
 wire _21527_;
 wire _21528_;
 wire _21529_;
 wire _21530_;
 wire _21531_;
 wire _21532_;
 wire _21533_;
 wire _21534_;
 wire _21535_;
 wire _21536_;
 wire _21537_;
 wire _21538_;
 wire _21539_;
 wire _21540_;
 wire _21541_;
 wire _21542_;
 wire _21543_;
 wire _21544_;
 wire _21545_;
 wire _21546_;
 wire _21547_;
 wire _21548_;
 wire _21549_;
 wire _21550_;
 wire _21551_;
 wire _21552_;
 wire _21553_;
 wire _21554_;
 wire _21555_;
 wire _21556_;
 wire _21557_;
 wire _21558_;
 wire _21559_;
 wire _21560_;
 wire _21561_;
 wire _21562_;
 wire _21563_;
 wire _21564_;
 wire _21565_;
 wire _21566_;
 wire _21567_;
 wire _21568_;
 wire _21569_;
 wire _21570_;
 wire _21571_;
 wire _21572_;
 wire _21573_;
 wire _21574_;
 wire _21575_;
 wire _21576_;
 wire _21577_;
 wire _21578_;
 wire _21579_;
 wire _21580_;
 wire _21581_;
 wire _21582_;
 wire _21583_;
 wire _21584_;
 wire _21585_;
 wire _21586_;
 wire _21587_;
 wire _21588_;
 wire _21589_;
 wire _21590_;
 wire _21591_;
 wire _21592_;
 wire _21593_;
 wire _21594_;
 wire _21595_;
 wire _21596_;
 wire _21597_;
 wire _21598_;
 wire _21599_;
 wire _21600_;
 wire _21601_;
 wire _21602_;
 wire _21603_;
 wire _21604_;
 wire _21605_;
 wire _21606_;
 wire _21607_;
 wire _21608_;
 wire _21609_;
 wire _21610_;
 wire _21611_;
 wire _21612_;
 wire _21613_;
 wire _21614_;
 wire _21615_;
 wire _21616_;
 wire _21617_;
 wire _21618_;
 wire _21619_;
 wire _21620_;
 wire _21621_;
 wire _21622_;
 wire _21623_;
 wire _21624_;
 wire _21625_;
 wire _21626_;
 wire _21627_;
 wire _21628_;
 wire _21629_;
 wire _21630_;
 wire _21631_;
 wire _21632_;
 wire _21633_;
 wire _21634_;
 wire _21635_;
 wire _21636_;
 wire _21637_;
 wire _21638_;
 wire _21639_;
 wire _21640_;
 wire _21641_;
 wire _21642_;
 wire _21643_;
 wire _21644_;
 wire _21645_;
 wire _21646_;
 wire _21647_;
 wire _21648_;
 wire _21649_;
 wire _21650_;
 wire _21651_;
 wire _21652_;
 wire _21653_;
 wire _21654_;
 wire _21655_;
 wire _21656_;
 wire _21657_;
 wire _21658_;
 wire _21659_;
 wire _21660_;
 wire _21661_;
 wire _21662_;
 wire _21663_;
 wire _21664_;
 wire _21665_;
 wire _21666_;
 wire _21667_;
 wire _21668_;
 wire _21669_;
 wire _21670_;
 wire _21671_;
 wire _21672_;
 wire _21673_;
 wire _21674_;
 wire _21675_;
 wire _21676_;
 wire _21677_;
 wire _21678_;
 wire _21679_;
 wire _21680_;
 wire _21681_;
 wire _21682_;
 wire _21683_;
 wire _21684_;
 wire _21685_;
 wire _21686_;
 wire _21687_;
 wire _21688_;
 wire _21689_;
 wire _21690_;
 wire _21691_;
 wire _21692_;
 wire _21693_;
 wire _21694_;
 wire _21695_;
 wire _21696_;
 wire _21697_;
 wire _21698_;
 wire _21699_;
 wire _21700_;
 wire _21701_;
 wire _21702_;
 wire _21703_;
 wire _21704_;
 wire _21705_;
 wire _21706_;
 wire _21707_;
 wire _21708_;
 wire _21709_;
 wire _21710_;
 wire _21711_;
 wire _21712_;
 wire _21713_;
 wire _21714_;
 wire _21715_;
 wire _21716_;
 wire _21717_;
 wire _21718_;
 wire _21719_;
 wire _21720_;
 wire _21721_;
 wire _21722_;
 wire _21723_;
 wire _21724_;
 wire _21725_;
 wire _21726_;
 wire _21727_;
 wire _21728_;
 wire _21729_;
 wire _21730_;
 wire _21731_;
 wire _21732_;
 wire _21733_;
 wire _21734_;
 wire _21735_;
 wire _21736_;
 wire _21737_;
 wire _21738_;
 wire _21739_;
 wire _21740_;
 wire _21741_;
 wire _21742_;
 wire _21743_;
 wire _21744_;
 wire _21745_;
 wire _21746_;
 wire _21747_;
 wire _21748_;
 wire _21749_;
 wire _21750_;
 wire _21751_;
 wire _21752_;
 wire _21753_;
 wire _21754_;
 wire _21755_;
 wire _21756_;
 wire _21757_;
 wire _21758_;
 wire _21759_;
 wire _21760_;
 wire _21761_;
 wire _21762_;
 wire _21763_;
 wire _21764_;
 wire _21765_;
 wire _21766_;
 wire _21767_;
 wire _21768_;
 wire _21769_;
 wire _21770_;
 wire _21771_;
 wire _21772_;
 wire _21773_;
 wire _21774_;
 wire _21775_;
 wire _21776_;
 wire _21777_;
 wire _21778_;
 wire _21779_;
 wire _21780_;
 wire _21781_;
 wire _21782_;
 wire _21783_;
 wire _21784_;
 wire _21785_;
 wire _21786_;
 wire _21787_;
 wire _21788_;
 wire _21789_;
 wire _21790_;
 wire _21791_;
 wire _21792_;
 wire _21793_;
 wire _21794_;
 wire _21795_;
 wire _21796_;
 wire _21797_;
 wire _21798_;
 wire _21799_;
 wire _21800_;
 wire _21801_;
 wire _21802_;
 wire _21803_;
 wire _21804_;
 wire _21805_;
 wire _21806_;
 wire _21807_;
 wire _21808_;
 wire _21809_;
 wire _21810_;
 wire _21811_;
 wire _21812_;
 wire _21813_;
 wire _21814_;
 wire _21815_;
 wire _21816_;
 wire _21817_;
 wire _21818_;
 wire _21819_;
 wire _21820_;
 wire _21821_;
 wire _21822_;
 wire _21823_;
 wire _21824_;
 wire _21825_;
 wire _21826_;
 wire _21827_;
 wire _21828_;
 wire _21829_;
 wire _21830_;
 wire _21831_;
 wire _21832_;
 wire _21833_;
 wire _21834_;
 wire _21835_;
 wire _21836_;
 wire _21837_;
 wire _21838_;
 wire _21839_;
 wire _21840_;
 wire _21841_;
 wire _21842_;
 wire _21843_;
 wire _21844_;
 wire _21845_;
 wire _21846_;
 wire _21847_;
 wire _21848_;
 wire _21849_;
 wire _21850_;
 wire _21851_;
 wire _21852_;
 wire _21853_;
 wire _21854_;
 wire _21855_;
 wire _21856_;
 wire _21857_;
 wire _21858_;
 wire _21859_;
 wire _21860_;
 wire _21861_;
 wire _21862_;
 wire _21863_;
 wire _21864_;
 wire _21865_;
 wire _21866_;
 wire _21867_;
 wire _21868_;
 wire _21869_;
 wire _21870_;
 wire _21871_;
 wire _21872_;
 wire _21873_;
 wire _21874_;
 wire _21875_;
 wire _21876_;
 wire _21877_;
 wire _21878_;
 wire _21879_;
 wire _21880_;
 wire _21881_;
 wire _21882_;
 wire _21883_;
 wire _21884_;
 wire _21885_;
 wire _21886_;
 wire _21887_;
 wire _21888_;
 wire _21889_;
 wire _21890_;
 wire _21891_;
 wire _21892_;
 wire _21893_;
 wire _21894_;
 wire _21895_;
 wire _21896_;
 wire _21897_;
 wire _21898_;
 wire _21899_;
 wire _21900_;
 wire _21901_;
 wire _21902_;
 wire _21903_;
 wire _21904_;
 wire _21905_;
 wire _21906_;
 wire _21907_;
 wire _21908_;
 wire _21909_;
 wire _21910_;
 wire _21911_;
 wire _21912_;
 wire _21913_;
 wire _21914_;
 wire _21915_;
 wire _21916_;
 wire _21917_;
 wire _21918_;
 wire _21919_;
 wire _21920_;
 wire _21921_;
 wire _21922_;
 wire _21923_;
 wire _21924_;
 wire _21925_;
 wire _21926_;
 wire _21927_;
 wire _21928_;
 wire _21929_;
 wire _21930_;
 wire _21931_;
 wire _21932_;
 wire _21933_;
 wire _21934_;
 wire _21935_;
 wire _21936_;
 wire _21937_;
 wire _21938_;
 wire _21939_;
 wire _21940_;
 wire _21941_;
 wire _21942_;
 wire _21943_;
 wire _21944_;
 wire _21945_;
 wire _21946_;
 wire _21947_;
 wire _21948_;
 wire _21949_;
 wire _21950_;
 wire _21951_;
 wire _21952_;
 wire _21953_;
 wire _21954_;
 wire _21955_;
 wire _21956_;
 wire _21957_;
 wire _21958_;
 wire _21959_;
 wire _21960_;
 wire _21961_;
 wire _21962_;
 wire _21963_;
 wire _21964_;
 wire _21965_;
 wire _21966_;
 wire _21967_;
 wire _21968_;
 wire _21969_;
 wire _21970_;
 wire _21971_;
 wire _21972_;
 wire _21973_;
 wire _21974_;
 wire _21975_;
 wire _21976_;
 wire _21977_;
 wire _21978_;
 wire _21979_;
 wire _21980_;
 wire _21981_;
 wire _21982_;
 wire _21983_;
 wire _21984_;
 wire _21985_;
 wire _21986_;
 wire _21987_;
 wire _21988_;
 wire _21989_;
 wire _21990_;
 wire _21991_;
 wire _21992_;
 wire _21993_;
 wire _21994_;
 wire _21995_;
 wire _21996_;
 wire _21997_;
 wire _21998_;
 wire _21999_;
 wire _22000_;
 wire _22001_;
 wire _22002_;
 wire _22003_;
 wire _22004_;
 wire _22005_;
 wire _22006_;
 wire _22007_;
 wire _22008_;
 wire _22009_;
 wire _22010_;
 wire _22011_;
 wire _22012_;
 wire _22013_;
 wire _22014_;
 wire _22015_;
 wire _22016_;
 wire _22017_;
 wire _22018_;
 wire _22019_;
 wire _22020_;
 wire _22021_;
 wire _22022_;
 wire _22023_;
 wire _22024_;
 wire _22025_;
 wire _22026_;
 wire _22027_;
 wire _22028_;
 wire _22029_;
 wire _22030_;
 wire _22031_;
 wire _22032_;
 wire _22033_;
 wire _22034_;
 wire _22035_;
 wire _22036_;
 wire _22037_;
 wire _22038_;
 wire _22039_;
 wire _22040_;
 wire _22041_;
 wire _22042_;
 wire _22043_;
 wire _22044_;
 wire _22045_;
 wire _22046_;
 wire _22047_;
 wire _22048_;
 wire _22049_;
 wire _22050_;
 wire _22051_;
 wire _22052_;
 wire _22053_;
 wire _22054_;
 wire _22055_;
 wire _22056_;
 wire _22057_;
 wire _22058_;
 wire _22059_;
 wire _22060_;
 wire _22061_;
 wire _22062_;
 wire _22063_;
 wire _22064_;
 wire _22065_;
 wire _22066_;
 wire _22067_;
 wire _22068_;
 wire _22069_;
 wire _22070_;
 wire _22071_;
 wire _22072_;
 wire _22073_;
 wire _22074_;
 wire _22075_;
 wire _22076_;
 wire _22077_;
 wire _22078_;
 wire _22079_;
 wire _22080_;
 wire _22081_;
 wire _22082_;
 wire _22083_;
 wire _22084_;
 wire _22085_;
 wire _22086_;
 wire _22087_;
 wire _22088_;
 wire _22089_;
 wire _22090_;
 wire _22091_;
 wire _22092_;
 wire _22093_;
 wire _22094_;
 wire _22095_;
 wire _22096_;
 wire _22097_;
 wire _22098_;
 wire _22099_;
 wire _22100_;
 wire _22101_;
 wire _22102_;
 wire _22103_;
 wire _22104_;
 wire _22105_;
 wire _22106_;
 wire _22107_;
 wire _22108_;
 wire _22109_;
 wire _22110_;
 wire _22111_;
 wire _22112_;
 wire _22113_;
 wire _22114_;
 wire _22115_;
 wire _22116_;
 wire _22117_;
 wire _22118_;
 wire _22119_;
 wire _22120_;
 wire _22121_;
 wire _22122_;
 wire _22123_;
 wire _22124_;
 wire _22125_;
 wire _22126_;
 wire _22127_;
 wire _22128_;
 wire _22129_;
 wire _22130_;
 wire _22131_;
 wire _22132_;
 wire _22133_;
 wire _22134_;
 wire _22135_;
 wire _22136_;
 wire _22137_;
 wire _22138_;
 wire _22139_;
 wire _22140_;
 wire _22141_;
 wire _22142_;
 wire _22143_;
 wire _22144_;
 wire _22145_;
 wire _22146_;
 wire _22147_;
 wire _22148_;
 wire _22149_;
 wire _22150_;
 wire _22151_;
 wire _22152_;
 wire _22153_;
 wire _22154_;
 wire _22155_;
 wire _22156_;
 wire _22157_;
 wire _22158_;
 wire _22159_;
 wire _22160_;
 wire _22161_;
 wire _22162_;
 wire _22163_;
 wire _22164_;
 wire _22165_;
 wire _22166_;
 wire _22167_;
 wire _22168_;
 wire _22169_;
 wire _22170_;
 wire _22171_;
 wire _22172_;
 wire _22173_;
 wire _22174_;
 wire _22175_;
 wire _22176_;
 wire _22177_;
 wire _22178_;
 wire _22179_;
 wire _22180_;
 wire _22181_;
 wire _22182_;
 wire _22183_;
 wire _22184_;
 wire _22185_;
 wire _22186_;
 wire _22187_;
 wire _22188_;
 wire _22189_;
 wire _22190_;
 wire _22191_;
 wire _22192_;
 wire _22193_;
 wire _22194_;
 wire _22195_;
 wire _22196_;
 wire _22197_;
 wire _22198_;
 wire _22199_;
 wire _22200_;
 wire _22201_;
 wire _22202_;
 wire _22203_;
 wire _22204_;
 wire _22205_;
 wire _22206_;
 wire _22207_;
 wire _22208_;
 wire _22209_;
 wire _22210_;
 wire _22211_;
 wire _22212_;
 wire _22213_;
 wire _22214_;
 wire _22215_;
 wire _22216_;
 wire _22217_;
 wire _22218_;
 wire _22219_;
 wire _22220_;
 wire _22221_;
 wire _22222_;
 wire _22223_;
 wire _22224_;
 wire _22225_;
 wire _22226_;
 wire _22227_;
 wire _22228_;
 wire _22229_;
 wire _22230_;
 wire _22231_;
 wire _22232_;
 wire _22233_;
 wire _22234_;
 wire _22235_;
 wire _22236_;
 wire _22237_;
 wire _22238_;
 wire _22239_;
 wire _22240_;
 wire _22241_;
 wire _22242_;
 wire _22243_;
 wire _22244_;
 wire _22245_;
 wire _22246_;
 wire _22247_;
 wire _22248_;
 wire _22249_;
 wire _22250_;
 wire _22251_;
 wire _22252_;
 wire _22253_;
 wire _22254_;
 wire _22255_;
 wire _22256_;
 wire _22257_;
 wire _22258_;
 wire _22259_;
 wire _22260_;
 wire _22261_;
 wire _22262_;
 wire _22263_;
 wire _22264_;
 wire _22265_;
 wire _22266_;
 wire _22267_;
 wire _22268_;
 wire _22269_;
 wire _22270_;
 wire _22271_;
 wire _22272_;
 wire _22273_;
 wire _22274_;
 wire _22275_;
 wire _22276_;
 wire _22277_;
 wire _22278_;
 wire _22279_;
 wire _22280_;
 wire _22281_;
 wire _22282_;
 wire _22283_;
 wire _22284_;
 wire _22285_;
 wire _22286_;
 wire _22287_;
 wire _22288_;
 wire _22289_;
 wire _22290_;
 wire _22291_;
 wire _22292_;
 wire _22293_;
 wire _22294_;
 wire _22295_;
 wire _22296_;
 wire _22297_;
 wire _22298_;
 wire _22299_;
 wire _22300_;
 wire _22301_;
 wire _22302_;
 wire _22303_;
 wire _22304_;
 wire _22305_;
 wire _22306_;
 wire _22307_;
 wire _22308_;
 wire _22309_;
 wire _22310_;
 wire _22311_;
 wire _22312_;
 wire _22313_;
 wire _22314_;
 wire _22315_;
 wire _22316_;
 wire _22317_;
 wire _22318_;
 wire _22319_;
 wire _22320_;
 wire _22321_;
 wire _22322_;
 wire _22323_;
 wire _22324_;
 wire _22325_;
 wire _22326_;
 wire _22327_;
 wire _22328_;
 wire _22329_;
 wire _22330_;
 wire _22331_;
 wire _22332_;
 wire _22333_;
 wire _22334_;
 wire _22335_;
 wire _22336_;
 wire _22337_;
 wire _22338_;
 wire _22339_;
 wire _22340_;
 wire _22341_;
 wire _22342_;
 wire _22343_;
 wire _22344_;
 wire _22345_;
 wire _22346_;
 wire _22347_;
 wire _22348_;
 wire _22349_;
 wire _22350_;
 wire _22351_;
 wire _22352_;
 wire _22353_;
 wire _22354_;
 wire _22355_;
 wire _22356_;
 wire _22357_;
 wire _22358_;
 wire _22359_;
 wire _22360_;
 wire _22361_;
 wire _22362_;
 wire _22363_;
 wire _22364_;
 wire _22365_;
 wire _22366_;
 wire _22367_;
 wire _22368_;
 wire _22369_;
 wire _22370_;
 wire _22371_;
 wire _22372_;
 wire _22373_;
 wire _22374_;
 wire _22375_;
 wire _22376_;
 wire _22377_;
 wire _22378_;
 wire _22379_;
 wire _22380_;
 wire _22381_;
 wire _22382_;
 wire _22383_;
 wire _22384_;
 wire _22385_;
 wire _22386_;
 wire _22387_;
 wire _22388_;
 wire _22389_;
 wire _22390_;
 wire _22391_;
 wire _22392_;
 wire _22393_;
 wire _22394_;
 wire _22395_;
 wire _22396_;
 wire _22397_;
 wire _22398_;
 wire _22399_;
 wire _22400_;
 wire _22401_;
 wire _22402_;
 wire _22403_;
 wire _22404_;
 wire _22405_;
 wire _22406_;
 wire _22407_;
 wire _22408_;
 wire _22409_;
 wire _22410_;
 wire _22411_;
 wire _22412_;
 wire _22413_;
 wire _22414_;
 wire _22415_;
 wire _22416_;
 wire _22417_;
 wire _22418_;
 wire _22419_;
 wire _22420_;
 wire _22421_;
 wire _22422_;
 wire _22423_;
 wire _22424_;
 wire _22425_;
 wire _22426_;
 wire _22427_;
 wire _22428_;
 wire _22429_;
 wire _22430_;
 wire _22431_;
 wire _22432_;
 wire _22433_;
 wire _22434_;
 wire _22435_;
 wire _22436_;
 wire _22437_;
 wire _22438_;
 wire _22439_;
 wire _22440_;
 wire _22441_;
 wire _22442_;
 wire _22443_;
 wire _22444_;
 wire _22445_;
 wire _22446_;
 wire _22447_;
 wire _22448_;
 wire _22449_;
 wire _22450_;
 wire _22451_;
 wire _22452_;
 wire _22453_;
 wire _22454_;
 wire _22455_;
 wire _22456_;
 wire _22457_;
 wire _22458_;
 wire _22459_;
 wire _22460_;
 wire _22461_;
 wire _22462_;
 wire _22463_;
 wire _22464_;
 wire _22465_;
 wire _22466_;
 wire _22467_;
 wire _22468_;
 wire _22469_;
 wire _22470_;
 wire _22471_;
 wire _22472_;
 wire _22473_;
 wire _22474_;
 wire _22475_;
 wire _22476_;
 wire _22477_;
 wire _22478_;
 wire _22479_;
 wire _22480_;
 wire _22481_;
 wire _22482_;
 wire _22483_;
 wire _22484_;
 wire _22485_;
 wire _22486_;
 wire _22487_;
 wire _22488_;
 wire _22489_;
 wire _22490_;
 wire _22491_;
 wire _22492_;
 wire _22493_;
 wire _22494_;
 wire _22495_;
 wire _22496_;
 wire _22497_;
 wire _22498_;
 wire _22499_;
 wire _22500_;
 wire _22501_;
 wire _22502_;
 wire _22503_;
 wire _22504_;
 wire _22505_;
 wire _22506_;
 wire _22507_;
 wire _22508_;
 wire _22509_;
 wire _22510_;
 wire _22511_;
 wire _22512_;
 wire _22513_;
 wire _22514_;
 wire _22515_;
 wire _22516_;
 wire _22517_;
 wire _22518_;
 wire _22519_;
 wire _22520_;
 wire _22521_;
 wire _22522_;
 wire _22523_;
 wire _22524_;
 wire _22525_;
 wire _22526_;
 wire _22527_;
 wire _22528_;
 wire _22529_;
 wire _22530_;
 wire _22531_;
 wire _22532_;
 wire _22533_;
 wire _22534_;
 wire _22535_;
 wire _22536_;
 wire _22537_;
 wire _22538_;
 wire _22539_;
 wire _22540_;
 wire _22541_;
 wire _22542_;
 wire _22543_;
 wire _22544_;
 wire _22545_;
 wire _22546_;
 wire _22547_;
 wire _22548_;
 wire _22549_;
 wire _22550_;
 wire _22551_;
 wire _22552_;
 wire _22553_;
 wire _22554_;
 wire _22555_;
 wire _22556_;
 wire _22557_;
 wire _22558_;
 wire _22559_;
 wire _22560_;
 wire _22561_;
 wire _22562_;
 wire _22563_;
 wire _22564_;
 wire _22565_;
 wire _22566_;
 wire _22567_;
 wire _22568_;
 wire _22569_;
 wire _22570_;
 wire _22571_;
 wire _22572_;
 wire _22573_;
 wire _22574_;
 wire _22575_;
 wire _22576_;
 wire _22577_;
 wire _22578_;
 wire _22579_;
 wire _22580_;
 wire _22581_;
 wire _22582_;
 wire _22583_;
 wire _22584_;
 wire _22585_;
 wire _22586_;
 wire _22587_;
 wire _22588_;
 wire _22589_;
 wire _22590_;
 wire _22591_;
 wire _22592_;
 wire _22593_;
 wire _22594_;
 wire _22595_;
 wire _22596_;
 wire _22597_;
 wire _22598_;
 wire _22599_;
 wire _22600_;
 wire _22601_;
 wire _22602_;
 wire _22603_;
 wire _22604_;
 wire _22605_;
 wire _22606_;
 wire _22607_;
 wire _22608_;
 wire _22609_;
 wire _22610_;
 wire _22611_;
 wire _22612_;
 wire _22613_;
 wire _22614_;
 wire _22615_;
 wire _22616_;
 wire _22617_;
 wire _22618_;
 wire _22619_;
 wire _22620_;
 wire _22621_;
 wire _22622_;
 wire _22623_;
 wire _22624_;
 wire _22625_;
 wire _22626_;
 wire _22627_;
 wire _22628_;
 wire _22629_;
 wire _22630_;
 wire _22631_;
 wire _22632_;
 wire _22633_;
 wire _22634_;
 wire _22635_;
 wire _22636_;
 wire _22637_;
 wire _22638_;
 wire _22639_;
 wire _22640_;
 wire _22641_;
 wire _22642_;
 wire _22643_;
 wire _22644_;
 wire _22645_;
 wire _22646_;
 wire _22647_;
 wire _22648_;
 wire _22649_;
 wire _22650_;
 wire _22651_;
 wire _22652_;
 wire _22653_;
 wire _22654_;
 wire _22655_;
 wire _22656_;
 wire _22657_;
 wire _22658_;
 wire _22659_;
 wire _22660_;
 wire _22661_;
 wire _22662_;
 wire _22663_;
 wire _22664_;
 wire _22665_;
 wire _22666_;
 wire _22667_;
 wire _22668_;
 wire _22669_;
 wire _22670_;
 wire _22671_;
 wire _22672_;
 wire _22673_;
 wire _22674_;
 wire _22675_;
 wire _22676_;
 wire _22677_;
 wire _22678_;
 wire _22679_;
 wire _22680_;
 wire _22681_;
 wire _22682_;
 wire _22683_;
 wire _22684_;
 wire _22685_;
 wire _22686_;
 wire _22687_;
 wire _22688_;
 wire _22689_;
 wire _22690_;
 wire _22691_;
 wire _22692_;
 wire _22693_;
 wire _22694_;
 wire _22695_;
 wire _22696_;
 wire _22697_;
 wire _22698_;
 wire _22699_;
 wire _22700_;
 wire _22701_;
 wire _22702_;
 wire _22703_;
 wire _22704_;
 wire _22705_;
 wire _22706_;
 wire _22707_;
 wire _22708_;
 wire _22709_;
 wire _22710_;
 wire _22711_;
 wire _22712_;
 wire _22713_;
 wire _22714_;
 wire _22715_;
 wire _22716_;
 wire _22717_;
 wire _22718_;
 wire _22719_;
 wire _22720_;
 wire _22721_;
 wire _22722_;
 wire _22723_;
 wire _22724_;
 wire _22725_;
 wire _22726_;
 wire _22727_;
 wire _22728_;
 wire _22729_;
 wire _22730_;
 wire _22731_;
 wire _22732_;
 wire _22733_;
 wire _22734_;
 wire _22735_;
 wire _22736_;
 wire _22737_;
 wire _22738_;
 wire _22739_;
 wire _22740_;
 wire _22741_;
 wire _22742_;
 wire _22743_;
 wire _22744_;
 wire _22745_;
 wire _22746_;
 wire _22747_;
 wire _22748_;
 wire _22749_;
 wire _22750_;
 wire _22751_;
 wire _22752_;
 wire _22753_;
 wire _22754_;
 wire _22755_;
 wire _22756_;
 wire _22757_;
 wire _22758_;
 wire _22759_;
 wire _22760_;
 wire _22761_;
 wire _22762_;
 wire _22763_;
 wire _22764_;
 wire _22765_;
 wire _22766_;
 wire _22767_;
 wire _22768_;
 wire _22769_;
 wire _22770_;
 wire _22771_;
 wire _22772_;
 wire _22773_;
 wire _22774_;
 wire _22775_;
 wire _22776_;
 wire _22777_;
 wire _22778_;
 wire _22779_;
 wire _22780_;
 wire _22781_;
 wire _22782_;
 wire _22783_;
 wire _22784_;
 wire _22785_;
 wire _22786_;
 wire _22787_;
 wire _22788_;
 wire _22789_;
 wire _22790_;
 wire _22791_;
 wire _22792_;
 wire _22793_;
 wire _22794_;
 wire _22795_;
 wire _22796_;
 wire _22797_;
 wire _22798_;
 wire _22799_;
 wire _22800_;
 wire _22801_;
 wire _22802_;
 wire _22803_;
 wire _22804_;
 wire _22805_;
 wire _22806_;
 wire _22807_;
 wire _22808_;
 wire _22809_;
 wire _22810_;
 wire _22811_;
 wire _22812_;
 wire _22813_;
 wire _22814_;
 wire _22815_;
 wire _22816_;
 wire _22817_;
 wire _22818_;
 wire _22819_;
 wire _22820_;
 wire _22821_;
 wire _22822_;
 wire _22823_;
 wire _22824_;
 wire _22825_;
 wire _22826_;
 wire _22827_;
 wire _22828_;
 wire _22829_;
 wire _22830_;
 wire _22831_;
 wire _22832_;
 wire _22833_;
 wire _22834_;
 wire _22835_;
 wire _22836_;
 wire _22837_;
 wire _22838_;
 wire _22839_;
 wire _22840_;
 wire _22841_;
 wire _22842_;
 wire _22843_;
 wire _22844_;
 wire _22845_;
 wire _22846_;
 wire _22847_;
 wire _22848_;
 wire _22849_;
 wire _22850_;
 wire _22851_;
 wire _22852_;
 wire _22853_;
 wire _22854_;
 wire _22855_;
 wire _22856_;
 wire _22857_;
 wire _22858_;
 wire _22859_;
 wire _22860_;
 wire _22861_;
 wire _22862_;
 wire _22863_;
 wire _22864_;
 wire _22865_;
 wire _22866_;
 wire _22867_;
 wire _22868_;
 wire _22869_;
 wire _22870_;
 wire _22871_;
 wire _22872_;
 wire _22873_;
 wire _22874_;
 wire _22875_;
 wire _22876_;
 wire _22877_;
 wire _22878_;
 wire _22879_;
 wire _22880_;
 wire _22881_;
 wire _22882_;
 wire _22883_;
 wire _22884_;
 wire _22885_;
 wire _22886_;
 wire _22887_;
 wire _22888_;
 wire _22889_;
 wire _22890_;
 wire _22891_;
 wire _22892_;
 wire _22893_;
 wire _22894_;
 wire _22895_;
 wire _22896_;
 wire _22897_;
 wire _22898_;
 wire _22899_;
 wire _22900_;
 wire _22901_;
 wire _22902_;
 wire _22903_;
 wire _22904_;
 wire _22905_;
 wire _22906_;
 wire _22907_;
 wire _22908_;
 wire _22909_;
 wire _22910_;
 wire _22911_;
 wire _22912_;
 wire _22913_;
 wire _22914_;
 wire _22915_;
 wire _22916_;
 wire _22917_;
 wire _22918_;
 wire _22919_;
 wire _22920_;
 wire _22921_;
 wire _22922_;
 wire _22923_;
 wire _22924_;
 wire _22925_;
 wire _22926_;
 wire _22927_;
 wire _22928_;
 wire _22929_;
 wire _22930_;
 wire _22931_;
 wire _22932_;
 wire _22933_;
 wire _22934_;
 wire _22935_;
 wire _22936_;
 wire _22937_;
 wire _22938_;
 wire _22939_;
 wire _22940_;
 wire _22941_;
 wire _22942_;
 wire _22943_;
 wire _22944_;
 wire _22945_;
 wire _22946_;
 wire _22947_;
 wire _22948_;
 wire _22949_;
 wire _22950_;
 wire _22951_;
 wire _22952_;
 wire _22953_;
 wire _22954_;
 wire _22955_;
 wire _22956_;
 wire _22957_;
 wire _22958_;
 wire _22959_;
 wire _22960_;
 wire _22961_;
 wire _22962_;
 wire _22963_;
 wire _22964_;
 wire _22965_;
 wire _22966_;
 wire _22967_;
 wire _22968_;
 wire _22969_;
 wire _22970_;
 wire _22971_;
 wire _22972_;
 wire _22973_;
 wire _22974_;
 wire _22975_;
 wire _22976_;
 wire _22977_;
 wire _22978_;
 wire _22979_;
 wire _22980_;
 wire _22981_;
 wire _22982_;
 wire _22983_;
 wire _22984_;
 wire _22985_;
 wire _22986_;
 wire _22987_;
 wire _22988_;
 wire _22989_;
 wire _22990_;
 wire _22991_;
 wire _22992_;
 wire _22993_;
 wire _22994_;
 wire _22995_;
 wire _22996_;
 wire _22997_;
 wire _22998_;
 wire _22999_;
 wire _23000_;
 wire _23001_;
 wire _23002_;
 wire _23003_;
 wire _23004_;
 wire _23005_;
 wire _23006_;
 wire _23007_;
 wire _23008_;
 wire _23009_;
 wire _23010_;
 wire _23011_;
 wire _23012_;
 wire _23013_;
 wire _23014_;
 wire _23015_;
 wire _23016_;
 wire _23017_;
 wire _23018_;
 wire _23019_;
 wire _23020_;
 wire _23021_;
 wire _23022_;
 wire _23023_;
 wire _23024_;
 wire _23025_;
 wire _23026_;
 wire _23027_;
 wire _23028_;
 wire _23029_;
 wire _23030_;
 wire _23031_;
 wire _23032_;
 wire _23033_;
 wire _23034_;
 wire _23035_;
 wire _23036_;
 wire _23037_;
 wire _23038_;
 wire _23039_;
 wire _23040_;
 wire _23041_;
 wire _23042_;
 wire _23043_;
 wire _23044_;
 wire _23045_;
 wire _23046_;
 wire _23047_;
 wire _23048_;
 wire _23049_;
 wire _23050_;
 wire _23051_;
 wire _23052_;
 wire _23053_;
 wire _23054_;
 wire _23055_;
 wire _23056_;
 wire _23057_;
 wire _23058_;
 wire _23059_;
 wire _23060_;
 wire _23061_;
 wire _23062_;
 wire _23063_;
 wire _23064_;
 wire _23065_;
 wire _23066_;
 wire _23067_;
 wire _23068_;
 wire _23069_;
 wire _23070_;
 wire _23071_;
 wire _23072_;
 wire _23073_;
 wire _23074_;
 wire _23075_;
 wire _23076_;
 wire _23077_;
 wire _23078_;
 wire _23079_;
 wire _23080_;
 wire _23081_;
 wire _23082_;
 wire _23083_;
 wire _23084_;
 wire _23085_;
 wire _23086_;
 wire _23087_;
 wire _23088_;
 wire _23089_;
 wire _23090_;
 wire _23091_;
 wire _23092_;
 wire _23093_;
 wire _23094_;
 wire _23095_;
 wire _23096_;
 wire _23097_;
 wire _23098_;
 wire _23099_;
 wire _23100_;
 wire _23101_;
 wire _23102_;
 wire _23103_;
 wire _23104_;
 wire _23105_;
 wire _23106_;
 wire _23107_;
 wire _23108_;
 wire _23109_;
 wire _23110_;
 wire _23111_;
 wire _23112_;
 wire _23113_;
 wire _23114_;
 wire _23115_;
 wire _23116_;
 wire _23117_;
 wire _23118_;
 wire _23119_;
 wire _23120_;
 wire _23121_;
 wire _23122_;
 wire _23123_;
 wire _23124_;
 wire _23125_;
 wire _23126_;
 wire _23127_;
 wire _23128_;
 wire _23129_;
 wire _23130_;
 wire _23131_;
 wire _23132_;
 wire _23133_;
 wire _23134_;
 wire _23135_;
 wire _23136_;
 wire _23137_;
 wire _23138_;
 wire _23139_;
 wire _23140_;
 wire _23141_;
 wire _23142_;
 wire _23143_;
 wire _23144_;
 wire _23145_;
 wire _23146_;
 wire _23147_;
 wire _23148_;
 wire _23149_;
 wire _23150_;
 wire _23151_;
 wire _23152_;
 wire _23153_;
 wire _23154_;
 wire _23155_;
 wire _23156_;
 wire _23157_;
 wire _23158_;
 wire _23159_;
 wire _23160_;
 wire _23161_;
 wire _23162_;
 wire _23163_;
 wire _23164_;
 wire _23165_;
 wire _23166_;
 wire _23167_;
 wire _23168_;
 wire _23169_;
 wire _23170_;
 wire _23171_;
 wire _23172_;
 wire _23173_;
 wire _23174_;
 wire _23175_;
 wire _23176_;
 wire _23177_;
 wire _23178_;
 wire _23179_;
 wire _23180_;
 wire _23181_;
 wire _23182_;
 wire _23183_;
 wire _23184_;
 wire _23185_;
 wire _23186_;
 wire _23187_;
 wire _23188_;
 wire _23189_;
 wire _23190_;
 wire _23191_;
 wire _23192_;
 wire _23193_;
 wire _23194_;
 wire _23195_;
 wire _23196_;
 wire _23197_;
 wire _23198_;
 wire _23199_;
 wire _23200_;
 wire _23201_;
 wire _23202_;
 wire _23203_;
 wire _23204_;
 wire _23205_;
 wire _23206_;
 wire _23207_;
 wire _23208_;
 wire _23209_;
 wire _23210_;
 wire _23211_;
 wire _23212_;
 wire _23213_;
 wire _23214_;
 wire _23215_;
 wire _23216_;
 wire _23217_;
 wire _23218_;
 wire _23219_;
 wire _23220_;
 wire _23221_;
 wire _23222_;
 wire _23223_;
 wire _23224_;
 wire _23225_;
 wire _23226_;
 wire _23227_;
 wire _23228_;
 wire _23229_;
 wire _23230_;
 wire _23231_;
 wire _23232_;
 wire _23233_;
 wire _23234_;
 wire _23235_;
 wire _23236_;
 wire _23237_;
 wire _23238_;
 wire _23239_;
 wire _23240_;
 wire _23241_;
 wire _23242_;
 wire _23243_;
 wire _23244_;
 wire _23245_;
 wire _23246_;
 wire _23247_;
 wire _23248_;
 wire _23249_;
 wire _23250_;
 wire _23251_;
 wire _23252_;
 wire _23253_;
 wire _23254_;
 wire _23255_;
 wire _23256_;
 wire _23257_;
 wire _23258_;
 wire _23259_;
 wire _23260_;
 wire _23261_;
 wire _23262_;
 wire _23263_;
 wire _23264_;
 wire _23265_;
 wire _23266_;
 wire _23267_;
 wire _23268_;
 wire _23269_;
 wire _23270_;
 wire _23271_;
 wire _23272_;
 wire _23273_;
 wire _23274_;
 wire _23275_;
 wire _23276_;
 wire _23277_;
 wire _23278_;
 wire _23279_;
 wire _23280_;
 wire _23281_;
 wire _23282_;
 wire _23283_;
 wire _23284_;
 wire _23285_;
 wire _23286_;
 wire _23287_;
 wire _23288_;
 wire _23289_;
 wire _23290_;
 wire _23291_;
 wire _23292_;
 wire _23293_;
 wire _23294_;
 wire _23295_;
 wire _23296_;
 wire _23297_;
 wire _23298_;
 wire _23299_;
 wire _23300_;
 wire _23301_;
 wire _23302_;
 wire _23303_;
 wire _23304_;
 wire _23305_;
 wire _23306_;
 wire _23307_;
 wire _23308_;
 wire _23309_;
 wire _23310_;
 wire _23311_;
 wire _23312_;
 wire _23313_;
 wire _23314_;
 wire _23315_;
 wire _23316_;
 wire _23317_;
 wire _23318_;
 wire _23319_;
 wire _23320_;
 wire _23321_;
 wire _23322_;
 wire _23323_;
 wire _23324_;
 wire _23325_;
 wire _23326_;
 wire _23327_;
 wire _23328_;
 wire _23329_;
 wire _23330_;
 wire _23331_;
 wire _23332_;
 wire _23333_;
 wire _23334_;
 wire _23335_;
 wire _23336_;
 wire _23337_;
 wire _23338_;
 wire _23339_;
 wire _23340_;
 wire _23341_;
 wire _23342_;
 wire _23343_;
 wire _23344_;
 wire _23345_;
 wire _23346_;
 wire _23347_;
 wire _23348_;
 wire _23349_;
 wire _23350_;
 wire _23351_;
 wire _23352_;
 wire _23353_;
 wire _23354_;
 wire _23355_;
 wire _23356_;
 wire _23357_;
 wire _23358_;
 wire _23359_;
 wire _23360_;
 wire _23361_;
 wire _23362_;
 wire _23363_;
 wire _23364_;
 wire _23365_;
 wire _23366_;
 wire _23367_;
 wire _23368_;
 wire _23369_;
 wire _23370_;
 wire _23371_;
 wire _23372_;
 wire _23373_;
 wire _23374_;
 wire _23375_;
 wire _23376_;
 wire _23377_;
 wire _23378_;
 wire _23379_;
 wire _23380_;
 wire _23381_;
 wire _23382_;
 wire _23383_;
 wire _23384_;
 wire _23385_;
 wire _23386_;
 wire _23387_;
 wire _23388_;
 wire _23389_;
 wire _23390_;
 wire _23391_;
 wire _23392_;
 wire _23393_;
 wire _23394_;
 wire _23395_;
 wire _23396_;
 wire _23397_;
 wire _23398_;
 wire _23399_;
 wire _23400_;
 wire _23401_;
 wire _23402_;
 wire _23403_;
 wire _23404_;
 wire _23405_;
 wire _23406_;
 wire _23407_;
 wire _23408_;
 wire _23409_;
 wire _23410_;
 wire _23411_;
 wire _23412_;
 wire _23413_;
 wire _23414_;
 wire _23415_;
 wire _23416_;
 wire _23417_;
 wire _23418_;
 wire _23419_;
 wire _23420_;
 wire _23421_;
 wire _23422_;
 wire _23423_;
 wire _23424_;
 wire _23425_;
 wire _23426_;
 wire _23427_;
 wire _23428_;
 wire _23429_;
 wire _23430_;
 wire _23431_;
 wire _23432_;
 wire _23433_;
 wire _23434_;
 wire _23435_;
 wire _23436_;
 wire _23437_;
 wire _23438_;
 wire _23439_;
 wire _23440_;
 wire _23441_;
 wire _23442_;
 wire _23443_;
 wire _23444_;
 wire _23445_;
 wire _23446_;
 wire _23447_;
 wire _23448_;
 wire _23449_;
 wire _23450_;
 wire _23451_;
 wire _23452_;
 wire _23453_;
 wire _23454_;
 wire _23455_;
 wire _23456_;
 wire _23457_;
 wire _23458_;
 wire _23459_;
 wire _23460_;
 wire _23461_;
 wire _23462_;
 wire _23463_;
 wire _23464_;
 wire _23465_;
 wire _23466_;
 wire _23467_;
 wire _23468_;
 wire _23469_;
 wire _23470_;
 wire _23471_;
 wire _23472_;
 wire _23473_;
 wire _23474_;
 wire _23475_;
 wire _23476_;
 wire _23477_;
 wire _23478_;
 wire _23479_;
 wire _23480_;
 wire _23481_;
 wire _23482_;
 wire _23483_;
 wire _23484_;
 wire _23485_;
 wire _23486_;
 wire _23487_;
 wire _23488_;
 wire _23489_;
 wire _23490_;
 wire _23491_;
 wire _23492_;
 wire _23493_;
 wire _23494_;
 wire _23495_;
 wire _23496_;
 wire _23497_;
 wire _23498_;
 wire _23499_;
 wire _23500_;
 wire _23501_;
 wire _23502_;
 wire _23503_;
 wire _23504_;
 wire _23505_;
 wire _23506_;
 wire _23507_;
 wire _23508_;
 wire _23509_;
 wire _23510_;
 wire _23511_;
 wire _23512_;
 wire _23513_;
 wire _23514_;
 wire _23515_;
 wire _23516_;
 wire _23517_;
 wire _23518_;
 wire _23519_;
 wire _23520_;
 wire _23521_;
 wire _23522_;
 wire _23523_;
 wire _23524_;
 wire _23525_;
 wire _23526_;
 wire _23527_;
 wire _23528_;
 wire _23529_;
 wire _23530_;
 wire _23531_;
 wire _23532_;
 wire _23533_;
 wire _23534_;
 wire _23535_;
 wire _23536_;
 wire _23537_;
 wire _23538_;
 wire _23539_;
 wire _23540_;
 wire _23541_;
 wire _23542_;
 wire _23543_;
 wire _23544_;
 wire _23545_;
 wire _23546_;
 wire _23547_;
 wire _23548_;
 wire _23549_;
 wire _23550_;
 wire _23551_;
 wire _23552_;
 wire _23553_;
 wire _23554_;
 wire _23555_;
 wire _23556_;
 wire _23557_;
 wire _23558_;
 wire _23559_;
 wire _23560_;
 wire _23561_;
 wire _23562_;
 wire _23563_;
 wire _23564_;
 wire _23565_;
 wire _23566_;
 wire _23567_;
 wire _23568_;
 wire _23569_;
 wire _23570_;
 wire _23571_;
 wire _23572_;
 wire _23573_;
 wire _23574_;
 wire _23575_;
 wire _23576_;
 wire _23577_;
 wire _23578_;
 wire _23579_;
 wire _23580_;
 wire _23581_;
 wire _23582_;
 wire _23583_;
 wire _23584_;
 wire _23585_;
 wire _23586_;
 wire _23587_;
 wire _23588_;
 wire _23589_;
 wire _23590_;
 wire _23591_;
 wire _23592_;
 wire _23593_;
 wire _23594_;
 wire _23595_;
 wire _23596_;
 wire _23597_;
 wire _23598_;
 wire _23599_;
 wire _23600_;
 wire _23601_;
 wire _23602_;
 wire _23603_;
 wire _23604_;
 wire _23605_;
 wire _23606_;
 wire _23607_;
 wire _23608_;
 wire _23609_;
 wire _23610_;
 wire _23611_;
 wire _23612_;
 wire _23613_;
 wire _23614_;
 wire _23615_;
 wire _23616_;
 wire _23617_;
 wire _23618_;
 wire _23619_;
 wire _23620_;
 wire _23621_;
 wire _23622_;
 wire _23623_;
 wire _23624_;
 wire _23625_;
 wire _23626_;
 wire _23627_;
 wire _23628_;
 wire _23629_;
 wire _23630_;
 wire _23631_;
 wire _23632_;
 wire _23633_;
 wire _23634_;
 wire _23635_;
 wire _23636_;
 wire _23637_;
 wire _23638_;
 wire _23639_;
 wire _23640_;
 wire _23641_;
 wire _23642_;
 wire _23643_;
 wire _23644_;
 wire _23645_;
 wire _23646_;
 wire _23647_;
 wire _23648_;
 wire _23649_;
 wire _23650_;
 wire _23651_;
 wire _23652_;
 wire _23653_;
 wire _23654_;
 wire _23655_;
 wire _23656_;
 wire _23657_;
 wire _23658_;
 wire _23659_;
 wire _23660_;
 wire _23661_;
 wire _23662_;
 wire _23663_;
 wire _23664_;
 wire _23665_;
 wire _23666_;
 wire _23667_;
 wire _23668_;
 wire _23669_;
 wire _23670_;
 wire _23671_;
 wire _23672_;
 wire _23673_;
 wire _23674_;
 wire _23675_;
 wire _23676_;
 wire _23677_;
 wire _23678_;
 wire _23679_;
 wire _23680_;
 wire _23681_;
 wire _23682_;
 wire _23683_;
 wire _23684_;
 wire _23685_;
 wire _23686_;
 wire _23687_;
 wire _23688_;
 wire _23689_;
 wire _23690_;
 wire _23691_;
 wire _23692_;
 wire _23693_;
 wire _23694_;
 wire _23695_;
 wire _23696_;
 wire _23697_;
 wire _23698_;
 wire _23699_;
 wire _23700_;
 wire _23701_;
 wire _23702_;
 wire _23703_;
 wire _23704_;
 wire _23705_;
 wire _23706_;
 wire _23707_;
 wire _23708_;
 wire _23709_;
 wire _23710_;
 wire _23711_;
 wire _23712_;
 wire _23713_;
 wire _23714_;
 wire _23715_;
 wire _23716_;
 wire _23717_;
 wire _23718_;
 wire _23719_;
 wire _23720_;
 wire _23721_;
 wire _23722_;
 wire _23723_;
 wire _23724_;
 wire _23725_;
 wire _23726_;
 wire _23727_;
 wire _23728_;
 wire _23729_;
 wire _23730_;
 wire _23731_;
 wire _23732_;
 wire _23733_;
 wire _23734_;
 wire _23735_;
 wire _23736_;
 wire _23737_;
 wire _23738_;
 wire _23739_;
 wire _23740_;
 wire _23741_;
 wire _23742_;
 wire _23743_;
 wire _23744_;
 wire _23745_;
 wire _23746_;
 wire _23747_;
 wire _23748_;
 wire _23749_;
 wire _23750_;
 wire _23751_;
 wire _23752_;
 wire _23753_;
 wire _23754_;
 wire _23755_;
 wire _23756_;
 wire _23757_;
 wire _23758_;
 wire _23759_;
 wire _23760_;
 wire _23761_;
 wire _23762_;
 wire _23763_;
 wire _23764_;
 wire _23765_;
 wire _23766_;
 wire _23767_;
 wire _23768_;
 wire _23769_;
 wire _23770_;
 wire _23771_;
 wire _23772_;
 wire _23773_;
 wire _23774_;
 wire _23775_;
 wire _23776_;
 wire _23777_;
 wire _23778_;
 wire _23779_;
 wire _23780_;
 wire _23781_;
 wire _23782_;
 wire _23783_;
 wire _23784_;
 wire _23785_;
 wire _23786_;
 wire _23787_;
 wire _23788_;
 wire _23789_;
 wire _23790_;
 wire _23791_;
 wire _23792_;
 wire _23793_;
 wire _23794_;
 wire _23795_;
 wire _23796_;
 wire _23797_;
 wire _23798_;
 wire _23799_;
 wire _23800_;
 wire _23801_;
 wire _23802_;
 wire _23803_;
 wire _23804_;
 wire _23805_;
 wire _23806_;
 wire _23807_;
 wire _23808_;
 wire _23809_;
 wire _23810_;
 wire _23811_;
 wire _23812_;
 wire _23813_;
 wire _23814_;
 wire _23815_;
 wire _23816_;
 wire _23817_;
 wire _23818_;
 wire _23819_;
 wire _23820_;
 wire _23821_;
 wire _23822_;
 wire _23823_;
 wire _23824_;
 wire _23825_;
 wire _23826_;
 wire _23827_;
 wire _23828_;
 wire _23829_;
 wire _23830_;
 wire _23831_;
 wire _23832_;
 wire _23833_;
 wire _23834_;
 wire _23835_;
 wire _23836_;
 wire _23837_;
 wire _23838_;
 wire _23839_;
 wire _23840_;
 wire _23841_;
 wire _23842_;
 wire _23843_;
 wire _23844_;
 wire _23845_;
 wire _23846_;
 wire _23847_;
 wire _23848_;
 wire _23849_;
 wire _23850_;
 wire _23851_;
 wire _23852_;
 wire _23853_;
 wire _23854_;
 wire _23855_;
 wire _23856_;
 wire _23857_;
 wire _23858_;
 wire _23859_;
 wire _23860_;
 wire _23861_;
 wire _23862_;
 wire _23863_;
 wire _23864_;
 wire _23865_;
 wire _23866_;
 wire _23867_;
 wire _23868_;
 wire _23869_;
 wire _23870_;
 wire _23871_;
 wire _23872_;
 wire _23873_;
 wire _23874_;
 wire _23875_;
 wire _23876_;
 wire _23877_;
 wire _23878_;
 wire _23879_;
 wire _23880_;
 wire _23881_;
 wire _23882_;
 wire _23883_;
 wire _23884_;
 wire _23885_;
 wire _23886_;
 wire _23887_;
 wire _23888_;
 wire _23889_;
 wire _23890_;
 wire _23891_;
 wire _23892_;
 wire _23893_;
 wire _23894_;
 wire _23895_;
 wire _23896_;
 wire _23897_;
 wire _23898_;
 wire _23899_;
 wire _23900_;
 wire _23901_;
 wire _23902_;
 wire _23903_;
 wire _23904_;
 wire _23905_;
 wire _23906_;
 wire _23907_;
 wire _23908_;
 wire _23909_;
 wire _23910_;
 wire _23911_;
 wire _23912_;
 wire _23913_;
 wire _23914_;
 wire _23915_;
 wire _23916_;
 wire _23917_;
 wire _23918_;
 wire _23919_;
 wire _23920_;
 wire _23921_;
 wire _23922_;
 wire _23923_;
 wire _23924_;
 wire _23925_;
 wire _23926_;
 wire _23927_;
 wire _23928_;
 wire _23929_;
 wire _23930_;
 wire _23931_;
 wire _23932_;
 wire _23933_;
 wire _23934_;
 wire _23935_;
 wire _23936_;
 wire _23937_;
 wire _23938_;
 wire _23939_;
 wire _23940_;
 wire _23941_;
 wire _23942_;
 wire _23943_;
 wire _23944_;
 wire _23945_;
 wire _23946_;
 wire _23947_;
 wire _23948_;
 wire _23949_;
 wire _23950_;
 wire _23951_;
 wire _23952_;
 wire _23953_;
 wire _23954_;
 wire _23955_;
 wire _23956_;
 wire _23957_;
 wire _23958_;
 wire _23959_;
 wire _23960_;
 wire _23961_;
 wire _23962_;
 wire _23963_;
 wire _23964_;
 wire _23965_;
 wire _23966_;
 wire _23967_;
 wire _23968_;
 wire _23969_;
 wire _23970_;
 wire _23971_;
 wire _23972_;
 wire _23973_;
 wire _23974_;
 wire _23975_;
 wire _23976_;
 wire _23977_;
 wire _23978_;
 wire _23979_;
 wire _23980_;
 wire _23981_;
 wire _23982_;
 wire _23983_;
 wire _23984_;
 wire _23985_;
 wire _23986_;
 wire _23987_;
 wire _23988_;
 wire _23989_;
 wire _23990_;
 wire _23991_;
 wire _23992_;
 wire _23993_;
 wire _23994_;
 wire _23995_;
 wire _23996_;
 wire _23997_;
 wire _23998_;
 wire _23999_;
 wire _24000_;
 wire _24001_;
 wire _24002_;
 wire _24003_;
 wire _24004_;
 wire _24005_;
 wire _24006_;
 wire _24007_;
 wire _24008_;
 wire _24009_;
 wire _24010_;
 wire _24011_;
 wire _24012_;
 wire _24013_;
 wire _24014_;
 wire _24015_;
 wire _24016_;
 wire _24017_;
 wire _24018_;
 wire _24019_;
 wire _24020_;
 wire _24021_;
 wire _24022_;
 wire _24023_;
 wire _24024_;
 wire _24025_;
 wire _24026_;
 wire _24027_;
 wire _24028_;
 wire _24029_;
 wire _24030_;
 wire _24031_;
 wire _24032_;
 wire _24033_;
 wire _24034_;
 wire _24035_;
 wire _24036_;
 wire _24037_;
 wire _24038_;
 wire _24039_;
 wire _24040_;
 wire _24041_;
 wire _24042_;
 wire _24043_;
 wire _24044_;
 wire _24045_;
 wire _24046_;
 wire _24047_;
 wire _24048_;
 wire _24049_;
 wire _24050_;
 wire _24051_;
 wire _24052_;
 wire _24053_;
 wire _24054_;
 wire _24055_;
 wire _24056_;
 wire _24057_;
 wire _24058_;
 wire _24059_;
 wire _24060_;
 wire _24061_;
 wire _24062_;
 wire _24063_;
 wire _24064_;
 wire _24065_;
 wire _24066_;
 wire _24067_;
 wire _24068_;
 wire _24069_;
 wire _24070_;
 wire _24071_;
 wire _24072_;
 wire _24073_;
 wire _24074_;
 wire _24075_;
 wire _24076_;
 wire _24077_;
 wire _24078_;
 wire _24079_;
 wire _24080_;
 wire _24081_;
 wire _24082_;
 wire _24083_;
 wire _24084_;
 wire _24085_;
 wire _24086_;
 wire _24087_;
 wire _24088_;
 wire _24089_;
 wire _24090_;
 wire _24091_;
 wire _24092_;
 wire _24093_;
 wire _24094_;
 wire _24095_;
 wire _24096_;
 wire _24097_;
 wire _24098_;
 wire _24099_;
 wire _24100_;
 wire _24101_;
 wire _24102_;
 wire _24103_;
 wire _24104_;
 wire _24105_;
 wire _24106_;
 wire _24107_;
 wire _24108_;
 wire _24109_;
 wire _24110_;
 wire _24111_;
 wire _24112_;
 wire _24113_;
 wire _24114_;
 wire _24115_;
 wire _24116_;
 wire _24117_;
 wire _24118_;
 wire _24119_;
 wire _24120_;
 wire _24121_;
 wire _24122_;
 wire _24123_;
 wire _24124_;
 wire _24125_;
 wire _24126_;
 wire _24127_;
 wire _24128_;
 wire _24129_;
 wire _24130_;
 wire _24131_;
 wire _24132_;
 wire _24133_;
 wire _24134_;
 wire _24135_;
 wire _24136_;
 wire _24137_;
 wire _24138_;
 wire _24139_;
 wire _24140_;
 wire _24141_;
 wire _24142_;
 wire _24143_;
 wire _24144_;
 wire _24145_;
 wire _24146_;
 wire _24147_;
 wire _24148_;
 wire _24149_;
 wire _24150_;
 wire _24151_;
 wire _24152_;
 wire _24153_;
 wire _24154_;
 wire _24155_;
 wire _24156_;
 wire _24157_;
 wire _24158_;
 wire _24159_;
 wire _24160_;
 wire _24161_;
 wire _24162_;
 wire _24163_;
 wire _24164_;
 wire _24165_;
 wire _24166_;
 wire _24167_;
 wire _24168_;
 wire _24169_;
 wire _24170_;
 wire _24171_;
 wire _24172_;
 wire _24173_;
 wire _24174_;
 wire _24175_;
 wire _24176_;
 wire _24177_;
 wire _24178_;
 wire _24179_;
 wire _24180_;
 wire _24181_;
 wire _24182_;
 wire _24183_;
 wire _24184_;
 wire _24185_;
 wire _24186_;
 wire _24187_;
 wire _24188_;
 wire _24189_;
 wire _24190_;
 wire _24191_;
 wire _24192_;
 wire _24193_;
 wire _24194_;
 wire _24195_;
 wire _24196_;
 wire _24197_;
 wire _24198_;
 wire _24199_;
 wire _24200_;
 wire _24201_;
 wire _24202_;
 wire _24203_;
 wire _24204_;
 wire _24205_;
 wire _24206_;
 wire _24207_;
 wire _24208_;
 wire _24209_;
 wire _24210_;
 wire _24211_;
 wire _24212_;
 wire _24213_;
 wire _24214_;
 wire _24215_;
 wire _24216_;
 wire _24217_;
 wire _24218_;
 wire _24219_;
 wire _24220_;
 wire _24221_;
 wire _24222_;
 wire _24223_;
 wire _24224_;
 wire _24225_;
 wire _24226_;
 wire _24227_;
 wire _24228_;
 wire _24229_;
 wire _24230_;
 wire _24231_;
 wire _24232_;
 wire _24233_;
 wire _24234_;
 wire _24235_;
 wire _24236_;
 wire _24237_;
 wire _24238_;
 wire _24239_;
 wire _24240_;
 wire _24241_;
 wire _24242_;
 wire _24243_;
 wire _24244_;
 wire _24245_;
 wire _24246_;
 wire _24247_;
 wire _24248_;
 wire _24249_;
 wire _24250_;
 wire _24251_;
 wire _24252_;
 wire _24253_;
 wire _24254_;
 wire _24255_;
 wire _24256_;
 wire _24257_;
 wire _24258_;
 wire _24259_;
 wire _24260_;
 wire _24261_;
 wire _24262_;
 wire _24263_;
 wire _24264_;
 wire _24265_;
 wire _24266_;
 wire _24267_;
 wire _24268_;
 wire _24269_;
 wire _24270_;
 wire _24271_;
 wire _24272_;
 wire _24273_;
 wire _24274_;
 wire _24275_;
 wire _24276_;
 wire _24277_;
 wire _24278_;
 wire _24279_;
 wire _24280_;
 wire _24281_;
 wire _24282_;
 wire _24283_;
 wire _24284_;
 wire _24285_;
 wire _24286_;
 wire _24287_;
 wire _24288_;
 wire _24289_;
 wire _24290_;
 wire _24291_;
 wire _24292_;
 wire _24293_;
 wire _24294_;
 wire _24295_;
 wire _24296_;
 wire _24297_;
 wire _24298_;
 wire _24299_;
 wire _24300_;
 wire _24301_;
 wire _24302_;
 wire _24303_;
 wire _24304_;
 wire _24305_;
 wire _24306_;
 wire _24307_;
 wire _24308_;
 wire _24309_;
 wire _24310_;
 wire _24311_;
 wire _24312_;
 wire _24313_;
 wire _24314_;
 wire _24315_;
 wire _24316_;
 wire _24317_;
 wire _24318_;
 wire _24319_;
 wire _24320_;
 wire _24321_;
 wire _24322_;
 wire _24323_;
 wire _24324_;
 wire _24325_;
 wire _24326_;
 wire _24327_;
 wire _24328_;
 wire _24329_;
 wire _24330_;
 wire _24331_;
 wire _24332_;
 wire _24333_;
 wire _24334_;
 wire _24335_;
 wire _24336_;
 wire _24337_;
 wire _24338_;
 wire _24339_;
 wire _24340_;
 wire _24341_;
 wire _24342_;
 wire _24343_;
 wire _24344_;
 wire _24345_;
 wire _24346_;
 wire _24347_;
 wire _24348_;
 wire _24349_;
 wire _24350_;
 wire _24351_;
 wire _24352_;
 wire _24353_;
 wire _24354_;
 wire _24355_;
 wire _24356_;
 wire _24357_;
 wire _24358_;
 wire _24359_;
 wire _24360_;
 wire _24361_;
 wire _24362_;
 wire _24363_;
 wire _24364_;
 wire _24365_;
 wire _24366_;
 wire _24367_;
 wire _24368_;
 wire _24369_;
 wire _24370_;
 wire _24371_;
 wire _24372_;
 wire _24373_;
 wire _24374_;
 wire _24375_;
 wire _24376_;
 wire _24377_;
 wire _24378_;
 wire _24379_;
 wire _24380_;
 wire _24381_;
 wire _24382_;
 wire _24383_;
 wire _24384_;
 wire _24385_;
 wire _24386_;
 wire _24387_;
 wire _24388_;
 wire _24389_;
 wire _24390_;
 wire _24391_;
 wire _24392_;
 wire _24393_;
 wire _24394_;
 wire _24395_;
 wire _24396_;
 wire _24397_;
 wire _24398_;
 wire _24399_;
 wire _24400_;
 wire _24401_;
 wire _24402_;
 wire _24403_;
 wire _24404_;
 wire _24405_;
 wire _24406_;
 wire _24407_;
 wire _24408_;
 wire _24409_;
 wire _24410_;
 wire _24411_;
 wire _24412_;
 wire _24413_;
 wire _24414_;
 wire _24415_;
 wire _24416_;
 wire _24417_;
 wire _24418_;
 wire _24419_;
 wire _24420_;
 wire _24421_;
 wire _24422_;
 wire _24423_;
 wire _24424_;
 wire _24425_;
 wire _24426_;
 wire _24427_;
 wire _24428_;
 wire _24429_;
 wire _24430_;
 wire _24431_;
 wire _24432_;
 wire _24433_;
 wire _24434_;
 wire _24435_;
 wire _24436_;
 wire _24437_;
 wire _24438_;
 wire _24439_;
 wire _24440_;
 wire _24441_;
 wire _24442_;
 wire _24443_;
 wire _24444_;
 wire _24445_;
 wire _24446_;
 wire _24447_;
 wire _24448_;
 wire _24449_;
 wire _24450_;
 wire _24451_;
 wire _24452_;
 wire _24453_;
 wire _24454_;
 wire _24455_;
 wire _24456_;
 wire _24457_;
 wire _24458_;
 wire _24459_;
 wire _24460_;
 wire _24461_;
 wire _24462_;
 wire _24463_;
 wire _24464_;
 wire _24465_;
 wire _24466_;
 wire _24467_;
 wire _24468_;
 wire _24469_;
 wire _24470_;
 wire _24471_;
 wire _24472_;
 wire _24473_;
 wire _24474_;
 wire _24475_;
 wire _24476_;
 wire _24477_;
 wire _24478_;
 wire _24479_;
 wire _24480_;
 wire _24481_;
 wire _24482_;
 wire _24483_;
 wire _24484_;
 wire _24485_;
 wire _24486_;
 wire _24487_;
 wire _24488_;
 wire _24489_;
 wire _24490_;
 wire _24491_;
 wire _24492_;
 wire _24493_;
 wire _24494_;
 wire _24495_;
 wire _24496_;
 wire _24497_;
 wire _24498_;
 wire _24499_;
 wire _24500_;
 wire _24501_;
 wire _24502_;
 wire _24503_;
 wire _24504_;
 wire _24505_;
 wire _24506_;
 wire _24507_;
 wire _24508_;
 wire _24509_;
 wire _24510_;
 wire _24511_;
 wire _24512_;
 wire _24513_;
 wire _24514_;
 wire _24515_;
 wire _24516_;
 wire _24517_;
 wire _24518_;
 wire _24519_;
 wire _24520_;
 wire _24521_;
 wire _24522_;
 wire _24523_;
 wire _24524_;
 wire _24525_;
 wire _24526_;
 wire _24527_;
 wire _24528_;
 wire _24529_;
 wire _24530_;
 wire _24531_;
 wire _24532_;
 wire _24533_;
 wire _24534_;
 wire _24535_;
 wire _24536_;
 wire _24537_;
 wire _24538_;
 wire _24539_;
 wire _24540_;
 wire _24541_;
 wire _24542_;
 wire _24543_;
 wire _24544_;
 wire _24545_;
 wire _24546_;
 wire _24547_;
 wire _24548_;
 wire _24549_;
 wire _24550_;
 wire _24551_;
 wire _24552_;
 wire _24553_;
 wire _24554_;
 wire _24555_;
 wire _24556_;
 wire _24557_;
 wire _24558_;
 wire _24559_;
 wire _24560_;
 wire _24561_;
 wire _24562_;
 wire _24563_;
 wire _24564_;
 wire _24565_;
 wire _24566_;
 wire _24567_;
 wire _24568_;
 wire _24569_;
 wire _24570_;
 wire _24571_;
 wire _24572_;
 wire _24573_;
 wire _24574_;
 wire _24575_;
 wire _24576_;
 wire _24577_;
 wire _24578_;
 wire _24579_;
 wire _24580_;
 wire _24581_;
 wire _24582_;
 wire _24583_;
 wire _24584_;
 wire _24585_;
 wire _24586_;
 wire _24587_;
 wire _24588_;
 wire _24589_;
 wire _24590_;
 wire _24591_;
 wire _24592_;
 wire _24593_;
 wire _24594_;
 wire _24595_;
 wire _24596_;
 wire _24597_;
 wire _24598_;
 wire _24599_;
 wire _24600_;
 wire _24601_;
 wire _24602_;
 wire _24603_;
 wire _24604_;
 wire _24605_;
 wire _24606_;
 wire _24607_;
 wire _24608_;
 wire _24609_;
 wire _24610_;
 wire _24611_;
 wire _24612_;
 wire _24613_;
 wire _24614_;
 wire _24615_;
 wire _24616_;
 wire _24617_;
 wire _24618_;
 wire _24619_;
 wire _24620_;
 wire _24621_;
 wire _24622_;
 wire _24623_;
 wire _24624_;
 wire _24625_;
 wire _24626_;
 wire _24627_;
 wire _24628_;
 wire _24629_;
 wire _24630_;
 wire _24631_;
 wire _24632_;
 wire _24633_;
 wire _24634_;
 wire _24635_;
 wire _24636_;
 wire _24637_;
 wire _24638_;
 wire _24639_;
 wire _24640_;
 wire _24641_;
 wire _24642_;
 wire _24643_;
 wire _24644_;
 wire _24645_;
 wire _24646_;
 wire _24647_;
 wire _24648_;
 wire _24649_;
 wire _24650_;
 wire _24651_;
 wire _24652_;
 wire _24653_;
 wire _24654_;
 wire _24655_;
 wire _24656_;
 wire _24657_;
 wire _24658_;
 wire _24659_;
 wire _24660_;
 wire _24661_;
 wire _24662_;
 wire _24663_;
 wire _24664_;
 wire _24665_;
 wire _24666_;
 wire _24667_;
 wire _24668_;
 wire _24669_;
 wire _24670_;
 wire _24671_;
 wire _24672_;
 wire _24673_;
 wire _24674_;
 wire _24675_;
 wire _24676_;
 wire _24677_;
 wire _24678_;
 wire _24679_;
 wire _24680_;
 wire _24681_;
 wire _24682_;
 wire _24683_;
 wire _24684_;
 wire _24685_;
 wire _24686_;
 wire _24687_;
 wire _24688_;
 wire _24689_;
 wire _24690_;
 wire _24691_;
 wire _24692_;
 wire _24693_;
 wire _24694_;
 wire _24695_;
 wire _24696_;
 wire _24697_;
 wire _24698_;
 wire _24699_;
 wire _24700_;
 wire _24701_;
 wire _24702_;
 wire _24703_;
 wire _24704_;
 wire _24705_;
 wire _24706_;
 wire _24707_;
 wire _24708_;
 wire _24709_;
 wire _24710_;
 wire _24711_;
 wire _24712_;
 wire _24713_;
 wire _24714_;
 wire _24715_;
 wire _24716_;
 wire _24717_;
 wire _24718_;
 wire _24719_;
 wire _24720_;
 wire _24721_;
 wire _24722_;
 wire _24723_;
 wire _24724_;
 wire _24725_;
 wire _24726_;
 wire _24727_;
 wire _24728_;
 wire _24729_;
 wire _24730_;
 wire _24731_;
 wire _24732_;
 wire _24733_;
 wire _24734_;
 wire _24735_;
 wire _24736_;
 wire _24737_;
 wire _24738_;
 wire _24739_;
 wire _24740_;
 wire _24741_;
 wire _24742_;
 wire _24743_;
 wire _24744_;
 wire _24745_;
 wire _24746_;
 wire _24747_;
 wire _24748_;
 wire _24749_;
 wire _24750_;
 wire _24751_;
 wire _24752_;
 wire _24753_;
 wire _24754_;
 wire _24755_;
 wire _24756_;
 wire _24757_;
 wire _24758_;
 wire _24759_;
 wire _24760_;
 wire _24761_;
 wire _24762_;
 wire _24763_;
 wire _24764_;
 wire _24765_;
 wire _24766_;
 wire _24767_;
 wire _24768_;
 wire _24769_;
 wire _24770_;
 wire _24771_;
 wire _24772_;
 wire _24773_;
 wire _24774_;
 wire _24775_;
 wire _24776_;
 wire _24777_;
 wire _24778_;
 wire _24779_;
 wire _24780_;
 wire _24781_;
 wire _24782_;
 wire _24783_;
 wire _24784_;
 wire _24785_;
 wire _24786_;
 wire _24787_;
 wire _24788_;
 wire _24789_;
 wire _24790_;
 wire _24791_;
 wire _24792_;
 wire _24793_;
 wire _24794_;
 wire _24795_;
 wire _24796_;
 wire _24797_;
 wire _24798_;
 wire _24799_;
 wire _24800_;
 wire _24801_;
 wire _24802_;
 wire _24803_;
 wire _24804_;
 wire _24805_;
 wire _24806_;
 wire _24807_;
 wire _24808_;
 wire _24809_;
 wire _24810_;
 wire _24811_;
 wire _24812_;
 wire _24813_;
 wire _24814_;
 wire _24815_;
 wire _24816_;
 wire _24817_;
 wire _24818_;
 wire _24819_;
 wire _24820_;
 wire _24821_;
 wire _24822_;
 wire _24823_;
 wire _24824_;
 wire _24825_;
 wire _24826_;
 wire _24827_;
 wire _24828_;
 wire _24829_;
 wire _24830_;
 wire _24831_;
 wire _24832_;
 wire _24833_;
 wire _24834_;
 wire _24835_;
 wire _24836_;
 wire _24837_;
 wire _24838_;
 wire _24839_;
 wire _24840_;
 wire _24841_;
 wire _24842_;
 wire _24843_;
 wire _24844_;
 wire _24845_;
 wire _24846_;
 wire _24847_;
 wire _24848_;
 wire _24849_;
 wire _24850_;
 wire _24851_;
 wire _24852_;
 wire _24853_;
 wire _24854_;
 wire _24855_;
 wire _24856_;
 wire _24857_;
 wire _24858_;
 wire _24859_;
 wire _24860_;
 wire _24861_;
 wire _24862_;
 wire _24863_;
 wire _24864_;
 wire _24865_;
 wire _24866_;
 wire _24867_;
 wire _24868_;
 wire _24869_;
 wire _24870_;
 wire _24871_;
 wire _24872_;
 wire _24873_;
 wire _24874_;
 wire _24875_;
 wire _24876_;
 wire _24877_;
 wire _24878_;
 wire _24879_;
 wire _24880_;
 wire _24881_;
 wire _24882_;
 wire _24883_;
 wire _24884_;
 wire _24885_;
 wire _24886_;
 wire _24887_;
 wire _24888_;
 wire _24889_;
 wire _24890_;
 wire _24891_;
 wire _24892_;
 wire _24893_;
 wire _24894_;
 wire _24895_;
 wire _24896_;
 wire _24897_;
 wire _24898_;
 wire _24899_;
 wire _24900_;
 wire _24901_;
 wire _24902_;
 wire _24903_;
 wire _24904_;
 wire _24905_;
 wire _24906_;
 wire _24907_;
 wire _24908_;
 wire _24909_;
 wire _24910_;
 wire _24911_;
 wire _24912_;
 wire _24913_;
 wire _24914_;
 wire _24915_;
 wire _24916_;
 wire _24917_;
 wire _24918_;
 wire _24919_;
 wire _24920_;
 wire _24921_;
 wire _24922_;
 wire _24923_;
 wire _24924_;
 wire _24925_;
 wire _24926_;
 wire _24927_;
 wire _24928_;
 wire _24929_;
 wire _24930_;
 wire _24931_;
 wire _24932_;
 wire _24933_;
 wire _24934_;
 wire _24935_;
 wire _24936_;
 wire _24937_;
 wire _24938_;
 wire _24939_;
 wire _24940_;
 wire _24941_;
 wire _24942_;
 wire _24943_;
 wire _24944_;
 wire _24945_;
 wire _24946_;
 wire _24947_;
 wire _24948_;
 wire _24949_;
 wire _24950_;
 wire _24951_;
 wire _24952_;
 wire _24953_;
 wire _24954_;
 wire _24955_;
 wire _24956_;
 wire _24957_;
 wire _24958_;
 wire _24959_;
 wire _24960_;
 wire _24961_;
 wire _24962_;
 wire _24963_;
 wire _24964_;
 wire _24965_;
 wire _24966_;
 wire _24967_;
 wire _24968_;
 wire _24969_;
 wire _24970_;
 wire _24971_;
 wire _24972_;
 wire _24973_;
 wire _24974_;
 wire _24975_;
 wire _24976_;
 wire _24977_;
 wire _24978_;
 wire _24979_;
 wire _24980_;
 wire _24981_;
 wire _24982_;
 wire _24983_;
 wire _24984_;
 wire _24985_;
 wire _24986_;
 wire _24987_;
 wire _24988_;
 wire _24989_;
 wire _24990_;
 wire _24991_;
 wire _24992_;
 wire _24993_;
 wire _24994_;
 wire _24995_;
 wire _24996_;
 wire _24997_;
 wire _24998_;
 wire _24999_;
 wire _25000_;
 wire _25001_;
 wire _25002_;
 wire _25003_;
 wire _25004_;
 wire _25005_;
 wire _25006_;
 wire _25007_;
 wire _25008_;
 wire _25009_;
 wire _25010_;
 wire _25011_;
 wire _25012_;
 wire _25013_;
 wire _25014_;
 wire _25015_;
 wire _25016_;
 wire _25017_;
 wire _25018_;
 wire _25019_;
 wire _25020_;
 wire _25021_;
 wire _25022_;
 wire _25023_;
 wire _25024_;
 wire _25025_;
 wire _25026_;
 wire _25027_;
 wire _25028_;
 wire _25029_;
 wire _25030_;
 wire _25031_;
 wire _25032_;
 wire _25033_;
 wire _25034_;
 wire _25035_;
 wire _25036_;
 wire _25037_;
 wire _25038_;
 wire _25039_;
 wire _25040_;
 wire _25041_;
 wire _25042_;
 wire _25043_;
 wire _25044_;
 wire _25045_;
 wire _25046_;
 wire _25047_;
 wire _25048_;
 wire _25049_;
 wire _25050_;
 wire _25051_;
 wire _25052_;
 wire _25053_;
 wire _25054_;
 wire _25055_;
 wire _25056_;
 wire _25057_;
 wire _25058_;
 wire _25059_;
 wire _25060_;
 wire _25061_;
 wire _25062_;
 wire _25063_;
 wire _25064_;
 wire _25065_;
 wire _25066_;
 wire _25067_;
 wire _25068_;
 wire _25069_;
 wire _25070_;
 wire _25071_;
 wire _25072_;
 wire _25073_;
 wire _25074_;
 wire _25075_;
 wire _25076_;
 wire _25077_;
 wire _25078_;
 wire _25079_;
 wire _25080_;
 wire _25081_;
 wire _25082_;
 wire _25083_;
 wire _25084_;
 wire _25085_;
 wire _25086_;
 wire _25087_;
 wire _25088_;
 wire _25089_;
 wire _25090_;
 wire _25091_;
 wire _25092_;
 wire _25093_;
 wire _25094_;
 wire _25095_;
 wire _25096_;
 wire _25097_;
 wire _25098_;
 wire _25099_;
 wire _25100_;
 wire _25101_;
 wire _25102_;
 wire _25103_;
 wire _25104_;
 wire _25105_;
 wire _25106_;
 wire _25107_;
 wire _25108_;
 wire _25109_;
 wire _25110_;
 wire _25111_;
 wire _25112_;
 wire _25113_;
 wire _25114_;
 wire _25115_;
 wire _25116_;
 wire _25117_;
 wire _25118_;
 wire _25119_;
 wire _25120_;
 wire _25121_;
 wire _25122_;
 wire _25123_;
 wire _25124_;
 wire _25125_;
 wire _25126_;
 wire _25127_;
 wire _25128_;
 wire _25129_;
 wire _25130_;
 wire _25131_;
 wire _25132_;
 wire _25133_;
 wire _25134_;
 wire _25135_;
 wire _25136_;
 wire _25137_;
 wire _25138_;
 wire _25139_;
 wire _25140_;
 wire _25141_;
 wire _25142_;
 wire _25143_;
 wire _25144_;
 wire _25145_;
 wire _25146_;
 wire _25147_;
 wire _25148_;
 wire _25149_;
 wire _25150_;
 wire _25151_;
 wire _25152_;
 wire _25153_;
 wire _25154_;
 wire _25155_;
 wire _25156_;
 wire _25157_;
 wire _25158_;
 wire _25159_;
 wire _25160_;
 wire _25161_;
 wire _25162_;
 wire _25163_;
 wire _25164_;
 wire _25165_;
 wire _25166_;
 wire _25167_;
 wire _25168_;
 wire _25169_;
 wire _25170_;
 wire _25171_;
 wire _25172_;
 wire _25173_;
 wire _25174_;
 wire _25175_;
 wire _25176_;
 wire _25177_;
 wire _25178_;
 wire _25179_;
 wire _25180_;
 wire _25181_;
 wire _25182_;
 wire _25183_;
 wire _25184_;
 wire _25185_;
 wire _25186_;
 wire _25187_;
 wire _25188_;
 wire _25189_;
 wire _25190_;
 wire _25191_;
 wire _25192_;
 wire _25193_;
 wire _25194_;
 wire _25195_;
 wire _25196_;
 wire _25197_;
 wire _25198_;
 wire _25199_;
 wire _25200_;
 wire _25201_;
 wire _25202_;
 wire _25203_;
 wire _25204_;
 wire _25205_;
 wire _25206_;
 wire _25207_;
 wire _25208_;
 wire _25209_;
 wire _25210_;
 wire _25211_;
 wire _25212_;
 wire _25213_;
 wire _25214_;
 wire _25215_;
 wire _25216_;
 wire _25217_;
 wire _25218_;
 wire _25219_;
 wire _25220_;
 wire _25221_;
 wire _25222_;
 wire _25223_;
 wire _25224_;
 wire _25225_;
 wire _25226_;
 wire _25227_;
 wire _25228_;
 wire _25229_;
 wire _25230_;
 wire _25231_;
 wire _25232_;
 wire _25233_;
 wire _25234_;
 wire _25235_;
 wire _25236_;
 wire _25237_;
 wire _25238_;
 wire _25239_;
 wire _25240_;
 wire _25241_;
 wire _25242_;
 wire _25243_;
 wire _25244_;
 wire _25245_;
 wire _25246_;
 wire _25247_;
 wire _25248_;
 wire _25249_;
 wire _25250_;
 wire _25251_;
 wire _25252_;
 wire _25253_;
 wire _25254_;
 wire _25255_;
 wire _25256_;
 wire _25257_;
 wire _25258_;
 wire _25259_;
 wire _25260_;
 wire _25261_;
 wire _25262_;
 wire _25263_;
 wire _25264_;
 wire _25265_;
 wire _25266_;
 wire _25267_;
 wire _25268_;
 wire _25269_;
 wire _25270_;
 wire _25271_;
 wire _25272_;
 wire _25273_;
 wire _25274_;
 wire _25275_;
 wire _25276_;
 wire _25277_;
 wire _25278_;
 wire _25279_;
 wire _25280_;
 wire _25281_;
 wire _25282_;
 wire _25283_;
 wire _25284_;
 wire _25285_;
 wire _25286_;
 wire _25287_;
 wire _25288_;
 wire _25289_;
 wire _25290_;
 wire _25291_;
 wire _25292_;
 wire _25293_;
 wire _25294_;
 wire _25295_;
 wire _25296_;
 wire _25297_;
 wire _25298_;
 wire _25299_;
 wire _25300_;
 wire _25301_;
 wire _25302_;
 wire _25303_;
 wire _25304_;
 wire _25305_;
 wire _25306_;
 wire _25307_;
 wire _25308_;
 wire _25309_;
 wire _25310_;
 wire _25311_;
 wire _25312_;
 wire _25313_;
 wire _25314_;
 wire _25315_;
 wire _25316_;
 wire _25317_;
 wire _25318_;
 wire _25319_;
 wire _25320_;
 wire _25321_;
 wire _25322_;
 wire _25323_;
 wire _25324_;
 wire _25325_;
 wire _25326_;
 wire _25327_;
 wire _25328_;
 wire _25329_;
 wire _25330_;
 wire _25331_;
 wire _25332_;
 wire _25333_;
 wire _25334_;
 wire _25335_;
 wire _25336_;
 wire _25337_;
 wire _25338_;
 wire _25339_;
 wire _25340_;
 wire _25341_;
 wire _25342_;
 wire _25343_;
 wire _25344_;
 wire _25345_;
 wire _25346_;
 wire _25347_;
 wire _25348_;
 wire _25349_;
 wire _25350_;
 wire _25351_;
 wire _25352_;
 wire _25353_;
 wire _25354_;
 wire _25355_;
 wire _25356_;
 wire _25357_;
 wire _25358_;
 wire _25359_;
 wire _25360_;
 wire _25361_;
 wire _25362_;
 wire _25363_;
 wire _25364_;
 wire _25365_;
 wire _25366_;
 wire _25367_;
 wire _25368_;
 wire _25369_;
 wire _25370_;
 wire _25371_;
 wire _25372_;
 wire _25373_;
 wire _25374_;
 wire _25375_;
 wire _25376_;
 wire _25377_;
 wire _25378_;
 wire _25379_;
 wire _25380_;
 wire _25381_;
 wire _25382_;
 wire _25383_;
 wire _25384_;
 wire _25385_;
 wire _25386_;
 wire _25387_;
 wire _25388_;
 wire _25389_;
 wire _25390_;
 wire _25391_;
 wire _25392_;
 wire _25393_;
 wire _25394_;
 wire _25395_;
 wire _25396_;
 wire _25397_;
 wire _25398_;
 wire _25399_;
 wire _25400_;
 wire _25401_;
 wire _25402_;
 wire _25403_;
 wire _25404_;
 wire _25405_;
 wire _25406_;
 wire _25407_;
 wire _25408_;
 wire _25409_;
 wire _25410_;
 wire _25411_;
 wire _25412_;
 wire _25413_;
 wire _25414_;
 wire _25415_;
 wire _25416_;
 wire _25417_;
 wire _25418_;
 wire _25419_;
 wire _25420_;
 wire _25421_;
 wire _25422_;
 wire _25423_;
 wire _25424_;
 wire _25425_;
 wire _25426_;
 wire _25427_;
 wire _25428_;
 wire _25429_;
 wire _25430_;
 wire _25431_;
 wire _25432_;
 wire _25433_;
 wire _25434_;
 wire _25435_;
 wire _25436_;
 wire _25437_;
 wire _25438_;
 wire _25439_;
 wire _25440_;
 wire _25441_;
 wire _25442_;
 wire _25443_;
 wire _25444_;
 wire _25445_;
 wire _25446_;
 wire \delay_line[0][0] ;
 wire \delay_line[0][10] ;
 wire \delay_line[0][11] ;
 wire \delay_line[0][12] ;
 wire \delay_line[0][13] ;
 wire \delay_line[0][14] ;
 wire \delay_line[0][15] ;
 wire \delay_line[0][1] ;
 wire \delay_line[0][2] ;
 wire \delay_line[0][3] ;
 wire \delay_line[0][4] ;
 wire \delay_line[0][5] ;
 wire \delay_line[0][6] ;
 wire \delay_line[0][7] ;
 wire \delay_line[0][8] ;
 wire \delay_line[0][9] ;
 wire \delay_line[10][0] ;
 wire \delay_line[10][10] ;
 wire \delay_line[10][11] ;
 wire \delay_line[10][12] ;
 wire \delay_line[10][13] ;
 wire \delay_line[10][14] ;
 wire \delay_line[10][15] ;
 wire \delay_line[10][1] ;
 wire \delay_line[10][2] ;
 wire \delay_line[10][3] ;
 wire \delay_line[10][4] ;
 wire \delay_line[10][5] ;
 wire \delay_line[10][6] ;
 wire \delay_line[10][7] ;
 wire \delay_line[10][8] ;
 wire \delay_line[10][9] ;
 wire \delay_line[11][0] ;
 wire \delay_line[11][10] ;
 wire \delay_line[11][11] ;
 wire \delay_line[11][12] ;
 wire \delay_line[11][13] ;
 wire \delay_line[11][14] ;
 wire \delay_line[11][15] ;
 wire \delay_line[11][1] ;
 wire \delay_line[11][2] ;
 wire \delay_line[11][3] ;
 wire \delay_line[11][4] ;
 wire \delay_line[11][5] ;
 wire \delay_line[11][6] ;
 wire \delay_line[11][7] ;
 wire \delay_line[11][8] ;
 wire \delay_line[11][9] ;
 wire \delay_line[12][0] ;
 wire \delay_line[12][10] ;
 wire \delay_line[12][11] ;
 wire \delay_line[12][12] ;
 wire \delay_line[12][13] ;
 wire \delay_line[12][14] ;
 wire \delay_line[12][15] ;
 wire \delay_line[12][1] ;
 wire \delay_line[12][2] ;
 wire \delay_line[12][3] ;
 wire \delay_line[12][4] ;
 wire \delay_line[12][5] ;
 wire \delay_line[12][6] ;
 wire \delay_line[12][7] ;
 wire \delay_line[12][8] ;
 wire \delay_line[12][9] ;
 wire \delay_line[13][0] ;
 wire \delay_line[13][10] ;
 wire \delay_line[13][11] ;
 wire \delay_line[13][12] ;
 wire \delay_line[13][13] ;
 wire \delay_line[13][14] ;
 wire \delay_line[13][15] ;
 wire \delay_line[13][1] ;
 wire \delay_line[13][2] ;
 wire \delay_line[13][3] ;
 wire \delay_line[13][4] ;
 wire \delay_line[13][5] ;
 wire \delay_line[13][6] ;
 wire \delay_line[13][7] ;
 wire \delay_line[13][8] ;
 wire \delay_line[13][9] ;
 wire \delay_line[14][0] ;
 wire \delay_line[14][10] ;
 wire \delay_line[14][11] ;
 wire \delay_line[14][12] ;
 wire \delay_line[14][13] ;
 wire \delay_line[14][14] ;
 wire \delay_line[14][15] ;
 wire \delay_line[14][1] ;
 wire \delay_line[14][2] ;
 wire \delay_line[14][3] ;
 wire \delay_line[14][4] ;
 wire \delay_line[14][5] ;
 wire \delay_line[14][6] ;
 wire \delay_line[14][7] ;
 wire \delay_line[14][8] ;
 wire \delay_line[14][9] ;
 wire \delay_line[15][0] ;
 wire \delay_line[15][10] ;
 wire \delay_line[15][11] ;
 wire \delay_line[15][12] ;
 wire \delay_line[15][13] ;
 wire \delay_line[15][14] ;
 wire \delay_line[15][15] ;
 wire \delay_line[15][1] ;
 wire \delay_line[15][2] ;
 wire \delay_line[15][3] ;
 wire \delay_line[15][4] ;
 wire \delay_line[15][5] ;
 wire \delay_line[15][6] ;
 wire \delay_line[15][7] ;
 wire \delay_line[15][8] ;
 wire \delay_line[15][9] ;
 wire \delay_line[16][0] ;
 wire \delay_line[16][10] ;
 wire \delay_line[16][11] ;
 wire \delay_line[16][12] ;
 wire \delay_line[16][13] ;
 wire \delay_line[16][14] ;
 wire \delay_line[16][15] ;
 wire \delay_line[16][1] ;
 wire \delay_line[16][2] ;
 wire \delay_line[16][3] ;
 wire \delay_line[16][4] ;
 wire \delay_line[16][5] ;
 wire \delay_line[16][6] ;
 wire \delay_line[16][7] ;
 wire \delay_line[16][8] ;
 wire \delay_line[16][9] ;
 wire \delay_line[17][0] ;
 wire \delay_line[17][10] ;
 wire \delay_line[17][11] ;
 wire \delay_line[17][12] ;
 wire \delay_line[17][13] ;
 wire \delay_line[17][14] ;
 wire \delay_line[17][15] ;
 wire \delay_line[17][1] ;
 wire \delay_line[17][2] ;
 wire \delay_line[17][3] ;
 wire \delay_line[17][4] ;
 wire \delay_line[17][5] ;
 wire \delay_line[17][6] ;
 wire \delay_line[17][7] ;
 wire \delay_line[17][8] ;
 wire \delay_line[17][9] ;
 wire \delay_line[18][0] ;
 wire \delay_line[18][10] ;
 wire \delay_line[18][11] ;
 wire \delay_line[18][12] ;
 wire \delay_line[18][13] ;
 wire \delay_line[18][14] ;
 wire \delay_line[18][15] ;
 wire \delay_line[18][1] ;
 wire \delay_line[18][2] ;
 wire \delay_line[18][3] ;
 wire \delay_line[18][4] ;
 wire \delay_line[18][5] ;
 wire \delay_line[18][6] ;
 wire \delay_line[18][7] ;
 wire \delay_line[18][8] ;
 wire \delay_line[18][9] ;
 wire \delay_line[19][0] ;
 wire \delay_line[19][10] ;
 wire \delay_line[19][11] ;
 wire \delay_line[19][12] ;
 wire \delay_line[19][13] ;
 wire \delay_line[19][14] ;
 wire \delay_line[19][15] ;
 wire \delay_line[19][1] ;
 wire \delay_line[19][2] ;
 wire \delay_line[19][3] ;
 wire \delay_line[19][4] ;
 wire \delay_line[19][5] ;
 wire \delay_line[19][6] ;
 wire \delay_line[19][7] ;
 wire \delay_line[19][8] ;
 wire \delay_line[19][9] ;
 wire \delay_line[1][0] ;
 wire \delay_line[1][10] ;
 wire \delay_line[1][11] ;
 wire \delay_line[1][12] ;
 wire \delay_line[1][13] ;
 wire \delay_line[1][14] ;
 wire \delay_line[1][15] ;
 wire \delay_line[1][1] ;
 wire \delay_line[1][2] ;
 wire \delay_line[1][3] ;
 wire \delay_line[1][4] ;
 wire \delay_line[1][5] ;
 wire \delay_line[1][6] ;
 wire \delay_line[1][7] ;
 wire \delay_line[1][8] ;
 wire \delay_line[1][9] ;
 wire \delay_line[20][0] ;
 wire \delay_line[20][10] ;
 wire \delay_line[20][11] ;
 wire \delay_line[20][12] ;
 wire \delay_line[20][13] ;
 wire \delay_line[20][14] ;
 wire \delay_line[20][15] ;
 wire \delay_line[20][1] ;
 wire \delay_line[20][2] ;
 wire \delay_line[20][3] ;
 wire \delay_line[20][4] ;
 wire \delay_line[20][5] ;
 wire \delay_line[20][6] ;
 wire \delay_line[20][7] ;
 wire \delay_line[20][8] ;
 wire \delay_line[20][9] ;
 wire \delay_line[21][0] ;
 wire \delay_line[21][10] ;
 wire \delay_line[21][11] ;
 wire \delay_line[21][12] ;
 wire \delay_line[21][13] ;
 wire \delay_line[21][14] ;
 wire \delay_line[21][15] ;
 wire \delay_line[21][1] ;
 wire \delay_line[21][2] ;
 wire \delay_line[21][3] ;
 wire \delay_line[21][4] ;
 wire \delay_line[21][5] ;
 wire \delay_line[21][6] ;
 wire \delay_line[21][7] ;
 wire \delay_line[21][8] ;
 wire \delay_line[21][9] ;
 wire \delay_line[22][0] ;
 wire \delay_line[22][10] ;
 wire \delay_line[22][11] ;
 wire \delay_line[22][12] ;
 wire \delay_line[22][13] ;
 wire \delay_line[22][14] ;
 wire \delay_line[22][15] ;
 wire \delay_line[22][1] ;
 wire \delay_line[22][2] ;
 wire \delay_line[22][3] ;
 wire \delay_line[22][4] ;
 wire \delay_line[22][5] ;
 wire \delay_line[22][6] ;
 wire \delay_line[22][7] ;
 wire \delay_line[22][8] ;
 wire \delay_line[22][9] ;
 wire \delay_line[23][0] ;
 wire \delay_line[23][10] ;
 wire \delay_line[23][11] ;
 wire \delay_line[23][12] ;
 wire \delay_line[23][13] ;
 wire \delay_line[23][14] ;
 wire \delay_line[23][15] ;
 wire \delay_line[23][1] ;
 wire \delay_line[23][2] ;
 wire \delay_line[23][3] ;
 wire \delay_line[23][4] ;
 wire \delay_line[23][5] ;
 wire \delay_line[23][6] ;
 wire \delay_line[23][7] ;
 wire \delay_line[23][8] ;
 wire \delay_line[23][9] ;
 wire \delay_line[24][0] ;
 wire \delay_line[24][10] ;
 wire \delay_line[24][11] ;
 wire \delay_line[24][12] ;
 wire \delay_line[24][13] ;
 wire \delay_line[24][14] ;
 wire \delay_line[24][15] ;
 wire \delay_line[24][1] ;
 wire \delay_line[24][2] ;
 wire \delay_line[24][3] ;
 wire \delay_line[24][4] ;
 wire \delay_line[24][5] ;
 wire \delay_line[24][6] ;
 wire \delay_line[24][7] ;
 wire \delay_line[24][8] ;
 wire \delay_line[24][9] ;
 wire \delay_line[25][0] ;
 wire \delay_line[25][10] ;
 wire \delay_line[25][11] ;
 wire \delay_line[25][12] ;
 wire \delay_line[25][13] ;
 wire \delay_line[25][14] ;
 wire \delay_line[25][15] ;
 wire \delay_line[25][1] ;
 wire \delay_line[25][2] ;
 wire \delay_line[25][3] ;
 wire \delay_line[25][4] ;
 wire \delay_line[25][5] ;
 wire \delay_line[25][6] ;
 wire \delay_line[25][7] ;
 wire \delay_line[25][8] ;
 wire \delay_line[25][9] ;
 wire \delay_line[26][0] ;
 wire \delay_line[26][10] ;
 wire \delay_line[26][11] ;
 wire \delay_line[26][12] ;
 wire \delay_line[26][13] ;
 wire \delay_line[26][14] ;
 wire \delay_line[26][15] ;
 wire \delay_line[26][1] ;
 wire \delay_line[26][2] ;
 wire \delay_line[26][3] ;
 wire \delay_line[26][4] ;
 wire \delay_line[26][5] ;
 wire \delay_line[26][6] ;
 wire \delay_line[26][7] ;
 wire \delay_line[26][8] ;
 wire \delay_line[26][9] ;
 wire \delay_line[27][0] ;
 wire \delay_line[27][10] ;
 wire \delay_line[27][11] ;
 wire \delay_line[27][12] ;
 wire \delay_line[27][13] ;
 wire \delay_line[27][14] ;
 wire \delay_line[27][15] ;
 wire \delay_line[27][1] ;
 wire \delay_line[27][2] ;
 wire \delay_line[27][3] ;
 wire \delay_line[27][4] ;
 wire \delay_line[27][5] ;
 wire \delay_line[27][6] ;
 wire \delay_line[27][7] ;
 wire \delay_line[27][8] ;
 wire \delay_line[27][9] ;
 wire \delay_line[28][0] ;
 wire \delay_line[28][10] ;
 wire \delay_line[28][11] ;
 wire \delay_line[28][12] ;
 wire \delay_line[28][13] ;
 wire \delay_line[28][14] ;
 wire \delay_line[28][15] ;
 wire \delay_line[28][1] ;
 wire \delay_line[28][2] ;
 wire \delay_line[28][3] ;
 wire \delay_line[28][4] ;
 wire \delay_line[28][5] ;
 wire \delay_line[28][6] ;
 wire \delay_line[28][7] ;
 wire \delay_line[28][8] ;
 wire \delay_line[28][9] ;
 wire \delay_line[29][0] ;
 wire \delay_line[29][10] ;
 wire \delay_line[29][11] ;
 wire \delay_line[29][12] ;
 wire \delay_line[29][13] ;
 wire \delay_line[29][14] ;
 wire \delay_line[29][15] ;
 wire \delay_line[29][1] ;
 wire \delay_line[29][2] ;
 wire \delay_line[29][3] ;
 wire \delay_line[29][4] ;
 wire \delay_line[29][5] ;
 wire \delay_line[29][6] ;
 wire \delay_line[29][7] ;
 wire \delay_line[29][8] ;
 wire \delay_line[29][9] ;
 wire \delay_line[2][0] ;
 wire \delay_line[2][10] ;
 wire \delay_line[2][11] ;
 wire \delay_line[2][12] ;
 wire \delay_line[2][13] ;
 wire \delay_line[2][14] ;
 wire \delay_line[2][15] ;
 wire \delay_line[2][1] ;
 wire \delay_line[2][2] ;
 wire \delay_line[2][3] ;
 wire \delay_line[2][4] ;
 wire \delay_line[2][5] ;
 wire \delay_line[2][6] ;
 wire \delay_line[2][7] ;
 wire \delay_line[2][8] ;
 wire \delay_line[2][9] ;
 wire \delay_line[30][0] ;
 wire \delay_line[30][10] ;
 wire \delay_line[30][11] ;
 wire \delay_line[30][12] ;
 wire \delay_line[30][13] ;
 wire \delay_line[30][14] ;
 wire \delay_line[30][15] ;
 wire \delay_line[30][1] ;
 wire \delay_line[30][2] ;
 wire \delay_line[30][3] ;
 wire \delay_line[30][4] ;
 wire \delay_line[30][5] ;
 wire \delay_line[30][6] ;
 wire \delay_line[30][7] ;
 wire \delay_line[30][8] ;
 wire \delay_line[30][9] ;
 wire \delay_line[31][0] ;
 wire \delay_line[31][10] ;
 wire \delay_line[31][11] ;
 wire \delay_line[31][12] ;
 wire \delay_line[31][13] ;
 wire \delay_line[31][14] ;
 wire \delay_line[31][15] ;
 wire \delay_line[31][1] ;
 wire \delay_line[31][2] ;
 wire \delay_line[31][3] ;
 wire \delay_line[31][4] ;
 wire \delay_line[31][5] ;
 wire \delay_line[31][6] ;
 wire \delay_line[31][7] ;
 wire \delay_line[31][8] ;
 wire \delay_line[31][9] ;
 wire \delay_line[32][0] ;
 wire \delay_line[32][10] ;
 wire \delay_line[32][11] ;
 wire \delay_line[32][12] ;
 wire \delay_line[32][13] ;
 wire \delay_line[32][14] ;
 wire \delay_line[32][15] ;
 wire \delay_line[32][1] ;
 wire \delay_line[32][2] ;
 wire \delay_line[32][3] ;
 wire \delay_line[32][4] ;
 wire \delay_line[32][5] ;
 wire \delay_line[32][6] ;
 wire \delay_line[32][7] ;
 wire \delay_line[32][8] ;
 wire \delay_line[32][9] ;
 wire \delay_line[33][0] ;
 wire \delay_line[33][10] ;
 wire \delay_line[33][11] ;
 wire \delay_line[33][12] ;
 wire \delay_line[33][13] ;
 wire \delay_line[33][14] ;
 wire \delay_line[33][15] ;
 wire \delay_line[33][1] ;
 wire \delay_line[33][2] ;
 wire \delay_line[33][3] ;
 wire \delay_line[33][4] ;
 wire \delay_line[33][5] ;
 wire \delay_line[33][6] ;
 wire \delay_line[33][7] ;
 wire \delay_line[33][8] ;
 wire \delay_line[33][9] ;
 wire \delay_line[34][0] ;
 wire \delay_line[34][10] ;
 wire \delay_line[34][11] ;
 wire \delay_line[34][12] ;
 wire \delay_line[34][13] ;
 wire \delay_line[34][14] ;
 wire \delay_line[34][15] ;
 wire \delay_line[34][1] ;
 wire \delay_line[34][2] ;
 wire \delay_line[34][3] ;
 wire \delay_line[34][4] ;
 wire \delay_line[34][5] ;
 wire \delay_line[34][6] ;
 wire \delay_line[34][7] ;
 wire \delay_line[34][8] ;
 wire \delay_line[34][9] ;
 wire \delay_line[35][0] ;
 wire \delay_line[35][10] ;
 wire \delay_line[35][11] ;
 wire \delay_line[35][12] ;
 wire \delay_line[35][13] ;
 wire \delay_line[35][14] ;
 wire \delay_line[35][15] ;
 wire \delay_line[35][1] ;
 wire \delay_line[35][2] ;
 wire \delay_line[35][3] ;
 wire \delay_line[35][4] ;
 wire \delay_line[35][5] ;
 wire \delay_line[35][6] ;
 wire \delay_line[35][7] ;
 wire \delay_line[35][8] ;
 wire \delay_line[35][9] ;
 wire \delay_line[36][0] ;
 wire \delay_line[36][10] ;
 wire \delay_line[36][11] ;
 wire \delay_line[36][12] ;
 wire \delay_line[36][13] ;
 wire \delay_line[36][14] ;
 wire \delay_line[36][15] ;
 wire \delay_line[36][1] ;
 wire \delay_line[36][2] ;
 wire \delay_line[36][3] ;
 wire \delay_line[36][4] ;
 wire \delay_line[36][5] ;
 wire \delay_line[36][6] ;
 wire \delay_line[36][7] ;
 wire \delay_line[36][8] ;
 wire \delay_line[36][9] ;
 wire \delay_line[37][0] ;
 wire \delay_line[37][10] ;
 wire \delay_line[37][11] ;
 wire \delay_line[37][12] ;
 wire \delay_line[37][13] ;
 wire \delay_line[37][14] ;
 wire \delay_line[37][15] ;
 wire \delay_line[37][1] ;
 wire \delay_line[37][2] ;
 wire \delay_line[37][3] ;
 wire \delay_line[37][4] ;
 wire \delay_line[37][5] ;
 wire \delay_line[37][6] ;
 wire \delay_line[37][7] ;
 wire \delay_line[37][8] ;
 wire \delay_line[37][9] ;
 wire \delay_line[38][0] ;
 wire \delay_line[38][10] ;
 wire \delay_line[38][11] ;
 wire \delay_line[38][12] ;
 wire \delay_line[38][13] ;
 wire \delay_line[38][14] ;
 wire \delay_line[38][15] ;
 wire \delay_line[38][1] ;
 wire \delay_line[38][2] ;
 wire \delay_line[38][3] ;
 wire \delay_line[38][4] ;
 wire \delay_line[38][5] ;
 wire \delay_line[38][6] ;
 wire \delay_line[38][7] ;
 wire \delay_line[38][8] ;
 wire \delay_line[38][9] ;
 wire \delay_line[39][0] ;
 wire \delay_line[39][10] ;
 wire \delay_line[39][11] ;
 wire \delay_line[39][12] ;
 wire \delay_line[39][13] ;
 wire \delay_line[39][14] ;
 wire \delay_line[39][15] ;
 wire \delay_line[39][1] ;
 wire \delay_line[39][2] ;
 wire \delay_line[39][3] ;
 wire \delay_line[39][4] ;
 wire \delay_line[39][5] ;
 wire \delay_line[39][6] ;
 wire \delay_line[39][7] ;
 wire \delay_line[39][8] ;
 wire \delay_line[39][9] ;
 wire \delay_line[3][0] ;
 wire \delay_line[3][10] ;
 wire \delay_line[3][11] ;
 wire \delay_line[3][12] ;
 wire \delay_line[3][13] ;
 wire \delay_line[3][14] ;
 wire \delay_line[3][15] ;
 wire \delay_line[3][1] ;
 wire \delay_line[3][2] ;
 wire \delay_line[3][3] ;
 wire \delay_line[3][4] ;
 wire \delay_line[3][5] ;
 wire \delay_line[3][6] ;
 wire \delay_line[3][7] ;
 wire \delay_line[3][8] ;
 wire \delay_line[3][9] ;
 wire \delay_line[40][0] ;
 wire \delay_line[40][10] ;
 wire \delay_line[40][11] ;
 wire \delay_line[40][12] ;
 wire \delay_line[40][13] ;
 wire \delay_line[40][14] ;
 wire \delay_line[40][15] ;
 wire \delay_line[40][1] ;
 wire \delay_line[40][2] ;
 wire \delay_line[40][3] ;
 wire \delay_line[40][4] ;
 wire \delay_line[40][5] ;
 wire \delay_line[40][6] ;
 wire \delay_line[40][7] ;
 wire \delay_line[40][8] ;
 wire \delay_line[40][9] ;
 wire \delay_line[4][0] ;
 wire \delay_line[4][10] ;
 wire \delay_line[4][11] ;
 wire \delay_line[4][12] ;
 wire \delay_line[4][13] ;
 wire \delay_line[4][14] ;
 wire \delay_line[4][15] ;
 wire \delay_line[4][1] ;
 wire \delay_line[4][2] ;
 wire \delay_line[4][3] ;
 wire \delay_line[4][4] ;
 wire \delay_line[4][5] ;
 wire \delay_line[4][6] ;
 wire \delay_line[4][7] ;
 wire \delay_line[4][8] ;
 wire \delay_line[4][9] ;
 wire \delay_line[5][0] ;
 wire \delay_line[5][10] ;
 wire \delay_line[5][11] ;
 wire \delay_line[5][12] ;
 wire \delay_line[5][13] ;
 wire \delay_line[5][14] ;
 wire \delay_line[5][15] ;
 wire \delay_line[5][1] ;
 wire \delay_line[5][2] ;
 wire \delay_line[5][3] ;
 wire \delay_line[5][4] ;
 wire \delay_line[5][5] ;
 wire \delay_line[5][6] ;
 wire \delay_line[5][7] ;
 wire \delay_line[5][8] ;
 wire \delay_line[5][9] ;
 wire \delay_line[6][0] ;
 wire \delay_line[6][10] ;
 wire \delay_line[6][11] ;
 wire \delay_line[6][12] ;
 wire \delay_line[6][13] ;
 wire \delay_line[6][14] ;
 wire \delay_line[6][15] ;
 wire \delay_line[6][1] ;
 wire \delay_line[6][2] ;
 wire \delay_line[6][3] ;
 wire \delay_line[6][4] ;
 wire \delay_line[6][5] ;
 wire \delay_line[6][6] ;
 wire \delay_line[6][7] ;
 wire \delay_line[6][8] ;
 wire \delay_line[6][9] ;
 wire \delay_line[7][0] ;
 wire \delay_line[7][10] ;
 wire \delay_line[7][11] ;
 wire \delay_line[7][12] ;
 wire \delay_line[7][13] ;
 wire \delay_line[7][14] ;
 wire \delay_line[7][15] ;
 wire \delay_line[7][1] ;
 wire \delay_line[7][2] ;
 wire \delay_line[7][3] ;
 wire \delay_line[7][4] ;
 wire \delay_line[7][5] ;
 wire \delay_line[7][6] ;
 wire \delay_line[7][7] ;
 wire \delay_line[7][8] ;
 wire \delay_line[7][9] ;
 wire \delay_line[8][0] ;
 wire \delay_line[8][10] ;
 wire \delay_line[8][11] ;
 wire \delay_line[8][12] ;
 wire \delay_line[8][13] ;
 wire \delay_line[8][14] ;
 wire \delay_line[8][15] ;
 wire \delay_line[8][1] ;
 wire \delay_line[8][2] ;
 wire \delay_line[8][3] ;
 wire \delay_line[8][4] ;
 wire \delay_line[8][5] ;
 wire \delay_line[8][6] ;
 wire \delay_line[8][7] ;
 wire \delay_line[8][8] ;
 wire \delay_line[8][9] ;
 wire \delay_line[9][0] ;
 wire \delay_line[9][10] ;
 wire \delay_line[9][11] ;
 wire \delay_line[9][12] ;
 wire \delay_line[9][13] ;
 wire \delay_line[9][14] ;
 wire \delay_line[9][15] ;
 wire \delay_line[9][1] ;
 wire \delay_line[9][2] ;
 wire \delay_line[9][3] ;
 wire \delay_line[9][4] ;
 wire \delay_line[9][5] ;
 wire \delay_line[9][6] ;
 wire \delay_line[9][7] ;
 wire \delay_line[9][8] ;
 wire \delay_line[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;

 sky130_fd_sc_hd__and3_2 _25447_ (.A(_22004_),
    .B(_22002_),
    .C(_22003_),
    .X(_22006_));
 sky130_fd_sc_hd__nor3_1 _25448_ (.A(_21905_),
    .B(_22005_),
    .C(_22006_),
    .Y(_22007_));
 sky130_fd_sc_hd__o21a_1 _25449_ (.A1(_22005_),
    .A2(_22006_),
    .B1(_21905_),
    .X(_22008_));
 sky130_fd_sc_hd__o2bb2ai_2 _25450_ (.A1_N(_21900_),
    .A2_N(_21904_),
    .B1(_22007_),
    .B2(_22008_),
    .Y(_22009_));
 sky130_fd_sc_hd__o21ba_1 _25451_ (.A1(_22005_),
    .A2(_22006_),
    .B1_N(_21905_),
    .X(_22010_));
 sky130_fd_sc_hd__a2111oi_4 _25452_ (.A1(_19881_),
    .A2(_19945_),
    .B1(_19947_),
    .C1(_22005_),
    .D1(_22006_),
    .Y(_22011_));
 sky130_fd_sc_hd__clkbuf_2 _25453_ (.A(_21900_),
    .X(_22012_));
 sky130_fd_sc_hd__o211ai_2 _25454_ (.A1(_22010_),
    .A2(_22011_),
    .B1(_22012_),
    .C1(_21904_),
    .Y(_22013_));
 sky130_fd_sc_hd__inv_2 _25455_ (.A(_20163_),
    .Y(_22014_));
 sky130_fd_sc_hd__a31o_1 _25456_ (.A1(_20167_),
    .A2(_20169_),
    .A3(_19955_),
    .B1(_22014_),
    .X(_22015_));
 sky130_fd_sc_hd__a21oi_1 _25457_ (.A1(_22009_),
    .A2(_22013_),
    .B1(_22015_),
    .Y(_22016_));
 sky130_fd_sc_hd__o21ai_2 _25458_ (.A1(_22010_),
    .A2(_22011_),
    .B1(_22012_),
    .Y(_22017_));
 sky130_fd_sc_hd__and3_2 _25459_ (.A(_21901_),
    .B(_21902_),
    .C(_21903_),
    .X(_22018_));
 sky130_fd_sc_hd__o211a_1 _25460_ (.A1(_22017_),
    .A2(_22018_),
    .B1(_22015_),
    .C1(_22009_),
    .X(_22019_));
 sky130_fd_sc_hd__a21oi_2 _25461_ (.A1(_20218_),
    .A2(_20184_),
    .B1(_20217_),
    .Y(_22020_));
 sky130_fd_sc_hd__nor2b_1 _25462_ (.A(_20191_),
    .B_N(net450),
    .Y(_22021_));
 sky130_fd_sc_hd__nor2_1 _25463_ (.A(_19051_),
    .B(_22021_),
    .Y(_22022_));
 sky130_fd_sc_hd__buf_1 _25464_ (.A(\delay_line[1][8] ),
    .X(_22023_));
 sky130_fd_sc_hd__buf_1 _25465_ (.A(\delay_line[1][7] ),
    .X(_22024_));
 sky130_fd_sc_hd__or2b_1 _25466_ (.A(_22023_),
    .B_N(_22024_),
    .X(_22025_));
 sky130_fd_sc_hd__nand2_1 _25467_ (.A(_22022_),
    .B(_22025_),
    .Y(_22026_));
 sky130_fd_sc_hd__nor2b_2 _25468_ (.A(net450),
    .B_N(_20191_),
    .Y(_22027_));
 sky130_fd_sc_hd__o21ai_1 _25469_ (.A1(_22027_),
    .A2(_22021_),
    .B1(_19051_),
    .Y(_22028_));
 sky130_fd_sc_hd__nand3b_1 _25470_ (.A_N(_20195_),
    .B(_22026_),
    .C(_22028_),
    .Y(_22029_));
 sky130_fd_sc_hd__a21bo_1 _25471_ (.A1(_22026_),
    .A2(_22028_),
    .B1_N(_20195_),
    .X(_22030_));
 sky130_fd_sc_hd__and2_1 _25472_ (.A(_19117_),
    .B(_19122_),
    .X(_22031_));
 sky130_fd_sc_hd__o21a_1 _25473_ (.A1(_19117_),
    .A2(_20186_),
    .B1(_19116_),
    .X(_22032_));
 sky130_fd_sc_hd__nor2_1 _25474_ (.A(_19117_),
    .B(_19121_),
    .Y(_22033_));
 sky130_fd_sc_hd__nand2_1 _25475_ (.A(_19117_),
    .B(_19121_),
    .Y(_22034_));
 sky130_fd_sc_hd__nand3b_1 _25476_ (.A_N(_22033_),
    .B(_22034_),
    .C(_20196_),
    .Y(_22035_));
 sky130_fd_sc_hd__o21ai_1 _25477_ (.A1(_22033_),
    .A2(_22031_),
    .B1(_20194_),
    .Y(_22036_));
 sky130_fd_sc_hd__o211ai_2 _25478_ (.A1(_22031_),
    .A2(_22032_),
    .B1(_22035_),
    .C1(_22036_),
    .Y(_22037_));
 sky130_fd_sc_hd__a211o_1 _25479_ (.A1(_22035_),
    .A2(_22036_),
    .B1(_22031_),
    .C1(_22032_),
    .X(_22038_));
 sky130_fd_sc_hd__nand4_1 _25480_ (.A(_22029_),
    .B(_22030_),
    .C(_22037_),
    .D(_22038_),
    .Y(_22039_));
 sky130_fd_sc_hd__nand2_1 _25481_ (.A(_22029_),
    .B(_22030_),
    .Y(_22040_));
 sky130_fd_sc_hd__nand2_1 _25482_ (.A(_22037_),
    .B(_22038_),
    .Y(_22041_));
 sky130_fd_sc_hd__nand2_1 _25483_ (.A(_22040_),
    .B(_22041_),
    .Y(_22042_));
 sky130_fd_sc_hd__nand2_1 _25484_ (.A(_20198_),
    .B(_20201_),
    .Y(_22043_));
 sky130_fd_sc_hd__a21oi_1 _25485_ (.A1(_22039_),
    .A2(_22042_),
    .B1(_22043_),
    .Y(_22044_));
 sky130_fd_sc_hd__and3_2 _25486_ (.A(_22043_),
    .B(_22039_),
    .C(_22042_),
    .X(_22045_));
 sky130_fd_sc_hd__o21ai_2 _25487_ (.A1(_18172_),
    .A2(_18174_),
    .B1(_19125_),
    .Y(_22046_));
 sky130_fd_sc_hd__o211a_1 _25488_ (.A1(_22044_),
    .A2(_22045_),
    .B1(_22046_),
    .C1(_20189_),
    .X(_22047_));
 sky130_fd_sc_hd__a211oi_2 _25489_ (.A1(_22046_),
    .A2(_20189_),
    .B1(_22044_),
    .C1(_22045_),
    .Y(_22048_));
 sky130_fd_sc_hd__o21bai_1 _25490_ (.A1(_19896_),
    .A2(_19897_),
    .B1_N(_19895_),
    .Y(_22049_));
 sky130_fd_sc_hd__o21bai_1 _25491_ (.A1(_22047_),
    .A2(_22048_),
    .B1_N(_22049_),
    .Y(_22050_));
 sky130_fd_sc_hd__a211o_1 _25492_ (.A1(_22046_),
    .A2(_20189_),
    .B1(_22044_),
    .C1(_22045_),
    .X(_22051_));
 sky130_fd_sc_hd__nand3b_1 _25493_ (.A_N(_22047_),
    .B(_22051_),
    .C(_22049_),
    .Y(_22052_));
 sky130_fd_sc_hd__nand2_1 _25494_ (.A(_22050_),
    .B(_22052_),
    .Y(_22053_));
 sky130_fd_sc_hd__nand2_1 _25495_ (.A(_20204_),
    .B(_20207_),
    .Y(_22054_));
 sky130_fd_sc_hd__xnor2_1 _25496_ (.A(_22053_),
    .B(_22054_),
    .Y(_22055_));
 sky130_fd_sc_hd__o311a_1 _25497_ (.A1(net237),
    .A2(_19076_),
    .A3(_19069_),
    .B1(net147),
    .C1(_19079_),
    .X(_22056_));
 sky130_fd_sc_hd__o21ai_1 _25498_ (.A1(_19900_),
    .A2(_22056_),
    .B1(_19942_),
    .Y(_22057_));
 sky130_fd_sc_hd__nand2_1 _25499_ (.A(_22055_),
    .B(_22057_),
    .Y(_22058_));
 sky130_fd_sc_hd__or2_1 _25500_ (.A(_22057_),
    .B(_22055_),
    .X(_22059_));
 sky130_fd_sc_hd__and2_1 _25501_ (.A(_20211_),
    .B(_20214_),
    .X(_22060_));
 sky130_fd_sc_hd__a21boi_1 _25502_ (.A1(_22058_),
    .A2(_22059_),
    .B1_N(_22060_),
    .Y(_22061_));
 sky130_fd_sc_hd__nand3b_1 _25503_ (.A_N(_22060_),
    .B(_22058_),
    .C(_22059_),
    .Y(_22062_));
 sky130_fd_sc_hd__or2b_1 _25504_ (.A(_22061_),
    .B_N(_22062_),
    .X(_22063_));
 sky130_fd_sc_hd__xor2_2 _25505_ (.A(_22020_),
    .B(_22063_),
    .X(_22064_));
 sky130_fd_sc_hd__xnor2_2 _25506_ (.A(_20175_),
    .B(_22064_),
    .Y(_22065_));
 sky130_fd_sc_hd__xnor2_1 _25507_ (.A(_20220_),
    .B(_22065_),
    .Y(_22066_));
 sky130_fd_sc_hd__o21ai_1 _25508_ (.A1(_22016_),
    .A2(_22019_),
    .B1(_22066_),
    .Y(_22067_));
 sky130_fd_sc_hd__a21o_1 _25509_ (.A1(_22009_),
    .A2(_22013_),
    .B1(_22015_),
    .X(_22068_));
 sky130_fd_sc_hd__nor2_2 _25510_ (.A(_20220_),
    .B(_22065_),
    .Y(_22069_));
 sky130_fd_sc_hd__o21a_1 _25511_ (.A1(_20221_),
    .A2(_20219_),
    .B1(_22065_),
    .X(_22070_));
 sky130_fd_sc_hd__nor2_1 _25512_ (.A(_22069_),
    .B(_22070_),
    .Y(_22071_));
 sky130_fd_sc_hd__o211ai_2 _25513_ (.A1(_22018_),
    .A2(_22017_),
    .B1(_22009_),
    .C1(_22015_),
    .Y(_22072_));
 sky130_fd_sc_hd__nand3_1 _25514_ (.A(_22068_),
    .B(_22071_),
    .C(_22072_),
    .Y(_22073_));
 sky130_fd_sc_hd__nand3_1 _25515_ (.A(_21677_),
    .B(_22067_),
    .C(_22073_),
    .Y(_22074_));
 sky130_fd_sc_hd__clkbuf_2 _25516_ (.A(_22074_),
    .X(_22075_));
 sky130_fd_sc_hd__o21ai_1 _25517_ (.A1(_22016_),
    .A2(_22019_),
    .B1(_22071_),
    .Y(_22076_));
 sky130_fd_sc_hd__a21oi_1 _25518_ (.A1(_20228_),
    .A2(_20182_),
    .B1(_20235_),
    .Y(_22077_));
 sky130_fd_sc_hd__nand3_1 _25519_ (.A(_22068_),
    .B(_22072_),
    .C(_22066_),
    .Y(_22078_));
 sky130_fd_sc_hd__nand3_4 _25520_ (.A(_22076_),
    .B(_22077_),
    .C(_22078_),
    .Y(_22079_));
 sky130_fd_sc_hd__o21ba_2 _25521_ (.A1(_19155_),
    .A2(_20223_),
    .B1_N(_20224_),
    .X(_22080_));
 sky130_fd_sc_hd__a21oi_2 _25522_ (.A1(_22075_),
    .A2(_22079_),
    .B1(_22080_),
    .Y(_22081_));
 sky130_fd_sc_hd__clkbuf_4 _25523_ (.A(_22081_),
    .X(_22082_));
 sky130_fd_sc_hd__a21boi_4 _25524_ (.A1(_20240_),
    .A2(_20244_),
    .B1_N(_20245_),
    .Y(_22083_));
 sky130_fd_sc_hd__a31o_4 _25525_ (.A1(_22075_),
    .A2(_22079_),
    .A3(_22080_),
    .B1(_22083_),
    .X(_22084_));
 sky130_fd_sc_hd__nor2_1 _25526_ (.A(_22082_),
    .B(_22084_),
    .Y(_22085_));
 sky130_fd_sc_hd__a21o_1 _25527_ (.A1(_22075_),
    .A2(_22079_),
    .B1(_22080_),
    .X(_22086_));
 sky130_fd_sc_hd__nand3_2 _25528_ (.A(_22075_),
    .B(_22079_),
    .C(_22080_),
    .Y(_22087_));
 sky130_fd_sc_hd__a21bo_1 _25529_ (.A1(_20240_),
    .A2(_20244_),
    .B1_N(_20245_),
    .X(_22088_));
 sky130_fd_sc_hd__a21oi_4 _25530_ (.A1(_22086_),
    .A2(_22087_),
    .B1(_22088_),
    .Y(_22089_));
 sky130_fd_sc_hd__a2bb2oi_4 _25531_ (.A1_N(_20241_),
    .A2_N(_20247_),
    .B1(_20256_),
    .B2(_20257_),
    .Y(_22090_));
 sky130_fd_sc_hd__o21ai_2 _25532_ (.A1(_22085_),
    .A2(_22089_),
    .B1(_22090_),
    .Y(_22091_));
 sky130_fd_sc_hd__and2_1 _25533_ (.A(net349),
    .B(\delay_line[23][8] ),
    .X(_22092_));
 sky130_fd_sc_hd__nor2_1 _25534_ (.A(net349),
    .B(\delay_line[23][8] ),
    .Y(_22093_));
 sky130_fd_sc_hd__nor2_1 _25535_ (.A(_22092_),
    .B(_22093_),
    .Y(_22094_));
 sky130_fd_sc_hd__and3_1 _25536_ (.A(_22074_),
    .B(_22079_),
    .C(_22080_),
    .X(_22095_));
 sky130_fd_sc_hd__o21ai_4 _25537_ (.A1(_22082_),
    .A2(_22095_),
    .B1(_22083_),
    .Y(_22096_));
 sky130_fd_sc_hd__o2bb2ai_4 _25538_ (.A1_N(_20256_),
    .A2_N(_20257_),
    .B1(_20241_),
    .B2(_20247_),
    .Y(_22097_));
 sky130_fd_sc_hd__o211ai_4 _25539_ (.A1(_22082_),
    .A2(_22084_),
    .B1(_22096_),
    .C1(_22097_),
    .Y(_22098_));
 sky130_fd_sc_hd__nand3_2 _25540_ (.A(_22091_),
    .B(_22094_),
    .C(_22098_),
    .Y(_22099_));
 sky130_fd_sc_hd__o21ai_2 _25541_ (.A1(_22085_),
    .A2(_22089_),
    .B1(_22097_),
    .Y(_22100_));
 sky130_fd_sc_hd__o211ai_4 _25542_ (.A1(_22082_),
    .A2(_22084_),
    .B1(_22096_),
    .C1(_22090_),
    .Y(_22101_));
 sky130_fd_sc_hd__o211ai_2 _25543_ (.A1(_22092_),
    .A2(_22093_),
    .B1(_22100_),
    .C1(_22101_),
    .Y(_22102_));
 sky130_fd_sc_hd__o211ai_4 _25544_ (.A1(_21676_),
    .A2(_20814_),
    .B1(_22099_),
    .C1(_22102_),
    .Y(_22103_));
 sky130_fd_sc_hd__o211ai_1 _25545_ (.A1(_22092_),
    .A2(_22093_),
    .B1(_22098_),
    .C1(_22091_),
    .Y(_22104_));
 sky130_fd_sc_hd__nor2_1 _25546_ (.A(_21676_),
    .B(_20814_),
    .Y(_22105_));
 sky130_fd_sc_hd__nand3_1 _25547_ (.A(_22100_),
    .B(_22101_),
    .C(_22094_),
    .Y(_22106_));
 sky130_fd_sc_hd__nand3_1 _25548_ (.A(_22104_),
    .B(_22105_),
    .C(_22106_),
    .Y(_22107_));
 sky130_fd_sc_hd__clkbuf_2 _25549_ (.A(_22107_),
    .X(_22108_));
 sky130_fd_sc_hd__clkbuf_2 _25550_ (.A(_19204_),
    .X(_22109_));
 sky130_fd_sc_hd__clkbuf_2 _25551_ (.A(_22109_),
    .X(_22110_));
 sky130_fd_sc_hd__clkbuf_2 _25552_ (.A(net349),
    .X(_22111_));
 sky130_fd_sc_hd__o211a_1 _25553_ (.A1(_22109_),
    .A2(_22111_),
    .B1(_20254_),
    .C1(_20258_),
    .X(_22112_));
 sky130_fd_sc_hd__a21o_1 _25554_ (.A1(_22110_),
    .A2(_22111_),
    .B1(_22112_),
    .X(_22113_));
 sky130_fd_sc_hd__a21oi_2 _25555_ (.A1(_22103_),
    .A2(_22108_),
    .B1(_22113_),
    .Y(_22114_));
 sky130_fd_sc_hd__o211a_1 _25556_ (.A1(_20266_),
    .A2(_22112_),
    .B1(_22103_),
    .C1(_22107_),
    .X(_22115_));
 sky130_fd_sc_hd__or2_1 _25557_ (.A(_20859_),
    .B(net103),
    .X(_22116_));
 sky130_fd_sc_hd__o21bai_2 _25558_ (.A1(_22114_),
    .A2(_22115_),
    .B1_N(_22116_),
    .Y(_22117_));
 sky130_fd_sc_hd__a21o_1 _25559_ (.A1(_22103_),
    .A2(_22108_),
    .B1(_22113_),
    .X(_22118_));
 sky130_fd_sc_hd__o211ai_2 _25560_ (.A1(_20266_),
    .A2(_22112_),
    .B1(_22103_),
    .C1(_22108_),
    .Y(_22119_));
 sky130_fd_sc_hd__nand3_1 _25561_ (.A(_22116_),
    .B(_22118_),
    .C(_22119_),
    .Y(_22120_));
 sky130_fd_sc_hd__a21o_1 _25562_ (.A1(_20269_),
    .A2(_20268_),
    .B1(_20275_),
    .X(_22121_));
 sky130_fd_sc_hd__a21oi_4 _25563_ (.A1(_22117_),
    .A2(_22120_),
    .B1(_22121_),
    .Y(_22122_));
 sky130_fd_sc_hd__o21ai_1 _25564_ (.A1(_20859_),
    .A2(net103),
    .B1(_22119_),
    .Y(_22123_));
 sky130_fd_sc_hd__o211a_4 _25565_ (.A1(_22123_),
    .A2(_22114_),
    .B1(_22121_),
    .C1(_22117_),
    .X(_22124_));
 sky130_fd_sc_hd__nor3_1 _25566_ (.A(_21675_),
    .B(_22122_),
    .C(_22124_),
    .Y(_22125_));
 sky130_fd_sc_hd__clkbuf_2 _25567_ (.A(_22125_),
    .X(_22126_));
 sky130_fd_sc_hd__nor2_1 _25568_ (.A(_17896_),
    .B(_22109_),
    .Y(_22127_));
 sky130_fd_sc_hd__and2_1 _25569_ (.A(_17896_),
    .B(_19204_),
    .X(_22128_));
 sky130_fd_sc_hd__buf_1 _25570_ (.A(_19216_),
    .X(_22129_));
 sky130_fd_sc_hd__clkbuf_2 _25571_ (.A(_22129_),
    .X(_22130_));
 sky130_fd_sc_hd__and4bb_1 _25572_ (.A_N(_22127_),
    .B_N(_22128_),
    .C(_15383_),
    .D(_22130_),
    .X(_22131_));
 sky130_fd_sc_hd__o2bb2a_1 _25573_ (.A1_N(_15427_),
    .A2_N(_22130_),
    .B1(_22127_),
    .B2(_22128_),
    .X(_22132_));
 sky130_fd_sc_hd__o21ai_1 _25574_ (.A1(_22122_),
    .A2(_22124_),
    .B1(_21675_),
    .Y(_22133_));
 sky130_fd_sc_hd__o21ai_2 _25575_ (.A1(_22131_),
    .A2(_22132_),
    .B1(_22133_),
    .Y(_22134_));
 sky130_fd_sc_hd__o21a_1 _25576_ (.A1(_20664_),
    .A2(_20867_),
    .B1(_20866_),
    .X(_22135_));
 sky130_fd_sc_hd__o21a_1 _25577_ (.A1(_22122_),
    .A2(_22124_),
    .B1(_21675_),
    .X(_22136_));
 sky130_fd_sc_hd__or2_1 _25578_ (.A(_22131_),
    .B(_22132_),
    .X(_22137_));
 sky130_fd_sc_hd__inv_2 _25579_ (.A(_22137_),
    .Y(_22138_));
 sky130_fd_sc_hd__o21ai_1 _25580_ (.A1(_22125_),
    .A2(_22136_),
    .B1(_22138_),
    .Y(_22140_));
 sky130_fd_sc_hd__o211ai_4 _25581_ (.A1(_22126_),
    .A2(_22134_),
    .B1(_22135_),
    .C1(_22140_),
    .Y(_22141_));
 sky130_fd_sc_hd__nand2_1 _25582_ (.A(_22133_),
    .B(_22138_),
    .Y(_22142_));
 sky130_fd_sc_hd__o21ai_2 _25583_ (.A1(_20664_),
    .A2(_20867_),
    .B1(_20866_),
    .Y(_22143_));
 sky130_fd_sc_hd__o21ai_1 _25584_ (.A1(_22126_),
    .A2(_22136_),
    .B1(_22137_),
    .Y(_22144_));
 sky130_fd_sc_hd__o211ai_2 _25585_ (.A1(_22142_),
    .A2(_22126_),
    .B1(_22143_),
    .C1(_22144_),
    .Y(_22145_));
 sky130_fd_sc_hd__clkbuf_2 _25586_ (.A(_22145_),
    .X(_22146_));
 sky130_fd_sc_hd__a31o_1 _25587_ (.A1(_20291_),
    .A2(_20292_),
    .A3(_20284_),
    .B1(_20871_),
    .X(_22147_));
 sky130_fd_sc_hd__a21oi_2 _25588_ (.A1(_22141_),
    .A2(_22146_),
    .B1(_22147_),
    .Y(_22148_));
 sky130_fd_sc_hd__and3_1 _25589_ (.A(_20291_),
    .B(_20292_),
    .C(_20284_),
    .X(_22149_));
 sky130_fd_sc_hd__o211a_1 _25590_ (.A1(_20871_),
    .A2(_22149_),
    .B1(_22141_),
    .C1(_22145_),
    .X(_22151_));
 sky130_fd_sc_hd__o22ai_4 _25591_ (.A1(_21673_),
    .A2(_21674_),
    .B1(_22148_),
    .B2(_22151_),
    .Y(_22152_));
 sky130_fd_sc_hd__a21o_1 _25592_ (.A1(_22141_),
    .A2(_22146_),
    .B1(_22147_),
    .X(_22153_));
 sky130_fd_sc_hd__o211ai_2 _25593_ (.A1(_20871_),
    .A2(_22149_),
    .B1(_22141_),
    .C1(_22146_),
    .Y(_22154_));
 sky130_fd_sc_hd__nor2_1 _25594_ (.A(_21673_),
    .B(_21674_),
    .Y(_22155_));
 sky130_fd_sc_hd__nand3_1 _25595_ (.A(_22153_),
    .B(_22154_),
    .C(_22155_),
    .Y(_22156_));
 sky130_fd_sc_hd__o21ai_2 _25596_ (.A1(_20300_),
    .A2(_20869_),
    .B1(_20877_),
    .Y(_22157_));
 sky130_fd_sc_hd__a21oi_1 _25597_ (.A1(_22152_),
    .A2(_22156_),
    .B1(_22157_),
    .Y(_22158_));
 sky130_fd_sc_hd__nand2_1 _25598_ (.A(_22154_),
    .B(_22155_),
    .Y(_22159_));
 sky130_fd_sc_hd__o211a_1 _25599_ (.A1(_22148_),
    .A2(_22159_),
    .B1(_22157_),
    .C1(_22152_),
    .X(_22160_));
 sky130_fd_sc_hd__o22ai_2 _25600_ (.A1(_20980_),
    .A2(_20981_),
    .B1(_22158_),
    .B2(_22160_),
    .Y(_22162_));
 sky130_fd_sc_hd__a21o_1 _25601_ (.A1(_20976_),
    .A2(_20977_),
    .B1(_20979_),
    .X(_22163_));
 sky130_fd_sc_hd__nand3_1 _25602_ (.A(_20976_),
    .B(_20977_),
    .C(_20979_),
    .Y(_22164_));
 sky130_fd_sc_hd__nand2_1 _25603_ (.A(_22163_),
    .B(_22164_),
    .Y(_22165_));
 sky130_fd_sc_hd__a21o_1 _25604_ (.A1(_22152_),
    .A2(_22156_),
    .B1(_22157_),
    .X(_22166_));
 sky130_fd_sc_hd__o211ai_2 _25605_ (.A1(_22148_),
    .A2(_22159_),
    .B1(_22157_),
    .C1(_22152_),
    .Y(_22167_));
 sky130_fd_sc_hd__nand3b_1 _25606_ (.A_N(_22165_),
    .B(_22166_),
    .C(_22167_),
    .Y(_22168_));
 sky130_fd_sc_hd__nand3_1 _25607_ (.A(_20925_),
    .B(_22162_),
    .C(_22168_),
    .Y(_22169_));
 sky130_fd_sc_hd__o21bai_1 _25608_ (.A1(_22158_),
    .A2(_22160_),
    .B1_N(_22165_),
    .Y(_22170_));
 sky130_fd_sc_hd__nand3_1 _25609_ (.A(_22165_),
    .B(_22166_),
    .C(_22167_),
    .Y(_22171_));
 sky130_fd_sc_hd__a21boi_1 _25610_ (.A1(_20887_),
    .A2(_20884_),
    .B1_N(_20880_),
    .Y(_22173_));
 sky130_fd_sc_hd__nand3_1 _25611_ (.A(_22170_),
    .B(_22171_),
    .C(_22173_),
    .Y(_22174_));
 sky130_fd_sc_hd__nand2_1 _25612_ (.A(_22169_),
    .B(_22174_),
    .Y(_22175_));
 sky130_fd_sc_hd__nand3_1 _25613_ (.A(_19840_),
    .B(_19836_),
    .C(_19839_),
    .Y(_22176_));
 sky130_fd_sc_hd__buf_1 _25614_ (.A(_11295_),
    .X(_22177_));
 sky130_fd_sc_hd__and2b_1 _25615_ (.A_N(_19827_),
    .B(_19825_),
    .X(_22178_));
 sky130_fd_sc_hd__and3_1 _25616_ (.A(_22177_),
    .B(_11361_),
    .C(_22178_),
    .X(_22179_));
 sky130_fd_sc_hd__nor2_1 _25617_ (.A(_18779_),
    .B(_19828_),
    .Y(_22180_));
 sky130_fd_sc_hd__o211a_1 _25618_ (.A1(_22179_),
    .A2(_22180_),
    .B1(_19823_),
    .C1(_19830_),
    .X(_22181_));
 sky130_fd_sc_hd__a211oi_4 _25619_ (.A1(_19823_),
    .A2(_19830_),
    .B1(_22179_),
    .C1(_22180_),
    .Y(_22182_));
 sky130_fd_sc_hd__o2111a_1 _25620_ (.A1(_22181_),
    .A2(_22182_),
    .B1(_20898_),
    .C1(_18779_),
    .D1(_18823_),
    .X(_22184_));
 sky130_fd_sc_hd__a311oi_4 _25621_ (.A1(_20898_),
    .A2(_18779_),
    .A3(_18823_),
    .B1(_22181_),
    .C1(_22182_),
    .Y(_22185_));
 sky130_fd_sc_hd__or4_1 _25622_ (.A(_19758_),
    .B(_20901_),
    .C(_22184_),
    .D(_22185_),
    .X(_22186_));
 sky130_fd_sc_hd__o22ai_4 _25623_ (.A1(_19758_),
    .A2(_20901_),
    .B1(_22184_),
    .B2(_22185_),
    .Y(_22187_));
 sky130_fd_sc_hd__and2_1 _25624_ (.A(_22186_),
    .B(_22187_),
    .X(_22188_));
 sky130_fd_sc_hd__a21o_1 _25625_ (.A1(_19839_),
    .A2(_22176_),
    .B1(_22188_),
    .X(_22189_));
 sky130_fd_sc_hd__nand3_1 _25626_ (.A(_19839_),
    .B(_22176_),
    .C(_22188_),
    .Y(_22190_));
 sky130_fd_sc_hd__o211a_1 _25627_ (.A1(_20902_),
    .A2(_20903_),
    .B1(_22190_),
    .C1(_20895_),
    .X(_22191_));
 sky130_fd_sc_hd__inv_2 _25628_ (.A(_20904_),
    .Y(_22192_));
 sky130_fd_sc_hd__a22oi_1 _25629_ (.A1(_20895_),
    .A2(_22192_),
    .B1(_22189_),
    .B2(_22190_),
    .Y(_22193_));
 sky130_fd_sc_hd__a21oi_1 _25630_ (.A1(_22189_),
    .A2(_22191_),
    .B1(_22193_),
    .Y(_22195_));
 sky130_fd_sc_hd__nand2_1 _25631_ (.A(_22175_),
    .B(_22195_),
    .Y(_22196_));
 sky130_fd_sc_hd__nand3b_1 _25632_ (.A_N(_22195_),
    .B(_22174_),
    .C(_22169_),
    .Y(_22197_));
 sky130_fd_sc_hd__a21boi_1 _25633_ (.A1(_20889_),
    .A2(_20907_),
    .B1_N(_20892_),
    .Y(_22198_));
 sky130_fd_sc_hd__a21bo_1 _25634_ (.A1(_22196_),
    .A2(_22197_),
    .B1_N(_22198_),
    .X(_22199_));
 sky130_fd_sc_hd__nand3b_1 _25635_ (.A_N(_22198_),
    .B(_22196_),
    .C(_22197_),
    .Y(_22200_));
 sky130_fd_sc_hd__inv_2 _25636_ (.A(_20906_),
    .Y(_22201_));
 sky130_fd_sc_hd__nand2_1 _25637_ (.A(_20893_),
    .B(_22201_),
    .Y(_22202_));
 sky130_fd_sc_hd__o21ai_2 _25638_ (.A1(_20894_),
    .A2(_20905_),
    .B1(_22202_),
    .Y(_22203_));
 sky130_fd_sc_hd__nand3_2 _25639_ (.A(_22199_),
    .B(_22200_),
    .C(_22203_),
    .Y(_22204_));
 sky130_fd_sc_hd__a32oi_2 _25640_ (.A1(_19787_),
    .A2(_20913_),
    .A3(_20914_),
    .B1(_20912_),
    .B2(_19764_),
    .Y(_22206_));
 sky130_fd_sc_hd__a21o_1 _25641_ (.A1(_22199_),
    .A2(_22200_),
    .B1(_22203_),
    .X(_22207_));
 sky130_fd_sc_hd__and2b_1 _25642_ (.A_N(_22206_),
    .B(_22207_),
    .X(_22208_));
 sky130_fd_sc_hd__a21bo_1 _25643_ (.A1(_22204_),
    .A2(_22207_),
    .B1_N(_22206_),
    .X(_22209_));
 sky130_fd_sc_hd__a21boi_1 _25644_ (.A1(_22204_),
    .A2(_22208_),
    .B1_N(_22209_),
    .Y(_22210_));
 sky130_fd_sc_hd__xor2_2 _25645_ (.A(_20924_),
    .B(_22210_),
    .X(_00039_));
 sky130_fd_sc_hd__a22oi_4 _25646_ (.A1(_22208_),
    .A2(_22204_),
    .B1(_20924_),
    .B2(_22209_),
    .Y(_22211_));
 sky130_fd_sc_hd__and3_1 _25647_ (.A(_22163_),
    .B(_22164_),
    .C(_22166_),
    .X(_22212_));
 sky130_fd_sc_hd__a31o_1 _25648_ (.A1(_22153_),
    .A2(_22154_),
    .A3(_22155_),
    .B1(_21673_),
    .X(_22213_));
 sky130_fd_sc_hd__o211a_2 _25649_ (.A1(_21676_),
    .A2(_20814_),
    .B1(_22099_),
    .C1(_22102_),
    .X(_22214_));
 sky130_fd_sc_hd__o21a_1 _25650_ (.A1(_20266_),
    .A2(_22112_),
    .B1(_22108_),
    .X(_22216_));
 sky130_fd_sc_hd__a21o_2 _25651_ (.A1(_21034_),
    .A2(_21082_),
    .B1(_21081_),
    .X(_22217_));
 sky130_fd_sc_hd__inv_2 _25652_ (.A(_22217_),
    .Y(_22218_));
 sky130_fd_sc_hd__a21boi_4 _25653_ (.A1(_21015_),
    .A2(_21030_),
    .B1_N(_21031_),
    .Y(_22219_));
 sky130_fd_sc_hd__inv_2 _25654_ (.A(_22219_),
    .Y(_22220_));
 sky130_fd_sc_hd__o22ai_4 _25655_ (.A1(_22081_),
    .A2(_22084_),
    .B1(_22089_),
    .B2(_22090_),
    .Y(_22221_));
 sky130_fd_sc_hd__or3b_2 _25656_ (.A(_22020_),
    .B(_22061_),
    .C_N(_22062_),
    .X(_22222_));
 sky130_fd_sc_hd__inv_2 _25657_ (.A(_22222_),
    .Y(_22223_));
 sky130_fd_sc_hd__inv_2 _25658_ (.A(_22006_),
    .Y(_22224_));
 sky130_fd_sc_hd__or2_1 _25659_ (.A(_21905_),
    .B(_22005_),
    .X(_22225_));
 sky130_fd_sc_hd__nand2_2 _25660_ (.A(_22058_),
    .B(_22062_),
    .Y(_22227_));
 sky130_fd_sc_hd__a21bo_1 _25661_ (.A1(_22050_),
    .A2(_22054_),
    .B1_N(_22052_),
    .X(_22228_));
 sky130_fd_sc_hd__nand2_1 _25662_ (.A(_22035_),
    .B(_22037_),
    .Y(_22229_));
 sky130_fd_sc_hd__or2b_1 _25663_ (.A(_19121_),
    .B_N(_22024_),
    .X(_22230_));
 sky130_fd_sc_hd__a21oi_2 _25664_ (.A1(_22034_),
    .A2(_22230_),
    .B1(_22027_),
    .Y(_22231_));
 sky130_fd_sc_hd__and2b_1 _25665_ (.A_N(_20186_),
    .B(_22024_),
    .X(_22232_));
 sky130_fd_sc_hd__a211oi_1 _25666_ (.A1(_22025_),
    .A2(_20186_),
    .B1(_22031_),
    .C1(_22232_),
    .Y(_22233_));
 sky130_fd_sc_hd__nor2_1 _25667_ (.A(net450),
    .B(\delay_line[1][9] ),
    .Y(_22234_));
 sky130_fd_sc_hd__buf_1 _25668_ (.A(\delay_line[1][9] ),
    .X(_22235_));
 sky130_fd_sc_hd__nand2_1 _25669_ (.A(_22023_),
    .B(_22235_),
    .Y(_22236_));
 sky130_fd_sc_hd__nand3b_2 _25670_ (.A_N(_22234_),
    .B(_22236_),
    .C(\delay_line[2][6] ),
    .Y(_22238_));
 sky130_fd_sc_hd__and2_2 _25671_ (.A(net450),
    .B(\delay_line[1][9] ),
    .X(_22239_));
 sky130_fd_sc_hd__o21bai_2 _25672_ (.A1(_22234_),
    .A2(_22239_),
    .B1_N(\delay_line[2][6] ),
    .Y(_22240_));
 sky130_fd_sc_hd__o2111ai_2 _25673_ (.A1(_22027_),
    .A2(_22021_),
    .B1(_19051_),
    .C1(_22238_),
    .D1(_22240_),
    .Y(_22241_));
 sky130_fd_sc_hd__a21bo_1 _25674_ (.A1(_22238_),
    .A2(_22240_),
    .B1_N(_22028_),
    .X(_22242_));
 sky130_fd_sc_hd__or4bb_1 _25675_ (.A(_22231_),
    .B(_22233_),
    .C_N(_22241_),
    .D_N(_22242_),
    .X(_22243_));
 sky130_fd_sc_hd__a2bb2o_1 _25676_ (.A1_N(_22231_),
    .A2_N(_22233_),
    .B1(_22241_),
    .B2(_22242_),
    .X(_22244_));
 sky130_fd_sc_hd__o21ai_1 _25677_ (.A1(_22040_),
    .A2(_22041_),
    .B1(_22029_),
    .Y(_22245_));
 sky130_fd_sc_hd__a21o_1 _25678_ (.A1(_22243_),
    .A2(_22244_),
    .B1(_22245_),
    .X(_22246_));
 sky130_fd_sc_hd__nand3_2 _25679_ (.A(_22245_),
    .B(_22243_),
    .C(_22244_),
    .Y(_22247_));
 sky130_fd_sc_hd__nand3_2 _25680_ (.A(_22229_),
    .B(_22246_),
    .C(_22247_),
    .Y(_22249_));
 sky130_fd_sc_hd__a21o_1 _25681_ (.A1(_22246_),
    .A2(_22247_),
    .B1(_22229_),
    .X(_22250_));
 sky130_fd_sc_hd__nor2_1 _25682_ (.A(_21950_),
    .B(_21951_),
    .Y(_22251_));
 sky130_fd_sc_hd__nand2_1 _25683_ (.A(_19891_),
    .B(_19893_),
    .Y(_22252_));
 sky130_fd_sc_hd__a221o_1 _25684_ (.A1(_22249_),
    .A2(_22250_),
    .B1(_22251_),
    .B2(_22252_),
    .C1(_21951_),
    .X(_22253_));
 sky130_fd_sc_hd__o211ai_2 _25685_ (.A1(_21951_),
    .A2(_21952_),
    .B1(_22249_),
    .C1(_22250_),
    .Y(_22254_));
 sky130_fd_sc_hd__a211oi_2 _25686_ (.A1(_22253_),
    .A2(_22254_),
    .B1(_22045_),
    .C1(_22048_),
    .Y(_22255_));
 sky130_fd_sc_hd__o211a_1 _25687_ (.A1(_22045_),
    .A2(_22048_),
    .B1(_22253_),
    .C1(_22254_),
    .X(_22256_));
 sky130_fd_sc_hd__o221ai_4 _25688_ (.A1(_21954_),
    .A2(_22000_),
    .B1(_22255_),
    .B2(_22256_),
    .C1(_21999_),
    .Y(_22257_));
 sky130_fd_sc_hd__inv_2 _25689_ (.A(_22256_),
    .Y(_22258_));
 sky130_fd_sc_hd__o21ai_1 _25690_ (.A1(_21954_),
    .A2(_22000_),
    .B1(_21999_),
    .Y(_22260_));
 sky130_fd_sc_hd__nand3b_1 _25691_ (.A_N(_22255_),
    .B(_22258_),
    .C(_22260_),
    .Y(_22261_));
 sky130_fd_sc_hd__nand2_1 _25692_ (.A(_22257_),
    .B(_22261_),
    .Y(_22262_));
 sky130_fd_sc_hd__xnor2_2 _25693_ (.A(_22228_),
    .B(_22262_),
    .Y(_22263_));
 sky130_fd_sc_hd__xnor2_1 _25694_ (.A(_22227_),
    .B(_22263_),
    .Y(_22264_));
 sky130_fd_sc_hd__a21oi_1 _25695_ (.A1(_22224_),
    .A2(_22225_),
    .B1(_22264_),
    .Y(_22265_));
 sky130_fd_sc_hd__and3_1 _25696_ (.A(_22224_),
    .B(_22225_),
    .C(_22264_),
    .X(_22266_));
 sky130_fd_sc_hd__or2_1 _25697_ (.A(_22265_),
    .B(_22266_),
    .X(_22267_));
 sky130_fd_sc_hd__nor2_1 _25698_ (.A(_22223_),
    .B(_22267_),
    .Y(_22268_));
 sky130_fd_sc_hd__o21a_1 _25699_ (.A1(_22265_),
    .A2(_22266_),
    .B1(_22223_),
    .X(_22269_));
 sky130_fd_sc_hd__inv_2 _25700_ (.A(_22012_),
    .Y(_22271_));
 sky130_fd_sc_hd__o211a_1 _25701_ (.A1(_22010_),
    .A2(_22011_),
    .B1(_22012_),
    .C1(_21904_),
    .X(_22272_));
 sky130_fd_sc_hd__o21ai_1 _25702_ (.A1(_21754_),
    .A2(_21749_),
    .B1(_21756_),
    .Y(_22273_));
 sky130_fd_sc_hd__inv_2 _25703_ (.A(_21731_),
    .Y(_22274_));
 sky130_fd_sc_hd__o21a_1 _25704_ (.A1(_21700_),
    .A2(_21705_),
    .B1(_21709_),
    .X(_22275_));
 sky130_fd_sc_hd__nand2b_1 _25705_ (.A_N(\delay_line[4][6] ),
    .B(_19993_),
    .Y(_22276_));
 sky130_fd_sc_hd__clkbuf_2 _25706_ (.A(\delay_line[4][6] ),
    .X(_22277_));
 sky130_fd_sc_hd__nand2b_2 _25707_ (.A_N(_19993_),
    .B(_22277_),
    .Y(_22278_));
 sky130_fd_sc_hd__o211ai_1 _25708_ (.A1(_21707_),
    .A2(_19996_),
    .B1(_22276_),
    .C1(_22278_),
    .Y(_22279_));
 sky130_fd_sc_hd__clkbuf_4 _25709_ (.A(\delay_line[4][5] ),
    .X(_22280_));
 sky130_fd_sc_hd__nand2_1 _25710_ (.A(_19990_),
    .B(_22280_),
    .Y(_22282_));
 sky130_fd_sc_hd__o21ai_1 _25711_ (.A1(_21707_),
    .A2(_19996_),
    .B1(_22282_),
    .Y(_22283_));
 sky130_fd_sc_hd__nand2_1 _25712_ (.A(_22278_),
    .B(_22276_),
    .Y(_22284_));
 sky130_fd_sc_hd__nand2_1 _25713_ (.A(_22283_),
    .B(_22284_),
    .Y(_22285_));
 sky130_fd_sc_hd__o21a_2 _25714_ (.A1(_21706_),
    .A2(_22279_),
    .B1(_22285_),
    .X(_22286_));
 sky130_fd_sc_hd__inv_2 _25715_ (.A(_21701_),
    .Y(_22287_));
 sky130_fd_sc_hd__or4_2 _25716_ (.A(_22287_),
    .B(_21704_),
    .C(_21699_),
    .D(_18930_),
    .X(_22288_));
 sky130_fd_sc_hd__and3_1 _25717_ (.A(_19994_),
    .B(_19991_),
    .C(_18929_),
    .X(_22289_));
 sky130_fd_sc_hd__nand2_1 _25718_ (.A(_21713_),
    .B(_22289_),
    .Y(_22290_));
 sky130_fd_sc_hd__o2111a_1 _25719_ (.A1(_20015_),
    .A2(_22275_),
    .B1(_22286_),
    .C1(_22288_),
    .D1(_22290_),
    .X(_22291_));
 sky130_fd_sc_hd__o21ai_1 _25720_ (.A1(_19990_),
    .A2(_22280_),
    .B1(_21699_),
    .Y(_22293_));
 sky130_fd_sc_hd__a21boi_2 _25721_ (.A1(_22282_),
    .A2(_22293_),
    .B1_N(_22284_),
    .Y(_22294_));
 sky130_fd_sc_hd__o2111a_1 _25722_ (.A1(_21707_),
    .A2(_19995_),
    .B1(_22282_),
    .C1(_22278_),
    .D1(_22276_),
    .X(_22295_));
 sky130_fd_sc_hd__nor2_1 _25723_ (.A(_21706_),
    .B(_21707_),
    .Y(_22296_));
 sky130_fd_sc_hd__o211ai_1 _25724_ (.A1(_18930_),
    .A2(_21704_),
    .B1(_19996_),
    .C1(_22296_),
    .Y(_22297_));
 sky130_fd_sc_hd__a21oi_1 _25725_ (.A1(_22297_),
    .A2(_21709_),
    .B1(_20015_),
    .Y(_22298_));
 sky130_fd_sc_hd__or3_1 _25726_ (.A(_21704_),
    .B(_21700_),
    .C(_18930_),
    .X(_22299_));
 sky130_fd_sc_hd__o2bb2ai_1 _25727_ (.A1_N(_22289_),
    .A2_N(_21714_),
    .B1(_22287_),
    .B2(_22299_),
    .Y(_22300_));
 sky130_fd_sc_hd__o22ai_1 _25728_ (.A1(_22294_),
    .A2(_22295_),
    .B1(_22298_),
    .B2(_22300_),
    .Y(_22301_));
 sky130_fd_sc_hd__clkbuf_2 _25729_ (.A(_22301_),
    .X(_22302_));
 sky130_fd_sc_hd__and2b_1 _25730_ (.A_N(_17937_),
    .B(\delay_line[11][7] ),
    .X(_22304_));
 sky130_fd_sc_hd__nor2b_1 _25731_ (.A(\delay_line[11][7] ),
    .B_N(_17937_),
    .Y(_22305_));
 sky130_fd_sc_hd__o22ai_4 _25732_ (.A1(_12262_),
    .A2(_21718_),
    .B1(_22304_),
    .B2(_22305_),
    .Y(_22306_));
 sky130_fd_sc_hd__inv_2 _25733_ (.A(\delay_line[11][3] ),
    .Y(_22307_));
 sky130_fd_sc_hd__clkbuf_4 _25734_ (.A(\delay_line[11][7] ),
    .X(_22308_));
 sky130_fd_sc_hd__nand2_2 _25735_ (.A(_22307_),
    .B(_22308_),
    .Y(_22309_));
 sky130_fd_sc_hd__or2b_2 _25736_ (.A(\delay_line[11][7] ),
    .B_N(\delay_line[11][3] ),
    .X(_22310_));
 sky130_fd_sc_hd__nand4_4 _25737_ (.A(_12361_),
    .B(_22309_),
    .C(_22310_),
    .D(_21720_),
    .Y(_22311_));
 sky130_fd_sc_hd__nand4_4 _25738_ (.A(_21722_),
    .B(_21725_),
    .C(_22306_),
    .D(_22311_),
    .Y(_22312_));
 sky130_fd_sc_hd__clkbuf_2 _25739_ (.A(_22309_),
    .X(_22313_));
 sky130_fd_sc_hd__nand3b_2 _25740_ (.A_N(_21725_),
    .B(_22313_),
    .C(_22310_),
    .Y(_22315_));
 sky130_fd_sc_hd__o21a_1 _25741_ (.A1(_08019_),
    .A2(_20004_),
    .B1(_20009_),
    .X(_22316_));
 sky130_fd_sc_hd__nor2_1 _25742_ (.A(_21723_),
    .B(_21724_),
    .Y(_22317_));
 sky130_fd_sc_hd__o2bb2ai_1 _25743_ (.A1_N(_22306_),
    .A2_N(_22311_),
    .B1(_22316_),
    .B2(_22317_),
    .Y(_22318_));
 sky130_fd_sc_hd__nand2_1 _25744_ (.A(_22315_),
    .B(_22318_),
    .Y(_22319_));
 sky130_fd_sc_hd__nand3b_1 _25745_ (.A_N(_20011_),
    .B(_21722_),
    .C(_21726_),
    .Y(_22320_));
 sky130_fd_sc_hd__a2bb2oi_2 _25746_ (.A1_N(_20012_),
    .A2_N(_22312_),
    .B1(_22319_),
    .B2(_22320_),
    .Y(_22321_));
 sky130_fd_sc_hd__nand2_1 _25747_ (.A(_22302_),
    .B(_22321_),
    .Y(_22322_));
 sky130_fd_sc_hd__clkbuf_2 _25748_ (.A(\delay_line[0][9] ),
    .X(_22323_));
 sky130_fd_sc_hd__nor2_1 _25749_ (.A(_20012_),
    .B(_22312_),
    .Y(_22324_));
 sky130_fd_sc_hd__o2bb2a_1 _25750_ (.A1_N(_22315_),
    .A2_N(_22318_),
    .B1(_20018_),
    .B2(_21732_),
    .X(_22326_));
 sky130_fd_sc_hd__and3_1 _25751_ (.A(_19995_),
    .B(_18924_),
    .C(_19992_),
    .X(_22327_));
 sky130_fd_sc_hd__a22oi_4 _25752_ (.A1(_22280_),
    .A2(_22327_),
    .B1(_21714_),
    .B2(_22289_),
    .Y(_22328_));
 sky130_fd_sc_hd__inv_2 _25753_ (.A(_20014_),
    .Y(_22329_));
 sky130_fd_sc_hd__nand2_2 _25754_ (.A(_21713_),
    .B(_22329_),
    .Y(_22330_));
 sky130_fd_sc_hd__a21oi_4 _25755_ (.A1(_22328_),
    .A2(_22330_),
    .B1(_22286_),
    .Y(_22331_));
 sky130_fd_sc_hd__o22ai_2 _25756_ (.A1(_22324_),
    .A2(_22326_),
    .B1(_22291_),
    .B2(_22331_),
    .Y(_22332_));
 sky130_fd_sc_hd__o211ai_4 _25757_ (.A1(_22291_),
    .A2(_22322_),
    .B1(_22323_),
    .C1(_22332_),
    .Y(_22333_));
 sky130_fd_sc_hd__o211ai_1 _25758_ (.A1(_22287_),
    .A2(_22299_),
    .B1(_22290_),
    .C1(_22286_),
    .Y(_22334_));
 sky130_fd_sc_hd__o211a_2 _25759_ (.A1(_22298_),
    .A2(_22334_),
    .B1(_22321_),
    .C1(_22302_),
    .X(_22335_));
 sky130_fd_sc_hd__o2111ai_1 _25760_ (.A1(_20016_),
    .A2(_22275_),
    .B1(_22286_),
    .C1(_22288_),
    .D1(_22290_),
    .Y(_22337_));
 sky130_fd_sc_hd__a21oi_1 _25761_ (.A1(_22337_),
    .A2(_22302_),
    .B1(_22321_),
    .Y(_22338_));
 sky130_fd_sc_hd__o21bai_4 _25762_ (.A1(_22335_),
    .A2(_22338_),
    .B1_N(_22323_),
    .Y(_22339_));
 sky130_fd_sc_hd__o211a_1 _25763_ (.A1(_22274_),
    .A2(_21740_),
    .B1(_22333_),
    .C1(_22339_),
    .X(_22340_));
 sky130_fd_sc_hd__a21o_1 _25764_ (.A1(_21736_),
    .A2(_21735_),
    .B1(_22274_),
    .X(_22341_));
 sky130_fd_sc_hd__a21oi_4 _25765_ (.A1(_22333_),
    .A2(_22339_),
    .B1(_22341_),
    .Y(_22342_));
 sky130_fd_sc_hd__buf_2 _25766_ (.A(_21736_),
    .X(_22343_));
 sky130_fd_sc_hd__o21ai_4 _25767_ (.A1(_22340_),
    .A2(_22342_),
    .B1(_22343_),
    .Y(_22344_));
 sky130_fd_sc_hd__o21ai_4 _25768_ (.A1(_22274_),
    .A2(_21740_),
    .B1(_22339_),
    .Y(_22345_));
 sky130_fd_sc_hd__inv_2 _25769_ (.A(_22333_),
    .Y(_22346_));
 sky130_fd_sc_hd__inv_2 _25770_ (.A(_21736_),
    .Y(_22348_));
 sky130_fd_sc_hd__a21o_1 _25771_ (.A1(_22333_),
    .A2(_22339_),
    .B1(_22341_),
    .X(_22349_));
 sky130_fd_sc_hd__o211ai_4 _25772_ (.A1(_22345_),
    .A2(_22346_),
    .B1(_22348_),
    .C1(_22349_),
    .Y(_22350_));
 sky130_fd_sc_hd__inv_2 _25773_ (.A(_21746_),
    .Y(_22351_));
 sky130_fd_sc_hd__o221a_1 _25774_ (.A1(_20019_),
    .A2(_20020_),
    .B1(_21737_),
    .B2(_21740_),
    .C1(_20022_),
    .X(_22352_));
 sky130_fd_sc_hd__o21a_2 _25775_ (.A1(_22351_),
    .A2(_22352_),
    .B1(_21744_),
    .X(_22353_));
 sky130_fd_sc_hd__nand3_4 _25776_ (.A(_22344_),
    .B(_22350_),
    .C(_22353_),
    .Y(_22354_));
 sky130_fd_sc_hd__nor2_1 _25777_ (.A(_22351_),
    .B(_22352_),
    .Y(_22355_));
 sky130_fd_sc_hd__o211ai_2 _25778_ (.A1(_22346_),
    .A2(_22345_),
    .B1(_22343_),
    .C1(_22349_),
    .Y(_22356_));
 sky130_fd_sc_hd__o21bai_1 _25779_ (.A1(_22340_),
    .A2(_22342_),
    .B1_N(_22343_),
    .Y(_22357_));
 sky130_fd_sc_hd__o211ai_4 _25780_ (.A1(_21750_),
    .A2(_22355_),
    .B1(_22356_),
    .C1(_22357_),
    .Y(_22359_));
 sky130_fd_sc_hd__xor2_2 _25781_ (.A(_17950_),
    .B(\delay_line[13][9] ),
    .X(_22360_));
 sky130_fd_sc_hd__and3_2 _25782_ (.A(_17956_),
    .B(net396),
    .C(_22360_),
    .X(_22361_));
 sky130_fd_sc_hd__clkbuf_2 _25783_ (.A(net396),
    .X(_22362_));
 sky130_fd_sc_hd__buf_2 _25784_ (.A(_22362_),
    .X(_22363_));
 sky130_fd_sc_hd__a21oi_2 _25785_ (.A1(_17956_),
    .A2(_22363_),
    .B1(_22360_),
    .Y(_22364_));
 sky130_fd_sc_hd__o2bb2ai_1 _25786_ (.A1_N(_22354_),
    .A2_N(_22359_),
    .B1(_22361_),
    .B2(_22364_),
    .Y(_22365_));
 sky130_fd_sc_hd__and2_1 _25787_ (.A(_22360_),
    .B(_21695_),
    .X(_22366_));
 sky130_fd_sc_hd__nor2_1 _25788_ (.A(_21695_),
    .B(_22360_),
    .Y(_22367_));
 sky130_fd_sc_hd__nor2_1 _25789_ (.A(_22366_),
    .B(_22367_),
    .Y(_22368_));
 sky130_fd_sc_hd__a31oi_4 _25790_ (.A1(_22344_),
    .A2(_22350_),
    .A3(_22353_),
    .B1(_22368_),
    .Y(_22370_));
 sky130_fd_sc_hd__nand2_1 _25791_ (.A(_22370_),
    .B(_22359_),
    .Y(_22371_));
 sky130_fd_sc_hd__nand3_2 _25792_ (.A(_22273_),
    .B(_22365_),
    .C(_22371_),
    .Y(_22372_));
 sky130_fd_sc_hd__o2bb2ai_4 _25793_ (.A1_N(_22354_),
    .A2_N(_22359_),
    .B1(_22366_),
    .B2(_22367_),
    .Y(_22373_));
 sky130_fd_sc_hd__o31a_2 _25794_ (.A1(_21697_),
    .A2(_21698_),
    .A3(_21749_),
    .B1(_21756_),
    .X(_22374_));
 sky130_fd_sc_hd__o211ai_4 _25795_ (.A1(_22361_),
    .A2(_22364_),
    .B1(_22354_),
    .C1(_22359_),
    .Y(_22375_));
 sky130_fd_sc_hd__nand3_1 _25796_ (.A(_22373_),
    .B(_22374_),
    .C(_22375_),
    .Y(_22376_));
 sky130_fd_sc_hd__buf_6 _25797_ (.A(_22376_),
    .X(_22377_));
 sky130_fd_sc_hd__xor2_1 _25798_ (.A(_08272_),
    .B(_20046_),
    .X(_22378_));
 sky130_fd_sc_hd__xnor2_1 _25799_ (.A(_21696_),
    .B(_22378_),
    .Y(_22379_));
 sky130_fd_sc_hd__a21oi_2 _25800_ (.A1(_21763_),
    .A2(_21766_),
    .B1(_22379_),
    .Y(_22381_));
 sky130_fd_sc_hd__and3_1 _25801_ (.A(_21763_),
    .B(_21766_),
    .C(_22379_),
    .X(_22382_));
 sky130_fd_sc_hd__or2_2 _25802_ (.A(_22381_),
    .B(_22382_),
    .X(_22383_));
 sky130_fd_sc_hd__a21oi_1 _25803_ (.A1(_22372_),
    .A2(_22377_),
    .B1(_22383_),
    .Y(_22384_));
 sky130_fd_sc_hd__nor2_1 _25804_ (.A(_21775_),
    .B(_21776_),
    .Y(_22385_));
 sky130_fd_sc_hd__a32o_1 _25805_ (.A1(_21693_),
    .A2(_21753_),
    .A3(_21757_),
    .B1(_21777_),
    .B2(_22385_),
    .X(_22386_));
 sky130_fd_sc_hd__a31o_1 _25806_ (.A1(_22372_),
    .A2(_22377_),
    .A3(_22383_),
    .B1(_22386_),
    .X(_22387_));
 sky130_fd_sc_hd__a31o_1 _25807_ (.A1(_19984_),
    .A2(_21766_),
    .A3(_21765_),
    .B1(_21775_),
    .X(_22388_));
 sky130_fd_sc_hd__nand3b_2 _25808_ (.A_N(net403),
    .B(net404),
    .C(net405),
    .Y(_22389_));
 sky130_fd_sc_hd__or2b_1 _25809_ (.A(net405),
    .B_N(net403),
    .X(_22390_));
 sky130_fd_sc_hd__buf_2 _25810_ (.A(_21679_),
    .X(_22392_));
 sky130_fd_sc_hd__and2b_1 _25811_ (.A_N(net404),
    .B(net403),
    .X(_22393_));
 sky130_fd_sc_hd__a311oi_4 _25812_ (.A1(_22389_),
    .A2(_22390_),
    .A3(_22392_),
    .B1(_22393_),
    .C1(_12130_),
    .Y(_22394_));
 sky130_fd_sc_hd__a31oi_1 _25813_ (.A1(_22389_),
    .A2(_22390_),
    .A3(_21679_),
    .B1(_22393_),
    .Y(_22395_));
 sky130_fd_sc_hd__nor2_1 _25814_ (.A(_12141_),
    .B(_22395_),
    .Y(_22396_));
 sky130_fd_sc_hd__clkbuf_2 _25815_ (.A(_22396_),
    .X(_22397_));
 sky130_fd_sc_hd__o21ai_1 _25816_ (.A1(_22394_),
    .A2(_22397_),
    .B1(_08393_),
    .Y(_22398_));
 sky130_fd_sc_hd__or3_1 _25817_ (.A(_25215_),
    .B(_22394_),
    .C(_22397_),
    .X(_22399_));
 sky130_fd_sc_hd__nand3_1 _25818_ (.A(_22388_),
    .B(_22398_),
    .C(_22399_),
    .Y(_22400_));
 sky130_fd_sc_hd__a21o_1 _25819_ (.A1(_22398_),
    .A2(_22399_),
    .B1(_22388_),
    .X(_22401_));
 sky130_fd_sc_hd__nand2_1 _25820_ (.A(_22400_),
    .B(_22401_),
    .Y(_22403_));
 sky130_fd_sc_hd__and2b_1 _25821_ (.A_N(_22403_),
    .B(_21686_),
    .X(_22404_));
 sky130_fd_sc_hd__and4b_1 _25822_ (.A_N(_21684_),
    .B(_08525_),
    .C(_21685_),
    .D(_22403_),
    .X(_22405_));
 sky130_fd_sc_hd__nor2_1 _25823_ (.A(_22404_),
    .B(_22405_),
    .Y(_22406_));
 sky130_fd_sc_hd__inv_2 _25824_ (.A(_22406_),
    .Y(_22407_));
 sky130_fd_sc_hd__o21ai_2 _25825_ (.A1(_22384_),
    .A2(_22387_),
    .B1(_22407_),
    .Y(_22408_));
 sky130_fd_sc_hd__nor2_1 _25826_ (.A(_22381_),
    .B(_22382_),
    .Y(_22409_));
 sky130_fd_sc_hd__nand2_1 _25827_ (.A(_22377_),
    .B(_22409_),
    .Y(_22410_));
 sky130_fd_sc_hd__a21oi_4 _25828_ (.A1(_22375_),
    .A2(_22373_),
    .B1(_22374_),
    .Y(_22411_));
 sky130_fd_sc_hd__o2bb2ai_2 _25829_ (.A1_N(_22372_),
    .A2_N(_22377_),
    .B1(_22381_),
    .B2(_22382_),
    .Y(_22412_));
 sky130_fd_sc_hd__o211a_1 _25830_ (.A1(_22410_),
    .A2(_22411_),
    .B1(_22386_),
    .C1(_22412_),
    .X(_22414_));
 sky130_fd_sc_hd__nor2_1 _25831_ (.A(net170),
    .B(_21789_),
    .Y(_22415_));
 sky130_fd_sc_hd__a32o_2 _25832_ (.A1(_21781_),
    .A2(_21782_),
    .A3(_21783_),
    .B1(_21787_),
    .B2(_22415_),
    .X(_22416_));
 sky130_fd_sc_hd__o211ai_4 _25833_ (.A1(_22410_),
    .A2(_22411_),
    .B1(_22386_),
    .C1(_22412_),
    .Y(_22417_));
 sky130_fd_sc_hd__a21o_1 _25834_ (.A1(_22372_),
    .A2(_22376_),
    .B1(_22383_),
    .X(_22418_));
 sky130_fd_sc_hd__a32oi_2 _25835_ (.A1(_21693_),
    .A2(_21753_),
    .A3(_21757_),
    .B1(_21777_),
    .B2(_22385_),
    .Y(_22419_));
 sky130_fd_sc_hd__o211ai_1 _25836_ (.A1(_22381_),
    .A2(_22382_),
    .B1(_22372_),
    .C1(_22377_),
    .Y(_22420_));
 sky130_fd_sc_hd__nand3_2 _25837_ (.A(_22418_),
    .B(_22419_),
    .C(_22420_),
    .Y(_22421_));
 sky130_fd_sc_hd__or4_1 _25838_ (.A(_20059_),
    .B(_21687_),
    .C(_21684_),
    .D(_22403_),
    .X(_22422_));
 sky130_fd_sc_hd__inv_2 _25839_ (.A(_22422_),
    .Y(_22423_));
 sky130_fd_sc_hd__o31a_1 _25840_ (.A1(_20059_),
    .A2(_21687_),
    .A3(_21684_),
    .B1(_22403_),
    .X(_22425_));
 sky130_fd_sc_hd__o2bb2ai_2 _25841_ (.A1_N(_22417_),
    .A2_N(_22421_),
    .B1(_22423_),
    .B2(_22425_),
    .Y(_22426_));
 sky130_fd_sc_hd__o211ai_4 _25842_ (.A1(_22408_),
    .A2(_22414_),
    .B1(_22416_),
    .C1(_22426_),
    .Y(_22427_));
 sky130_fd_sc_hd__o2bb2ai_1 _25843_ (.A1_N(_22417_),
    .A2_N(_22421_),
    .B1(_22404_),
    .B2(_22405_),
    .Y(_22428_));
 sky130_fd_sc_hd__a21oi_1 _25844_ (.A1(_21787_),
    .A2(_22415_),
    .B1(_21784_),
    .Y(_22429_));
 sky130_fd_sc_hd__o221ai_1 _25845_ (.A1(_22423_),
    .A2(_22425_),
    .B1(_22384_),
    .B2(_22387_),
    .C1(_22417_),
    .Y(_22430_));
 sky130_fd_sc_hd__nand3_1 _25846_ (.A(_22428_),
    .B(_22429_),
    .C(_22430_),
    .Y(_22431_));
 sky130_fd_sc_hd__buf_2 _25847_ (.A(_22431_),
    .X(_22432_));
 sky130_fd_sc_hd__a32o_1 _25848_ (.A1(_19969_),
    .A2(_21804_),
    .A3(_21806_),
    .B1(_21810_),
    .B2(_21827_),
    .X(_22433_));
 sky130_fd_sc_hd__or2b_1 _25849_ (.A(\delay_line[10][1] ),
    .B_N(\delay_line[9][9] ),
    .X(_22434_));
 sky130_fd_sc_hd__inv_2 _25850_ (.A(\delay_line[9][9] ),
    .Y(_22436_));
 sky130_fd_sc_hd__nand2_1 _25851_ (.A(_22436_),
    .B(_25040_),
    .Y(_22437_));
 sky130_fd_sc_hd__a22o_1 _25852_ (.A1(_02821_),
    .A2(_08701_),
    .B1(_22434_),
    .B2(_22437_),
    .X(_22438_));
 sky130_fd_sc_hd__buf_2 _25853_ (.A(net419),
    .X(_22439_));
 sky130_fd_sc_hd__clkbuf_2 _25854_ (.A(_22439_),
    .X(_22440_));
 sky130_fd_sc_hd__nand4_2 _25855_ (.A(_22434_),
    .B(_22437_),
    .C(_02832_),
    .D(_08712_),
    .Y(_22441_));
 sky130_fd_sc_hd__nand4_2 _25856_ (.A(_11691_),
    .B(_22438_),
    .C(_22440_),
    .D(_22441_),
    .Y(_22442_));
 sky130_fd_sc_hd__a22o_1 _25857_ (.A1(_22440_),
    .A2(_11691_),
    .B1(_22438_),
    .B2(_22441_),
    .X(_22443_));
 sky130_fd_sc_hd__or2_1 _25858_ (.A(net413),
    .B(_21817_),
    .X(_22444_));
 sky130_fd_sc_hd__nand2_1 _25859_ (.A(_13042_),
    .B(_08701_),
    .Y(_22445_));
 sky130_fd_sc_hd__clkbuf_2 _25860_ (.A(\delay_line[10][6] ),
    .X(_22447_));
 sky130_fd_sc_hd__clkbuf_2 _25861_ (.A(_22447_),
    .X(_22448_));
 sky130_fd_sc_hd__a21o_1 _25862_ (.A1(_22444_),
    .A2(_22445_),
    .B1(_22448_),
    .X(_22449_));
 sky130_fd_sc_hd__nand3_1 _25863_ (.A(_22444_),
    .B(_22445_),
    .C(_19964_),
    .Y(_22450_));
 sky130_fd_sc_hd__nand3b_2 _25864_ (.A_N(_21823_),
    .B(_22449_),
    .C(_22450_),
    .Y(_22451_));
 sky130_fd_sc_hd__a21bo_1 _25865_ (.A1(_22449_),
    .A2(_22450_),
    .B1_N(_21823_),
    .X(_22452_));
 sky130_fd_sc_hd__nand4_4 _25866_ (.A(_22442_),
    .B(_22443_),
    .C(_22451_),
    .D(_22452_),
    .Y(_22453_));
 sky130_fd_sc_hd__a22o_1 _25867_ (.A1(_22442_),
    .A2(_22443_),
    .B1(_22451_),
    .B2(_22452_),
    .X(_22454_));
 sky130_fd_sc_hd__nand2_1 _25868_ (.A(_21808_),
    .B(_21804_),
    .Y(_22455_));
 sky130_fd_sc_hd__buf_2 _25869_ (.A(\delay_line[10][8] ),
    .X(_22456_));
 sky130_fd_sc_hd__buf_2 _25870_ (.A(_22456_),
    .X(_22458_));
 sky130_fd_sc_hd__nor2_1 _25871_ (.A(net407),
    .B(\delay_line[10][9] ),
    .Y(_22459_));
 sky130_fd_sc_hd__and2_1 _25872_ (.A(\delay_line[12][3] ),
    .B(\delay_line[10][9] ),
    .X(_22460_));
 sky130_fd_sc_hd__or4bb_1 _25873_ (.A(_22459_),
    .B(_22460_),
    .C_N(\delay_line[12][2] ),
    .D_N(\delay_line[10][8] ),
    .X(_22461_));
 sky130_fd_sc_hd__a2bb2o_1 _25874_ (.A1_N(_22459_),
    .A2_N(_22460_),
    .B1(\delay_line[12][2] ),
    .B2(\delay_line[10][8] ),
    .X(_22462_));
 sky130_fd_sc_hd__nand2_1 _25875_ (.A(_22461_),
    .B(_22462_),
    .Y(_22463_));
 sky130_fd_sc_hd__a21o_1 _25876_ (.A1(_21680_),
    .A2(_21685_),
    .B1(_22463_),
    .X(_22464_));
 sky130_fd_sc_hd__buf_2 _25877_ (.A(_22392_),
    .X(_22465_));
 sky130_fd_sc_hd__o211ai_1 _25878_ (.A1(_22465_),
    .A2(_20061_),
    .B1(_21685_),
    .C1(_22463_),
    .Y(_22466_));
 sky130_fd_sc_hd__a2bb2o_1 _25879_ (.A1_N(_13031_),
    .A2_N(_22458_),
    .B1(_22464_),
    .B2(_22466_),
    .X(_22467_));
 sky130_fd_sc_hd__nor2_1 _25880_ (.A(_22456_),
    .B(_13031_),
    .Y(_22469_));
 sky130_fd_sc_hd__nand3_1 _25881_ (.A(_22466_),
    .B(_22464_),
    .C(_22469_),
    .Y(_22470_));
 sky130_fd_sc_hd__clkbuf_2 _25882_ (.A(_22470_),
    .X(_22471_));
 sky130_fd_sc_hd__nand4_2 _25883_ (.A(_21806_),
    .B(_22455_),
    .C(_22467_),
    .D(_22471_),
    .Y(_22472_));
 sky130_fd_sc_hd__a22o_1 _25884_ (.A1(_21806_),
    .A2(_22455_),
    .B1(_22467_),
    .B2(_22471_),
    .X(_22473_));
 sky130_fd_sc_hd__a22o_1 _25885_ (.A1(_22453_),
    .A2(_22454_),
    .B1(_22472_),
    .B2(_22473_),
    .X(_22474_));
 sky130_fd_sc_hd__a22oi_2 _25886_ (.A1(_21806_),
    .A2(_22455_),
    .B1(_22467_),
    .B2(_22471_),
    .Y(_22475_));
 sky130_fd_sc_hd__nand2_1 _25887_ (.A(_22453_),
    .B(_22454_),
    .Y(_22476_));
 sky130_fd_sc_hd__or3b_1 _25888_ (.A(_22475_),
    .B(_22476_),
    .C_N(_22472_),
    .X(_22477_));
 sky130_fd_sc_hd__nand2_1 _25889_ (.A(_22474_),
    .B(_22477_),
    .Y(_22478_));
 sky130_fd_sc_hd__a31o_1 _25890_ (.A1(_20052_),
    .A2(_21686_),
    .A3(_21688_),
    .B1(_21788_),
    .X(_22480_));
 sky130_fd_sc_hd__and2b_1 _25891_ (.A_N(_22478_),
    .B(_22480_),
    .X(_22481_));
 sky130_fd_sc_hd__and2b_1 _25892_ (.A_N(_22480_),
    .B(_22478_),
    .X(_22482_));
 sky130_fd_sc_hd__nor2_1 _25893_ (.A(_22481_),
    .B(_22482_),
    .Y(_22483_));
 sky130_fd_sc_hd__inv_2 _25894_ (.A(_22483_),
    .Y(_22484_));
 sky130_fd_sc_hd__nor2_1 _25895_ (.A(_22433_),
    .B(_22484_),
    .Y(_22485_));
 sky130_fd_sc_hd__and2_1 _25896_ (.A(_22433_),
    .B(_22484_),
    .X(_22486_));
 sky130_fd_sc_hd__o2bb2ai_1 _25897_ (.A1_N(_22427_),
    .A2_N(_22432_),
    .B1(_22485_),
    .B2(_22486_),
    .Y(_22487_));
 sky130_fd_sc_hd__a21o_2 _25898_ (.A1(_21795_),
    .A2(_21892_),
    .B1(_21894_),
    .X(_22488_));
 sky130_fd_sc_hd__inv_2 _25899_ (.A(_22488_),
    .Y(_22489_));
 sky130_fd_sc_hd__and2_2 _25900_ (.A(_22483_),
    .B(_22433_),
    .X(_22491_));
 sky130_fd_sc_hd__nor2_2 _25901_ (.A(_22433_),
    .B(_22483_),
    .Y(_22492_));
 sky130_fd_sc_hd__o211ai_4 _25902_ (.A1(_22491_),
    .A2(_22492_),
    .B1(_22427_),
    .C1(_22432_),
    .Y(_22493_));
 sky130_fd_sc_hd__nand3_4 _25903_ (.A(_22487_),
    .B(_22489_),
    .C(_22493_),
    .Y(_22494_));
 sky130_fd_sc_hd__nor2_1 _25904_ (.A(_22491_),
    .B(_22492_),
    .Y(_22495_));
 sky130_fd_sc_hd__nand2_1 _25905_ (.A(_22432_),
    .B(_22495_),
    .Y(_22496_));
 sky130_fd_sc_hd__o211a_2 _25906_ (.A1(_22408_),
    .A2(_22414_),
    .B1(_22416_),
    .C1(_22426_),
    .X(_22497_));
 sky130_fd_sc_hd__o2bb2ai_2 _25907_ (.A1_N(_22427_),
    .A2_N(_22432_),
    .B1(_22491_),
    .B2(_22492_),
    .Y(_22498_));
 sky130_fd_sc_hd__o211ai_4 _25908_ (.A1(_22496_),
    .A2(_22497_),
    .B1(_22488_),
    .C1(_22498_),
    .Y(_22499_));
 sky130_fd_sc_hd__and2b_1 _25909_ (.A_N(\delay_line[9][1] ),
    .B(\delay_line[8][9] ),
    .X(_22500_));
 sky130_fd_sc_hd__buf_1 _25910_ (.A(_22500_),
    .X(_22502_));
 sky130_fd_sc_hd__buf_1 _25911_ (.A(\delay_line[8][9] ),
    .X(_22503_));
 sky130_fd_sc_hd__and2b_1 _25912_ (.A_N(_22503_),
    .B(\delay_line[9][1] ),
    .X(_22504_));
 sky130_fd_sc_hd__or3_1 _25913_ (.A(_22502_),
    .B(_22504_),
    .C(_21868_),
    .X(_22505_));
 sky130_fd_sc_hd__o21ai_1 _25914_ (.A1(_22502_),
    .A2(_22504_),
    .B1(_21868_),
    .Y(_22506_));
 sky130_fd_sc_hd__o21ai_2 _25915_ (.A1(_20104_),
    .A2(net424),
    .B1(_20099_),
    .Y(_22507_));
 sky130_fd_sc_hd__and2_1 _25916_ (.A(_20104_),
    .B(net424),
    .X(_22508_));
 sky130_fd_sc_hd__clkbuf_2 _25917_ (.A(_20104_),
    .X(_22509_));
 sky130_fd_sc_hd__nor2_1 _25918_ (.A(_22509_),
    .B(_21867_),
    .Y(_22510_));
 sky130_fd_sc_hd__o21bai_2 _25919_ (.A1(_22508_),
    .A2(_22510_),
    .B1_N(_20099_),
    .Y(_22511_));
 sky130_fd_sc_hd__o211ai_4 _25920_ (.A1(_22507_),
    .A2(_22508_),
    .B1(_20103_),
    .C1(_22511_),
    .Y(_22513_));
 sky130_fd_sc_hd__a21o_1 _25921_ (.A1(_22509_),
    .A2(_21867_),
    .B1(_22507_),
    .X(_22514_));
 sky130_fd_sc_hd__a21o_1 _25922_ (.A1(_22514_),
    .A2(_22511_),
    .B1(_20103_),
    .X(_22515_));
 sky130_fd_sc_hd__a21o_1 _25923_ (.A1(_22513_),
    .A2(_22515_),
    .B1(_09020_),
    .X(_22516_));
 sky130_fd_sc_hd__nand3_2 _25924_ (.A(_22515_),
    .B(_09020_),
    .C(_22513_),
    .Y(_22517_));
 sky130_fd_sc_hd__a22oi_2 _25925_ (.A1(_22505_),
    .A2(_22506_),
    .B1(_22516_),
    .B2(_22517_),
    .Y(_22518_));
 sky130_fd_sc_hd__and4_1 _25926_ (.A(_22505_),
    .B(_22506_),
    .C(_22516_),
    .D(_22517_),
    .X(_22519_));
 sky130_fd_sc_hd__or3b_1 _25927_ (.A(_22518_),
    .B(_22519_),
    .C_N(_21875_),
    .X(_22520_));
 sky130_fd_sc_hd__o21bai_1 _25928_ (.A1(_22518_),
    .A2(_22519_),
    .B1_N(_21875_),
    .Y(_22521_));
 sky130_fd_sc_hd__and2_1 _25929_ (.A(_20105_),
    .B(_21872_),
    .X(_22522_));
 sky130_fd_sc_hd__or2b_1 _25930_ (.A(_03150_),
    .B_N(net425),
    .X(_22524_));
 sky130_fd_sc_hd__clkbuf_2 _25931_ (.A(net425),
    .X(_22525_));
 sky130_fd_sc_hd__or2b_1 _25932_ (.A(_22525_),
    .B_N(_03161_),
    .X(_22526_));
 sky130_fd_sc_hd__clkbuf_2 _25933_ (.A(\delay_line[7][8] ),
    .X(_22527_));
 sky130_fd_sc_hd__nand4_2 _25934_ (.A(_22996_),
    .B(_22524_),
    .C(_22526_),
    .D(_22527_),
    .Y(_22528_));
 sky130_fd_sc_hd__a22o_1 _25935_ (.A1(_22996_),
    .A2(_22527_),
    .B1(_22524_),
    .B2(_22526_),
    .X(_22529_));
 sky130_fd_sc_hd__nand2_1 _25936_ (.A(_22528_),
    .B(_22529_),
    .Y(_22530_));
 sky130_fd_sc_hd__xnor2_1 _25937_ (.A(_22522_),
    .B(_22530_),
    .Y(_22531_));
 sky130_fd_sc_hd__a21oi_1 _25938_ (.A1(_22520_),
    .A2(_22521_),
    .B1(_22531_),
    .Y(_22532_));
 sky130_fd_sc_hd__nand3_1 _25939_ (.A(_22531_),
    .B(_22520_),
    .C(_22521_),
    .Y(_22533_));
 sky130_fd_sc_hd__and2b_2 _25940_ (.A_N(_22532_),
    .B(_22533_),
    .X(_22535_));
 sky130_fd_sc_hd__o211ai_1 _25941_ (.A1(_18869_),
    .A2(_18870_),
    .B1(_18052_),
    .C1(_11669_),
    .Y(_22536_));
 sky130_fd_sc_hd__nor2_1 _25942_ (.A(_21853_),
    .B(net207),
    .Y(_22537_));
 sky130_fd_sc_hd__and4b_1 _25943_ (.A_N(_22536_),
    .B(_22537_),
    .C(_20133_),
    .D(_20131_),
    .X(_22538_));
 sky130_fd_sc_hd__a41o_1 _25944_ (.A1(_25062_),
    .A2(_08723_),
    .A3(_21845_),
    .A4(_21846_),
    .B1(_21850_),
    .X(_22539_));
 sky130_fd_sc_hd__o21ai_2 _25945_ (.A1(_21816_),
    .A2(_21826_),
    .B1(_21824_),
    .Y(_22540_));
 sky130_fd_sc_hd__inv_2 _25946_ (.A(net421),
    .Y(_22541_));
 sky130_fd_sc_hd__a21o_1 _25947_ (.A1(_22541_),
    .A2(_21843_),
    .B1(net419),
    .X(_22542_));
 sky130_fd_sc_hd__buf_2 _25948_ (.A(_22541_),
    .X(_22543_));
 sky130_fd_sc_hd__nand3_1 _25949_ (.A(_22543_),
    .B(_21843_),
    .C(_22439_),
    .Y(_22544_));
 sky130_fd_sc_hd__nand3_1 _25950_ (.A(_22542_),
    .B(_22544_),
    .C(_08657_),
    .Y(_22546_));
 sky130_fd_sc_hd__a21oi_1 _25951_ (.A1(_22543_),
    .A2(_21843_),
    .B1(_22439_),
    .Y(_22547_));
 sky130_fd_sc_hd__and3_1 _25952_ (.A(_22541_),
    .B(_20125_),
    .C(net419),
    .X(_22548_));
 sky130_fd_sc_hd__o21bai_2 _25953_ (.A1(_22547_),
    .A2(_22548_),
    .B1_N(_08657_),
    .Y(_22549_));
 sky130_fd_sc_hd__a21bo_1 _25954_ (.A1(_22546_),
    .A2(_22549_),
    .B1_N(_21814_),
    .X(_22550_));
 sky130_fd_sc_hd__nand3b_2 _25955_ (.A_N(_21814_),
    .B(_22546_),
    .C(_22549_),
    .Y(_22551_));
 sky130_fd_sc_hd__o2111ai_4 _25956_ (.A1(_20128_),
    .A2(_21844_),
    .B1(_21845_),
    .C1(_22550_),
    .D1(_22551_),
    .Y(_22552_));
 sky130_fd_sc_hd__a22o_1 _25957_ (.A1(_20127_),
    .A2(_21845_),
    .B1(_22550_),
    .B2(_22551_),
    .X(_22553_));
 sky130_fd_sc_hd__and3_1 _25958_ (.A(_22540_),
    .B(_22552_),
    .C(_22553_),
    .X(_22554_));
 sky130_fd_sc_hd__a21oi_1 _25959_ (.A1(_22552_),
    .A2(_22553_),
    .B1(_22540_),
    .Y(_22555_));
 sky130_fd_sc_hd__nor2_1 _25960_ (.A(_22554_),
    .B(_22555_),
    .Y(_22557_));
 sky130_fd_sc_hd__xnor2_1 _25961_ (.A(_22539_),
    .B(_22557_),
    .Y(_22558_));
 sky130_fd_sc_hd__o21bai_2 _25962_ (.A1(_21854_),
    .A2(_22538_),
    .B1_N(_22558_),
    .Y(_22559_));
 sky130_fd_sc_hd__o311a_1 _25963_ (.A1(_21852_),
    .A2(_21850_),
    .A3(_21851_),
    .B1(_21855_),
    .C1(_22558_),
    .X(_22560_));
 sky130_fd_sc_hd__inv_2 _25964_ (.A(_22560_),
    .Y(_22561_));
 sky130_fd_sc_hd__nand2_1 _25965_ (.A(_22559_),
    .B(_22561_),
    .Y(_22562_));
 sky130_fd_sc_hd__xnor2_1 _25966_ (.A(_22535_),
    .B(_22562_),
    .Y(_22563_));
 sky130_fd_sc_hd__o21ai_1 _25967_ (.A1(_21798_),
    .A2(_21828_),
    .B1(_21835_),
    .Y(_22564_));
 sky130_fd_sc_hd__nand2_1 _25968_ (.A(_22563_),
    .B(_22564_),
    .Y(_22565_));
 sky130_fd_sc_hd__and2_1 _25969_ (.A(_22535_),
    .B(_22562_),
    .X(_22566_));
 sky130_fd_sc_hd__or3b_1 _25970_ (.A(_22560_),
    .B(_22535_),
    .C_N(_22559_),
    .X(_22568_));
 sky130_fd_sc_hd__or3b_2 _25971_ (.A(_22564_),
    .B(_22566_),
    .C_N(_22568_),
    .X(_22569_));
 sky130_fd_sc_hd__a21o_1 _25972_ (.A1(_21859_),
    .A2(_21881_),
    .B1(_21857_),
    .X(_22570_));
 sky130_fd_sc_hd__a21oi_2 _25973_ (.A1(_22565_),
    .A2(_22569_),
    .B1(_22570_),
    .Y(_22571_));
 sky130_fd_sc_hd__and3_1 _25974_ (.A(_22570_),
    .B(_22565_),
    .C(_22569_),
    .X(_22572_));
 sky130_fd_sc_hd__o2bb2ai_1 _25975_ (.A1_N(_22494_),
    .A2_N(_22499_),
    .B1(_22571_),
    .B2(_22572_),
    .Y(_22573_));
 sky130_fd_sc_hd__inv_2 _25976_ (.A(_22570_),
    .Y(_22574_));
 sky130_fd_sc_hd__a21oi_2 _25977_ (.A1(_22565_),
    .A2(_22569_),
    .B1(_22574_),
    .Y(_22575_));
 sky130_fd_sc_hd__and3_1 _25978_ (.A(_22569_),
    .B(_22574_),
    .C(_22565_),
    .X(_22576_));
 sky130_fd_sc_hd__o211ai_2 _25979_ (.A1(_22575_),
    .A2(_22576_),
    .B1(_22494_),
    .C1(_22499_),
    .Y(_22577_));
 sky130_fd_sc_hd__a21oi_2 _25980_ (.A1(_21840_),
    .A2(_21890_),
    .B1(_21896_),
    .Y(_22579_));
 sky130_fd_sc_hd__nand3_4 _25981_ (.A(_22573_),
    .B(_22577_),
    .C(_22579_),
    .Y(_22580_));
 sky130_fd_sc_hd__o2bb2ai_2 _25982_ (.A1_N(_22494_),
    .A2_N(_22499_),
    .B1(_22575_),
    .B2(_22576_),
    .Y(_22581_));
 sky130_fd_sc_hd__o211ai_4 _25983_ (.A1(_22571_),
    .A2(_22572_),
    .B1(_22494_),
    .C1(_22499_),
    .Y(_22582_));
 sky130_fd_sc_hd__a21o_1 _25984_ (.A1(_21840_),
    .A2(_21890_),
    .B1(_21896_),
    .X(_22583_));
 sky130_fd_sc_hd__nand3_2 _25985_ (.A(_22581_),
    .B(_22582_),
    .C(_22583_),
    .Y(_22584_));
 sky130_fd_sc_hd__a21bo_1 _25986_ (.A1(_21937_),
    .A2(_22001_),
    .B1_N(_21935_),
    .X(_22585_));
 sky130_fd_sc_hd__nor2_1 _25987_ (.A(_21887_),
    .B(_21885_),
    .Y(_22586_));
 sky130_fd_sc_hd__a31o_1 _25988_ (.A1(_20091_),
    .A2(_21883_),
    .A3(_21884_),
    .B1(_22586_),
    .X(_22587_));
 sky130_fd_sc_hd__a21o_1 _25989_ (.A1(_20114_),
    .A2(_20118_),
    .B1(_21930_),
    .X(_22588_));
 sky130_fd_sc_hd__a21o_1 _25990_ (.A1(_21915_),
    .A2(_21920_),
    .B1(_21914_),
    .X(_22590_));
 sky130_fd_sc_hd__buf_2 _25991_ (.A(_21911_),
    .X(_22591_));
 sky130_fd_sc_hd__nor2_1 _25992_ (.A(_11954_),
    .B(\delay_line[7][5] ),
    .Y(_22592_));
 sky130_fd_sc_hd__nand2_1 _25993_ (.A(_11954_),
    .B(_18025_),
    .Y(_22593_));
 sky130_fd_sc_hd__or2b_1 _25994_ (.A(_22592_),
    .B_N(_22593_),
    .X(_22594_));
 sky130_fd_sc_hd__xor2_1 _25995_ (.A(_22591_),
    .B(_22594_),
    .X(_22595_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _25996_ (.A(\delay_line[6][9] ),
    .X(_22596_));
 sky130_fd_sc_hd__nand2_1 _25997_ (.A(_00051_),
    .B(_22596_),
    .Y(_22597_));
 sky130_fd_sc_hd__or2_1 _25998_ (.A(_00051_),
    .B(\delay_line[6][9] ),
    .X(_22598_));
 sky130_fd_sc_hd__nand4_2 _25999_ (.A(_21909_),
    .B(_21907_),
    .C(_22597_),
    .D(_22598_),
    .Y(_22599_));
 sky130_fd_sc_hd__and2_1 _26000_ (.A(\delay_line[7][1] ),
    .B(\delay_line[6][9] ),
    .X(_22601_));
 sky130_fd_sc_hd__nor2_1 _26001_ (.A(_00051_),
    .B(_22596_),
    .Y(_22602_));
 sky130_fd_sc_hd__o2bb2ai_4 _26002_ (.A1_N(_21909_),
    .A2_N(_21907_),
    .B1(_22601_),
    .B2(_22602_),
    .Y(_22603_));
 sky130_fd_sc_hd__buf_2 _26003_ (.A(\delay_line[6][8] ),
    .X(_22604_));
 sky130_fd_sc_hd__nand4_4 _26004_ (.A(_22974_),
    .B(_22599_),
    .C(_22603_),
    .D(_22604_),
    .Y(_22605_));
 sky130_fd_sc_hd__clkbuf_2 _26005_ (.A(\delay_line[6][8] ),
    .X(_22606_));
 sky130_fd_sc_hd__a22o_1 _26006_ (.A1(_22963_),
    .A2(_22606_),
    .B1(_22599_),
    .B2(_22603_),
    .X(_22607_));
 sky130_fd_sc_hd__and3_1 _26007_ (.A(_22595_),
    .B(_22605_),
    .C(_22607_),
    .X(_22608_));
 sky130_fd_sc_hd__a21oi_1 _26008_ (.A1(_22605_),
    .A2(_22607_),
    .B1(_22595_),
    .Y(_22609_));
 sky130_fd_sc_hd__o211ai_1 _26009_ (.A1(_22608_),
    .A2(_22609_),
    .B1(_21863_),
    .C1(_21861_),
    .Y(_22610_));
 sky130_fd_sc_hd__a211o_1 _26010_ (.A1(_21861_),
    .A2(_21863_),
    .B1(_22609_),
    .C1(_22608_),
    .X(_22612_));
 sky130_fd_sc_hd__nand3b_1 _26011_ (.A_N(_22590_),
    .B(_22610_),
    .C(_22612_),
    .Y(_22613_));
 sky130_fd_sc_hd__a21bo_1 _26012_ (.A1(_22610_),
    .A2(_22612_),
    .B1_N(_22590_),
    .X(_22614_));
 sky130_fd_sc_hd__o21ai_1 _26013_ (.A1(_21875_),
    .A2(_21876_),
    .B1(_21877_),
    .Y(_22615_));
 sky130_fd_sc_hd__a21oi_1 _26014_ (.A1(_22615_),
    .A2(_21866_),
    .B1(_21879_),
    .Y(_22616_));
 sky130_fd_sc_hd__a21boi_1 _26015_ (.A1(_22613_),
    .A2(_22614_),
    .B1_N(_22616_),
    .Y(_22617_));
 sky130_fd_sc_hd__nand3b_2 _26016_ (.A_N(_22616_),
    .B(_22613_),
    .C(_22614_),
    .Y(_22618_));
 sky130_fd_sc_hd__nand3_1 _26017_ (.A(_21928_),
    .B(_21929_),
    .C(_22618_),
    .Y(_22619_));
 sky130_fd_sc_hd__a21bo_1 _26018_ (.A1(_22613_),
    .A2(_22614_),
    .B1_N(_22616_),
    .X(_22620_));
 sky130_fd_sc_hd__a22o_1 _26019_ (.A1(_21928_),
    .A2(_21929_),
    .B1(_22620_),
    .B2(_22618_),
    .X(_22621_));
 sky130_fd_sc_hd__o21a_1 _26020_ (.A1(_22617_),
    .A2(_22619_),
    .B1(_22621_),
    .X(_22623_));
 sky130_fd_sc_hd__a21o_1 _26021_ (.A1(_22588_),
    .A2(_21934_),
    .B1(_22623_),
    .X(_22624_));
 sky130_fd_sc_hd__inv_2 _26022_ (.A(_22624_),
    .Y(_22625_));
 sky130_fd_sc_hd__and3_1 _26023_ (.A(_22623_),
    .B(_21934_),
    .C(_22588_),
    .X(_22626_));
 sky130_fd_sc_hd__and2_1 _26024_ (.A(_21978_),
    .B(_19904_),
    .X(_22627_));
 sky130_fd_sc_hd__nor2_1 _26025_ (.A(_21978_),
    .B(_21979_),
    .Y(_22628_));
 sky130_fd_sc_hd__o21bai_2 _26026_ (.A1(_22627_),
    .A2(_22628_),
    .B1_N(_18080_),
    .Y(_22629_));
 sky130_fd_sc_hd__a21o_1 _26027_ (.A1(_19905_),
    .A2(_22629_),
    .B1(net273),
    .X(_22630_));
 sky130_fd_sc_hd__nand3_1 _26028_ (.A(net273),
    .B(_22629_),
    .C(_19905_),
    .Y(_22631_));
 sky130_fd_sc_hd__a21bo_1 _26029_ (.A1(_21983_),
    .A2(_21956_),
    .B1_N(_21980_),
    .X(_22632_));
 sky130_fd_sc_hd__a21oi_1 _26030_ (.A1(_22630_),
    .A2(_22631_),
    .B1(_22632_),
    .Y(_22634_));
 sky130_fd_sc_hd__and3_1 _26031_ (.A(_22632_),
    .B(_22630_),
    .C(_22631_),
    .X(_22635_));
 sky130_fd_sc_hd__a211o_1 _26032_ (.A1(_21986_),
    .A2(_21988_),
    .B1(_22634_),
    .C1(_22635_),
    .X(_22636_));
 sky130_fd_sc_hd__o211ai_2 _26033_ (.A1(_22634_),
    .A2(_22635_),
    .B1(_21986_),
    .C1(_21988_),
    .Y(_22637_));
 sky130_fd_sc_hd__inv_2 _26034_ (.A(\delay_line[3][9] ),
    .Y(_22638_));
 sky130_fd_sc_hd__nor2_1 _26035_ (.A(_18101_),
    .B(_22638_),
    .Y(_22639_));
 sky130_fd_sc_hd__clkbuf_2 _26036_ (.A(_22638_),
    .X(_22640_));
 sky130_fd_sc_hd__and2_1 _26037_ (.A(_22640_),
    .B(_18098_),
    .X(_22641_));
 sky130_fd_sc_hd__buf_2 _26038_ (.A(_19927_),
    .X(_22642_));
 sky130_fd_sc_hd__clkbuf_2 _26039_ (.A(_22642_),
    .X(_22643_));
 sky130_fd_sc_hd__o21ai_1 _26040_ (.A1(_22639_),
    .A2(_22641_),
    .B1(_22643_),
    .Y(_22645_));
 sky130_fd_sc_hd__or3_1 _26041_ (.A(_22643_),
    .B(_22639_),
    .C(_22641_),
    .X(_22646_));
 sky130_fd_sc_hd__and3_1 _26042_ (.A(_21961_),
    .B(_21963_),
    .C(\delay_line[5][7] ),
    .X(_22647_));
 sky130_fd_sc_hd__nand2b_1 _26043_ (.A_N(_19062_),
    .B(\delay_line[5][9] ),
    .Y(_22648_));
 sky130_fd_sc_hd__or2b_1 _26044_ (.A(\delay_line[5][9] ),
    .B_N(_19062_),
    .X(_22649_));
 sky130_fd_sc_hd__nand3_1 _26045_ (.A(_22648_),
    .B(_22649_),
    .C(_21958_),
    .Y(_22650_));
 sky130_fd_sc_hd__buf_2 _26046_ (.A(_22650_),
    .X(_22651_));
 sky130_fd_sc_hd__a21o_2 _26047_ (.A1(_22648_),
    .A2(_22649_),
    .B1(_21958_),
    .X(_22652_));
 sky130_fd_sc_hd__o211ai_4 _26048_ (.A1(_21957_),
    .A2(_22647_),
    .B1(_22651_),
    .C1(_22652_),
    .Y(_22653_));
 sky130_fd_sc_hd__o21ai_2 _26049_ (.A1(_19927_),
    .A2(_21959_),
    .B1(_21961_),
    .Y(_22654_));
 sky130_fd_sc_hd__a21o_1 _26050_ (.A1(_22651_),
    .A2(_22652_),
    .B1(_22654_),
    .X(_22656_));
 sky130_fd_sc_hd__o2111ai_4 _26051_ (.A1(_19928_),
    .A2(_21969_),
    .B1(_22653_),
    .C1(_22656_),
    .D1(_21965_),
    .Y(_22657_));
 sky130_fd_sc_hd__o21a_1 _26052_ (.A1(_22919_),
    .A2(_22642_),
    .B1(_21966_),
    .X(_22658_));
 sky130_fd_sc_hd__nand2_1 _26053_ (.A(_22653_),
    .B(_22656_),
    .Y(_22659_));
 sky130_fd_sc_hd__o21ai_1 _26054_ (.A1(_21968_),
    .A2(_22658_),
    .B1(_22659_),
    .Y(_22660_));
 sky130_fd_sc_hd__nand4_2 _26055_ (.A(_22645_),
    .B(_22646_),
    .C(_22657_),
    .D(_22660_),
    .Y(_22661_));
 sky130_fd_sc_hd__a22o_1 _26056_ (.A1(_22645_),
    .A2(_22646_),
    .B1(_22657_),
    .B2(_22660_),
    .X(_22662_));
 sky130_fd_sc_hd__nand2_1 _26057_ (.A(_22661_),
    .B(_22662_),
    .Y(_22663_));
 sky130_fd_sc_hd__a21o_1 _26058_ (.A1(_22636_),
    .A2(_22637_),
    .B1(_22663_),
    .X(_22664_));
 sky130_fd_sc_hd__nand3_1 _26059_ (.A(_22663_),
    .B(_22636_),
    .C(_22637_),
    .Y(_22665_));
 sky130_fd_sc_hd__a22o_1 _26060_ (.A1(_21993_),
    .A2(_21994_),
    .B1(_22664_),
    .B2(_22665_),
    .X(_22667_));
 sky130_fd_sc_hd__nand4_1 _26061_ (.A(_21993_),
    .B(_21994_),
    .C(_22664_),
    .D(_22665_),
    .Y(_22668_));
 sky130_fd_sc_hd__nand2_1 _26062_ (.A(_22667_),
    .B(_22668_),
    .Y(_22669_));
 sky130_fd_sc_hd__nand2_1 _26063_ (.A(_21945_),
    .B(_21947_),
    .Y(_22670_));
 sky130_fd_sc_hd__or2b_1 _26064_ (.A(_19885_),
    .B_N(net441),
    .X(_22671_));
 sky130_fd_sc_hd__or2b_1 _26065_ (.A(net441),
    .B_N(_19885_),
    .X(_22672_));
 sky130_fd_sc_hd__nand4_2 _26066_ (.A(_03568_),
    .B(_22671_),
    .C(_22672_),
    .D(_21971_),
    .Y(_22673_));
 sky130_fd_sc_hd__inv_2 _26067_ (.A(\delay_line[3][8] ),
    .Y(_22674_));
 sky130_fd_sc_hd__o2bb2ai_1 _26068_ (.A1_N(_22671_),
    .A2_N(_22672_),
    .B1(_03546_),
    .B2(_22674_),
    .Y(_22675_));
 sky130_fd_sc_hd__and2b_1 _26069_ (.A_N(_19047_),
    .B(net442),
    .X(_22676_));
 sky130_fd_sc_hd__a21oi_2 _26070_ (.A1(_22673_),
    .A2(_22675_),
    .B1(_22676_),
    .Y(_22678_));
 sky130_fd_sc_hd__o21ai_2 _26071_ (.A1(_18104_),
    .A2(_21972_),
    .B1(_19882_),
    .Y(_22679_));
 sky130_fd_sc_hd__a31oi_1 _26072_ (.A1(_22676_),
    .A2(_22673_),
    .A3(_22675_),
    .B1(_22679_),
    .Y(_22680_));
 sky130_fd_sc_hd__or2b_1 _26073_ (.A(_22678_),
    .B_N(_22680_),
    .X(_22681_));
 sky130_fd_sc_hd__and3_1 _26074_ (.A(_22675_),
    .B(_22676_),
    .C(_22673_),
    .X(_22682_));
 sky130_fd_sc_hd__o21ai_1 _26075_ (.A1(_22678_),
    .A2(_22682_),
    .B1(_22679_),
    .Y(_22683_));
 sky130_fd_sc_hd__nand3b_4 _26076_ (.A_N(_21942_),
    .B(_22681_),
    .C(_22683_),
    .Y(_22684_));
 sky130_fd_sc_hd__nor3_1 _26077_ (.A(_22679_),
    .B(_22678_),
    .C(_22682_),
    .Y(_22685_));
 sky130_fd_sc_hd__o21a_1 _26078_ (.A1(_22678_),
    .A2(_22682_),
    .B1(_22679_),
    .X(_22686_));
 sky130_fd_sc_hd__o21ai_2 _26079_ (.A1(_22685_),
    .A2(_22686_),
    .B1(_21942_),
    .Y(_22687_));
 sky130_fd_sc_hd__and3_1 _26080_ (.A(_21965_),
    .B(_21966_),
    .C(_19930_),
    .X(_22689_));
 sky130_fd_sc_hd__a21oi_2 _26081_ (.A1(_21967_),
    .A2(_21970_),
    .B1(_21973_),
    .Y(_22690_));
 sky130_fd_sc_hd__a211o_1 _26082_ (.A1(_22684_),
    .A2(_22687_),
    .B1(_22689_),
    .C1(_22690_),
    .X(_22691_));
 sky130_fd_sc_hd__o211ai_4 _26083_ (.A1(_22690_),
    .A2(_22689_),
    .B1(_22687_),
    .C1(_22684_),
    .Y(_22692_));
 sky130_fd_sc_hd__and3_1 _26084_ (.A(_22670_),
    .B(_22691_),
    .C(_22692_),
    .X(_22693_));
 sky130_fd_sc_hd__a21oi_1 _26085_ (.A1(_22691_),
    .A2(_22692_),
    .B1(_22670_),
    .Y(_22694_));
 sky130_fd_sc_hd__nor2_1 _26086_ (.A(_22693_),
    .B(_22694_),
    .Y(_22695_));
 sky130_fd_sc_hd__xor2_2 _26087_ (.A(_22669_),
    .B(_22695_),
    .X(_22696_));
 sky130_fd_sc_hd__o21a_1 _26088_ (.A1(_22625_),
    .A2(_22626_),
    .B1(_22696_),
    .X(_22697_));
 sky130_fd_sc_hd__inv_2 _26089_ (.A(_22697_),
    .Y(_22698_));
 sky130_fd_sc_hd__or3_2 _26090_ (.A(_22696_),
    .B(_22626_),
    .C(_22625_),
    .X(_22700_));
 sky130_fd_sc_hd__nand3_2 _26091_ (.A(_22587_),
    .B(_22698_),
    .C(_22700_),
    .Y(_22701_));
 sky130_fd_sc_hd__a21o_1 _26092_ (.A1(_22698_),
    .A2(_22700_),
    .B1(_22587_),
    .X(_22702_));
 sky130_fd_sc_hd__and3_1 _26093_ (.A(_22585_),
    .B(_22701_),
    .C(_22702_),
    .X(_22703_));
 sky130_fd_sc_hd__a21oi_2 _26094_ (.A1(_22701_),
    .A2(_22702_),
    .B1(_22585_),
    .Y(_22704_));
 sky130_fd_sc_hd__nor2_2 _26095_ (.A(_22703_),
    .B(_22704_),
    .Y(_22705_));
 sky130_fd_sc_hd__nand3_2 _26096_ (.A(_22580_),
    .B(_22584_),
    .C(_22705_),
    .Y(_22706_));
 sky130_fd_sc_hd__o2bb2ai_4 _26097_ (.A1_N(_22580_),
    .A2_N(_22584_),
    .B1(_22703_),
    .B2(_22704_),
    .Y(_22707_));
 sky130_fd_sc_hd__o211a_1 _26098_ (.A1(_22271_),
    .A2(_22272_),
    .B1(_22706_),
    .C1(_22707_),
    .X(_22708_));
 sky130_fd_sc_hd__o21ai_1 _26099_ (.A1(_22018_),
    .A2(_22017_),
    .B1(_22012_),
    .Y(_22709_));
 sky130_fd_sc_hd__a21oi_1 _26100_ (.A1(_22706_),
    .A2(_22707_),
    .B1(_22709_),
    .Y(_22711_));
 sky130_fd_sc_hd__o22ai_1 _26101_ (.A1(_22268_),
    .A2(_22269_),
    .B1(_22708_),
    .B2(_22711_),
    .Y(_22712_));
 sky130_fd_sc_hd__o21ai_2 _26102_ (.A1(_22016_),
    .A2(_22066_),
    .B1(_22072_),
    .Y(_22713_));
 sky130_fd_sc_hd__inv_2 _26103_ (.A(_22713_),
    .Y(_22714_));
 sky130_fd_sc_hd__a21o_1 _26104_ (.A1(_22706_),
    .A2(_22707_),
    .B1(_22709_),
    .X(_22715_));
 sky130_fd_sc_hd__nor2_1 _26105_ (.A(_22268_),
    .B(_22269_),
    .Y(_22716_));
 sky130_fd_sc_hd__o211ai_2 _26106_ (.A1(_22271_),
    .A2(_22272_),
    .B1(_22706_),
    .C1(_22707_),
    .Y(_22717_));
 sky130_fd_sc_hd__nand3_1 _26107_ (.A(_22715_),
    .B(_22716_),
    .C(_22717_),
    .Y(_22718_));
 sky130_fd_sc_hd__and3_2 _26108_ (.A(_22712_),
    .B(_22714_),
    .C(_22718_),
    .X(_22719_));
 sky130_fd_sc_hd__clkbuf_2 _26109_ (.A(_22265_),
    .X(_22720_));
 sky130_fd_sc_hd__o21a_1 _26110_ (.A1(_22720_),
    .A2(_22266_),
    .B1(_22222_),
    .X(_22722_));
 sky130_fd_sc_hd__nor2_1 _26111_ (.A(_22222_),
    .B(_22267_),
    .Y(_22723_));
 sky130_fd_sc_hd__o22ai_2 _26112_ (.A1(_22722_),
    .A2(_22723_),
    .B1(_22708_),
    .B2(_22711_),
    .Y(_22724_));
 sky130_fd_sc_hd__o211ai_2 _26113_ (.A1(_22268_),
    .A2(_22269_),
    .B1(_22717_),
    .C1(_22715_),
    .Y(_22725_));
 sky130_fd_sc_hd__a2bb2o_2 _26114_ (.A1_N(_20220_),
    .A2_N(_22065_),
    .B1(_22064_),
    .B2(_20175_),
    .X(_22726_));
 sky130_fd_sc_hd__a31o_1 _26115_ (.A1(_22713_),
    .A2(_22724_),
    .A3(_22725_),
    .B1(_22726_),
    .X(_22727_));
 sky130_fd_sc_hd__nand2_2 _26116_ (.A(_22075_),
    .B(_22087_),
    .Y(_22728_));
 sky130_fd_sc_hd__inv_2 _26117_ (.A(_22728_),
    .Y(_22729_));
 sky130_fd_sc_hd__and2_2 _26118_ (.A(_22064_),
    .B(_20175_),
    .X(_22730_));
 sky130_fd_sc_hd__nand3_1 _26119_ (.A(_22712_),
    .B(_22714_),
    .C(_22718_),
    .Y(_22731_));
 sky130_fd_sc_hd__nand3_1 _26120_ (.A(_22713_),
    .B(_22724_),
    .C(_22725_),
    .Y(_22733_));
 sky130_fd_sc_hd__nand2_1 _26121_ (.A(_22731_),
    .B(_22733_),
    .Y(_22734_));
 sky130_fd_sc_hd__o21ai_1 _26122_ (.A1(_22730_),
    .A2(_22069_),
    .B1(_22734_),
    .Y(_22735_));
 sky130_fd_sc_hd__o211ai_4 _26123_ (.A1(_22719_),
    .A2(_22727_),
    .B1(_22729_),
    .C1(_22735_),
    .Y(_22736_));
 sky130_fd_sc_hd__inv_2 _26124_ (.A(_22726_),
    .Y(_22737_));
 sky130_fd_sc_hd__nand2_1 _26125_ (.A(_22734_),
    .B(_22737_),
    .Y(_22738_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26126_ (.A(_22731_),
    .X(_22739_));
 sky130_fd_sc_hd__o211ai_2 _26127_ (.A1(_22730_),
    .A2(_22069_),
    .B1(_22739_),
    .C1(_22733_),
    .Y(_22740_));
 sky130_fd_sc_hd__nand3_2 _26128_ (.A(_22728_),
    .B(_22738_),
    .C(_22740_),
    .Y(_22741_));
 sky130_fd_sc_hd__nand3_4 _26129_ (.A(_22221_),
    .B(_22736_),
    .C(_22741_),
    .Y(_22742_));
 sky130_fd_sc_hd__nand2_1 _26130_ (.A(_22736_),
    .B(_22741_),
    .Y(_22744_));
 sky130_fd_sc_hd__o22a_1 _26131_ (.A1(_22082_),
    .A2(_22084_),
    .B1(_22089_),
    .B2(_22090_),
    .X(_22745_));
 sky130_fd_sc_hd__nand2_2 _26132_ (.A(_22744_),
    .B(_22745_),
    .Y(_22746_));
 sky130_fd_sc_hd__buf_1 _26133_ (.A(\delay_line[23][8] ),
    .X(_22747_));
 sky130_fd_sc_hd__and2_1 _26134_ (.A(_22747_),
    .B(\delay_line[23][9] ),
    .X(_22748_));
 sky130_fd_sc_hd__clkbuf_2 _26135_ (.A(\delay_line[23][9] ),
    .X(_22749_));
 sky130_fd_sc_hd__nor2_1 _26136_ (.A(_22747_),
    .B(_22749_),
    .Y(_22750_));
 sky130_fd_sc_hd__o2bb2ai_1 _26137_ (.A1_N(_22742_),
    .A2_N(_22746_),
    .B1(_22748_),
    .B2(_22750_),
    .Y(_22751_));
 sky130_fd_sc_hd__and2b_1 _26138_ (.A_N(\delay_line[23][9] ),
    .B(_22747_),
    .X(_22752_));
 sky130_fd_sc_hd__and2b_1 _26139_ (.A_N(_22747_),
    .B(_22749_),
    .X(_22753_));
 sky130_fd_sc_hd__o211ai_2 _26140_ (.A1(_22752_),
    .A2(_22753_),
    .B1(_22742_),
    .C1(_22746_),
    .Y(_22755_));
 sky130_fd_sc_hd__nand3_2 _26141_ (.A(_22220_),
    .B(_22751_),
    .C(_22755_),
    .Y(_22756_));
 sky130_fd_sc_hd__o2bb2ai_1 _26142_ (.A1_N(_22742_),
    .A2_N(_22746_),
    .B1(_22752_),
    .B2(_22753_),
    .Y(_22757_));
 sky130_fd_sc_hd__o211ai_1 _26143_ (.A1(_22748_),
    .A2(_22750_),
    .B1(_22742_),
    .C1(_22746_),
    .Y(_22758_));
 sky130_fd_sc_hd__nand3_2 _26144_ (.A(_22757_),
    .B(_22758_),
    .C(_22219_),
    .Y(_22759_));
 sky130_fd_sc_hd__clkbuf_2 _26145_ (.A(_22111_),
    .X(_22760_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26146_ (.A(\delay_line[23][8] ),
    .X(_22761_));
 sky130_fd_sc_hd__o211a_1 _26147_ (.A1(_22760_),
    .A2(_22747_),
    .B1(_22098_),
    .C1(_22091_),
    .X(_22762_));
 sky130_fd_sc_hd__a21o_1 _26148_ (.A1(_22760_),
    .A2(_22761_),
    .B1(_22762_),
    .X(_22763_));
 sky130_fd_sc_hd__a21oi_2 _26149_ (.A1(_22756_),
    .A2(_22759_),
    .B1(_22763_),
    .Y(_22764_));
 sky130_fd_sc_hd__and3_1 _26150_ (.A(_22763_),
    .B(_22756_),
    .C(_22759_),
    .X(_22766_));
 sky130_fd_sc_hd__nor3_2 _26151_ (.A(_22218_),
    .B(_22764_),
    .C(_22766_),
    .Y(_22767_));
 sky130_fd_sc_hd__a21o_1 _26152_ (.A1(_22756_),
    .A2(_22759_),
    .B1(_22763_),
    .X(_22768_));
 sky130_fd_sc_hd__nand3_2 _26153_ (.A(_22763_),
    .B(_22756_),
    .C(_22759_),
    .Y(_22769_));
 sky130_fd_sc_hd__a21oi_4 _26154_ (.A1(_22768_),
    .A2(_22769_),
    .B1(_22217_),
    .Y(_22770_));
 sky130_fd_sc_hd__o22ai_4 _26155_ (.A1(_22214_),
    .A2(_22216_),
    .B1(_22767_),
    .B2(_22770_),
    .Y(_22771_));
 sky130_fd_sc_hd__o21ai_2 _26156_ (.A1(_22764_),
    .A2(_22766_),
    .B1(_22218_),
    .Y(_22772_));
 sky130_fd_sc_hd__a21oi_4 _26157_ (.A1(_22113_),
    .A2(_22108_),
    .B1(_22214_),
    .Y(_22773_));
 sky130_fd_sc_hd__nand3_2 _26158_ (.A(_22217_),
    .B(_22768_),
    .C(_22769_),
    .Y(_22774_));
 sky130_fd_sc_hd__nand3_2 _26159_ (.A(_22772_),
    .B(_22773_),
    .C(_22774_),
    .Y(_22775_));
 sky130_fd_sc_hd__o2bb2a_2 _26160_ (.A1_N(_22121_),
    .A2_N(_22117_),
    .B1(_22123_),
    .B2(_22114_),
    .X(_22777_));
 sky130_fd_sc_hd__and2_1 _26161_ (.A(_19236_),
    .B(_22760_),
    .X(_22778_));
 sky130_fd_sc_hd__nor2_1 _26162_ (.A(_19236_),
    .B(_22760_),
    .Y(_22779_));
 sky130_fd_sc_hd__or3b_2 _26163_ (.A(_22778_),
    .B(_22779_),
    .C_N(_22128_),
    .X(_22780_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26164_ (.A(_17897_),
    .X(_22781_));
 sky130_fd_sc_hd__clkbuf_2 _26165_ (.A(_22110_),
    .X(_22782_));
 sky130_fd_sc_hd__a2bb2o_1 _26166_ (.A1_N(_22778_),
    .A2_N(_22779_),
    .B1(_22781_),
    .B2(_22782_),
    .X(_22783_));
 sky130_fd_sc_hd__and3b_1 _26167_ (.A_N(_00755_),
    .B(_22780_),
    .C(_22783_),
    .X(_22784_));
 sky130_fd_sc_hd__a21boi_1 _26168_ (.A1(_22780_),
    .A2(_22783_),
    .B1_N(_00755_),
    .Y(_22785_));
 sky130_fd_sc_hd__nor2_1 _26169_ (.A(_22784_),
    .B(_22785_),
    .Y(_22786_));
 sky130_fd_sc_hd__a31o_1 _26170_ (.A1(_22771_),
    .A2(_22775_),
    .A3(_22777_),
    .B1(_22786_),
    .X(_22788_));
 sky130_fd_sc_hd__and3_1 _26171_ (.A(_22116_),
    .B(_22118_),
    .C(_22119_),
    .X(_22789_));
 sky130_fd_sc_hd__o211ai_2 _26172_ (.A1(_22214_),
    .A2(_22216_),
    .B1(_22774_),
    .C1(_22772_),
    .Y(_22790_));
 sky130_fd_sc_hd__o21ai_1 _26173_ (.A1(_22767_),
    .A2(_22770_),
    .B1(_22773_),
    .Y(_22791_));
 sky130_fd_sc_hd__o211ai_4 _26174_ (.A1(_22789_),
    .A2(_22124_),
    .B1(_22790_),
    .C1(_22791_),
    .Y(_22792_));
 sky130_fd_sc_hd__inv_2 _26175_ (.A(_22792_),
    .Y(_22793_));
 sky130_fd_sc_hd__o21a_2 _26176_ (.A1(_21196_),
    .A2(_21197_),
    .B1(_21200_),
    .X(_22794_));
 sky130_fd_sc_hd__inv_2 _26177_ (.A(_22794_),
    .Y(_22795_));
 sky130_fd_sc_hd__nand3_1 _26178_ (.A(_22771_),
    .B(_22775_),
    .C(_22777_),
    .Y(_22796_));
 sky130_fd_sc_hd__nand2_1 _26179_ (.A(_22796_),
    .B(_22792_),
    .Y(_22797_));
 sky130_fd_sc_hd__nand2_1 _26180_ (.A(_22797_),
    .B(_22786_),
    .Y(_22799_));
 sky130_fd_sc_hd__o211ai_2 _26181_ (.A1(_22788_),
    .A2(_22793_),
    .B1(_22795_),
    .C1(_22799_),
    .Y(_22800_));
 sky130_fd_sc_hd__o21ai_1 _26182_ (.A1(_22784_),
    .A2(_22785_),
    .B1(_22797_),
    .Y(_22801_));
 sky130_fd_sc_hd__nand3_1 _26183_ (.A(_22792_),
    .B(_22786_),
    .C(_22796_),
    .Y(_22802_));
 sky130_fd_sc_hd__nand3_2 _26184_ (.A(_22801_),
    .B(_22794_),
    .C(_22802_),
    .Y(_22803_));
 sky130_fd_sc_hd__o32a_1 _26185_ (.A1(_21675_),
    .A2(_22122_),
    .A3(_22124_),
    .B1(_22137_),
    .B2(_22136_),
    .X(_22804_));
 sky130_fd_sc_hd__a21boi_2 _26186_ (.A1(_22800_),
    .A2(_22803_),
    .B1_N(_22804_),
    .Y(_22805_));
 sky130_fd_sc_hd__nor2_1 _26187_ (.A(_22137_),
    .B(_22136_),
    .Y(_22806_));
 sky130_fd_sc_hd__buf_1 _26188_ (.A(_22800_),
    .X(_22807_));
 sky130_fd_sc_hd__o211a_1 _26189_ (.A1(_22126_),
    .A2(_22806_),
    .B1(_22807_),
    .C1(_22803_),
    .X(_22808_));
 sky130_fd_sc_hd__o21ai_1 _26190_ (.A1(_21353_),
    .A2(_21663_),
    .B1(_21661_),
    .Y(_22810_));
 sky130_fd_sc_hd__a21boi_1 _26191_ (.A1(_21576_),
    .A2(_21579_),
    .B1_N(_21573_),
    .Y(_22811_));
 sky130_fd_sc_hd__and2_1 _26192_ (.A(\delay_line[25][7] ),
    .B(\delay_line[25][9] ),
    .X(_22812_));
 sky130_fd_sc_hd__clkbuf_2 _26193_ (.A(_22812_),
    .X(_22813_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26194_ (.A(\delay_line[25][9] ),
    .X(_22814_));
 sky130_fd_sc_hd__o211ai_2 _26195_ (.A1(_20483_),
    .A2(_22814_),
    .B1(_21562_),
    .C1(_19488_),
    .Y(_22815_));
 sky130_fd_sc_hd__nor2_1 _26196_ (.A(\delay_line[25][7] ),
    .B(_22814_),
    .Y(_22816_));
 sky130_fd_sc_hd__o21bai_2 _26197_ (.A1(_22812_),
    .A2(_22816_),
    .B1_N(_21560_),
    .Y(_22817_));
 sky130_fd_sc_hd__o211a_1 _26198_ (.A1(_22813_),
    .A2(_22815_),
    .B1(_17204_),
    .C1(_22817_),
    .X(_22818_));
 sky130_fd_sc_hd__clkbuf_2 _26199_ (.A(_22814_),
    .X(_22819_));
 sky130_fd_sc_hd__a21o_1 _26200_ (.A1(_21565_),
    .A2(_22819_),
    .B1(_22815_),
    .X(_22821_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26201_ (.A(_17204_),
    .X(_22822_));
 sky130_fd_sc_hd__a21o_1 _26202_ (.A1(_22821_),
    .A2(_22817_),
    .B1(_22822_),
    .X(_22823_));
 sky130_fd_sc_hd__o2bb2ai_1 _26203_ (.A1_N(_06766_),
    .A2_N(_21567_),
    .B1(_21564_),
    .B2(_21561_),
    .Y(_22824_));
 sky130_fd_sc_hd__nand3b_2 _26204_ (.A_N(_22818_),
    .B(_22823_),
    .C(_22824_),
    .Y(_22825_));
 sky130_fd_sc_hd__a21oi_1 _26205_ (.A1(_22821_),
    .A2(_22817_),
    .B1(_22822_),
    .Y(_22826_));
 sky130_fd_sc_hd__o21bai_2 _26206_ (.A1(_22818_),
    .A2(_22826_),
    .B1_N(_22824_),
    .Y(_22827_));
 sky130_fd_sc_hd__o21a_1 _26207_ (.A1(_01501_),
    .A2(_01512_),
    .B1(\delay_line[25][1] ),
    .X(_22828_));
 sky130_fd_sc_hd__a21o_1 _26208_ (.A1(_06810_),
    .A2(_17226_),
    .B1(_22828_),
    .X(_22829_));
 sky130_fd_sc_hd__and3_1 _26209_ (.A(_22825_),
    .B(_22827_),
    .C(_22829_),
    .X(_22830_));
 sky130_fd_sc_hd__a21oi_1 _26210_ (.A1(_22825_),
    .A2(_22827_),
    .B1(_22829_),
    .Y(_22832_));
 sky130_fd_sc_hd__nor3_1 _26211_ (.A(_22811_),
    .B(_22830_),
    .C(_22832_),
    .Y(_22833_));
 sky130_fd_sc_hd__o21ai_1 _26212_ (.A1(_22830_),
    .A2(_22832_),
    .B1(_22811_),
    .Y(_22834_));
 sky130_fd_sc_hd__nand3b_2 _26213_ (.A_N(_22833_),
    .B(_22380_),
    .C(_22834_),
    .Y(_22835_));
 sky130_fd_sc_hd__and2_1 _26214_ (.A(_06810_),
    .B(_01490_),
    .X(_22836_));
 sky130_fd_sc_hd__o211ai_1 _26215_ (.A1(_22836_),
    .A2(_22828_),
    .B1(_22825_),
    .C1(_22827_),
    .Y(_22837_));
 sky130_fd_sc_hd__a21o_1 _26216_ (.A1(_22825_),
    .A2(_22827_),
    .B1(_22829_),
    .X(_22838_));
 sky130_fd_sc_hd__a21boi_1 _26217_ (.A1(_22837_),
    .A2(_22838_),
    .B1_N(_22811_),
    .Y(_22839_));
 sky130_fd_sc_hd__o21bai_2 _26218_ (.A1(_22839_),
    .A2(_22833_),
    .B1_N(_22369_),
    .Y(_22840_));
 sky130_fd_sc_hd__o2111ai_2 _26219_ (.A1(_21586_),
    .A2(_21583_),
    .B1(_21591_),
    .C1(_22835_),
    .D1(_22840_),
    .Y(_22841_));
 sky130_fd_sc_hd__o21a_1 _26220_ (.A1(_21586_),
    .A2(_21583_),
    .B1(_21591_),
    .X(_22843_));
 sky130_fd_sc_hd__a21o_1 _26221_ (.A1(_22835_),
    .A2(_22840_),
    .B1(_22843_),
    .X(_22844_));
 sky130_fd_sc_hd__nand4_1 _26222_ (.A(_21585_),
    .B(_20496_),
    .C(_21592_),
    .D(_20482_),
    .Y(_22845_));
 sky130_fd_sc_hd__o2111a_1 _26223_ (.A1(_20502_),
    .A2(_21595_),
    .B1(_22841_),
    .C1(_22844_),
    .D1(_22845_),
    .X(_22846_));
 sky130_fd_sc_hd__nand2_1 _26224_ (.A(_22841_),
    .B(_22844_),
    .Y(_22847_));
 sky130_fd_sc_hd__o21a_1 _26225_ (.A1(_21593_),
    .A2(_21597_),
    .B1(_22847_),
    .X(_22848_));
 sky130_fd_sc_hd__and4_1 _26226_ (.A(_21605_),
    .B(_20451_),
    .C(_19504_),
    .D(_21606_),
    .X(_22849_));
 sky130_fd_sc_hd__or2_1 _26227_ (.A(\delay_line[22][0] ),
    .B(_01402_),
    .X(_22850_));
 sky130_fd_sc_hd__nand2_1 _26228_ (.A(\delay_line[22][0] ),
    .B(\delay_line[22][1] ),
    .Y(_22851_));
 sky130_fd_sc_hd__clkbuf_2 _26229_ (.A(_22851_),
    .X(_22852_));
 sky130_fd_sc_hd__nor2_1 _26230_ (.A(_18316_),
    .B(\delay_line[22][8] ),
    .Y(_22854_));
 sky130_fd_sc_hd__nand2_1 _26231_ (.A(_18316_),
    .B(\delay_line[22][8] ),
    .Y(_22855_));
 sky130_fd_sc_hd__nand3b_2 _26232_ (.A_N(_22854_),
    .B(_22855_),
    .C(_21603_),
    .Y(_22856_));
 sky130_fd_sc_hd__and2_1 _26233_ (.A(\delay_line[22][4] ),
    .B(\delay_line[22][8] ),
    .X(_22857_));
 sky130_fd_sc_hd__o21ai_1 _26234_ (.A1(_22854_),
    .A2(_22857_),
    .B1(_21601_),
    .Y(_22858_));
 sky130_fd_sc_hd__a22o_1 _26235_ (.A1(_22850_),
    .A2(_22852_),
    .B1(_22856_),
    .B2(_22858_),
    .X(_22859_));
 sky130_fd_sc_hd__nor2_1 _26236_ (.A(\delay_line[22][0] ),
    .B(_01402_),
    .Y(_22860_));
 sky130_fd_sc_hd__nand4b_2 _26237_ (.A_N(_22860_),
    .B(_22852_),
    .C(_22856_),
    .D(_22858_),
    .Y(_22861_));
 sky130_fd_sc_hd__nand2_1 _26238_ (.A(_21602_),
    .B(_21606_),
    .Y(_22862_));
 sky130_fd_sc_hd__nand3_1 _26239_ (.A(_22859_),
    .B(_22861_),
    .C(_22862_),
    .Y(_22863_));
 sky130_fd_sc_hd__a21o_1 _26240_ (.A1(_22859_),
    .A2(_22861_),
    .B1(_22862_),
    .X(_22865_));
 sky130_fd_sc_hd__nand2_1 _26241_ (.A(_22863_),
    .B(_22865_),
    .Y(_22866_));
 sky130_fd_sc_hd__a311oi_2 _26242_ (.A1(_19507_),
    .A2(_21608_),
    .A3(_20452_),
    .B1(_22849_),
    .C1(_22866_),
    .Y(_22867_));
 sky130_fd_sc_hd__o21a_1 _26243_ (.A1(_22849_),
    .A2(_21610_),
    .B1(_22866_),
    .X(_22868_));
 sky130_fd_sc_hd__nand4_2 _26244_ (.A(_21643_),
    .B(_20456_),
    .C(_21640_),
    .D(_20474_),
    .Y(_22869_));
 sky130_fd_sc_hd__o21a_1 _26245_ (.A1(_01446_),
    .A2(_06920_),
    .B1(_23687_),
    .X(_22870_));
 sky130_fd_sc_hd__clkbuf_2 _26246_ (.A(_20467_),
    .X(_22871_));
 sky130_fd_sc_hd__o22a_1 _26247_ (.A1(_22871_),
    .A2(_21614_),
    .B1(_21627_),
    .B2(_21629_),
    .X(_22872_));
 sky130_fd_sc_hd__o21ai_1 _26248_ (.A1(_21613_),
    .A2(_22872_),
    .B1(_21634_),
    .Y(_22873_));
 sky130_fd_sc_hd__inv_2 _26249_ (.A(net343),
    .Y(_22874_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26250_ (.A(_22874_),
    .X(_22876_));
 sky130_fd_sc_hd__inv_2 _26251_ (.A(_19512_),
    .Y(_22877_));
 sky130_fd_sc_hd__o21a_1 _26252_ (.A1(_21616_),
    .A2(_19513_),
    .B1(_20458_),
    .X(_22878_));
 sky130_fd_sc_hd__o21ai_1 _26253_ (.A1(_22876_),
    .A2(_22877_),
    .B1(_22878_),
    .Y(_22879_));
 sky130_fd_sc_hd__and2_2 _26254_ (.A(\delay_line[24][4] ),
    .B(_19512_),
    .X(_22880_));
 sky130_fd_sc_hd__nor2_1 _26255_ (.A(_21616_),
    .B(_19513_),
    .Y(_22881_));
 sky130_fd_sc_hd__o21bai_2 _26256_ (.A1(_22880_),
    .A2(_22881_),
    .B1_N(_20458_),
    .Y(_22882_));
 sky130_fd_sc_hd__clkbuf_2 _26257_ (.A(net342),
    .X(_22883_));
 sky130_fd_sc_hd__clkbuf_2 _26258_ (.A(_22883_),
    .X(_22884_));
 sky130_fd_sc_hd__a21o_1 _26259_ (.A1(_22879_),
    .A2(_22882_),
    .B1(_22884_),
    .X(_22885_));
 sky130_fd_sc_hd__o21ai_2 _26260_ (.A1(_21616_),
    .A2(_19513_),
    .B1(_17007_),
    .Y(_22887_));
 sky130_fd_sc_hd__o211ai_2 _26261_ (.A1(_22880_),
    .A2(_22887_),
    .B1(_22884_),
    .C1(_22882_),
    .Y(_22888_));
 sky130_fd_sc_hd__nand3_2 _26262_ (.A(_22885_),
    .B(_21627_),
    .C(_22888_),
    .Y(_22889_));
 sky130_fd_sc_hd__o211a_1 _26263_ (.A1(_22880_),
    .A2(_22887_),
    .B1(_22884_),
    .C1(_22882_),
    .X(_22890_));
 sky130_fd_sc_hd__clkbuf_2 _26264_ (.A(_22884_),
    .X(_22891_));
 sky130_fd_sc_hd__a21oi_1 _26265_ (.A1(_22879_),
    .A2(_22882_),
    .B1(_22891_),
    .Y(_22892_));
 sky130_fd_sc_hd__o21ai_2 _26266_ (.A1(_22890_),
    .A2(_22892_),
    .B1(_21623_),
    .Y(_22893_));
 sky130_fd_sc_hd__o21a_1 _26267_ (.A1(_06909_),
    .A2(_21615_),
    .B1(_21618_),
    .X(_22894_));
 sky130_fd_sc_hd__a21o_1 _26268_ (.A1(_22889_),
    .A2(_22893_),
    .B1(_22894_),
    .X(_22895_));
 sky130_fd_sc_hd__o2111ai_1 _26269_ (.A1(_06920_),
    .A2(_21615_),
    .B1(_21618_),
    .C1(_22889_),
    .D1(_22893_),
    .Y(_22896_));
 sky130_fd_sc_hd__nand3_2 _26270_ (.A(_22873_),
    .B(_22895_),
    .C(_22896_),
    .Y(_22898_));
 sky130_fd_sc_hd__a21oi_1 _26271_ (.A1(_22889_),
    .A2(_22893_),
    .B1(_22894_),
    .Y(_22899_));
 sky130_fd_sc_hd__and3_1 _26272_ (.A(_22893_),
    .B(_22894_),
    .C(_22889_),
    .X(_22900_));
 sky130_fd_sc_hd__o21bai_2 _26273_ (.A1(_22899_),
    .A2(_22900_),
    .B1_N(_22873_),
    .Y(_22901_));
 sky130_fd_sc_hd__nor2_1 _26274_ (.A(_17040_),
    .B(_06920_),
    .Y(_22902_));
 sky130_fd_sc_hd__o2bb2ai_1 _26275_ (.A1_N(_22898_),
    .A2_N(_22901_),
    .B1(_19508_),
    .B2(_22902_),
    .Y(_22903_));
 sky130_fd_sc_hd__o2111ai_4 _26276_ (.A1(_17040_),
    .A2(_06931_),
    .B1(_01457_),
    .C1(_22898_),
    .D1(_22901_),
    .Y(_22904_));
 sky130_fd_sc_hd__a221o_1 _26277_ (.A1(_21639_),
    .A2(_22870_),
    .B1(_22903_),
    .B2(_22904_),
    .C1(_21642_),
    .X(_22905_));
 sky130_fd_sc_hd__and3_1 _26278_ (.A(_21639_),
    .B(_22870_),
    .C(_21638_),
    .X(_22906_));
 sky130_fd_sc_hd__o211ai_2 _26279_ (.A1(_21642_),
    .A2(_22906_),
    .B1(_22904_),
    .C1(_22903_),
    .Y(_22907_));
 sky130_fd_sc_hd__and4_1 _26280_ (.A(_22869_),
    .B(_21647_),
    .C(_22905_),
    .D(_22907_),
    .X(_22909_));
 sky130_fd_sc_hd__a22oi_2 _26281_ (.A1(_22869_),
    .A2(_21647_),
    .B1(_22905_),
    .B2(_22907_),
    .Y(_22910_));
 sky130_fd_sc_hd__nor4_1 _26282_ (.A(_22867_),
    .B(_22868_),
    .C(_22909_),
    .D(_22910_),
    .Y(_22911_));
 sky130_fd_sc_hd__o22a_1 _26283_ (.A1(_22867_),
    .A2(_22868_),
    .B1(_22909_),
    .B2(_22910_),
    .X(_22912_));
 sky130_fd_sc_hd__nor4_1 _26284_ (.A(_22846_),
    .B(_22848_),
    .C(net137),
    .D(_22912_),
    .Y(_22913_));
 sky130_fd_sc_hd__o22a_1 _26285_ (.A1(_22846_),
    .A2(_22848_),
    .B1(net137),
    .B2(_22912_),
    .X(_22914_));
 sky130_fd_sc_hd__or2_1 _26286_ (.A(net112),
    .B(_22914_),
    .X(_22915_));
 sky130_fd_sc_hd__and3_1 _26287_ (.A(_21406_),
    .B(_21443_),
    .C(_22915_),
    .X(_22916_));
 sky130_fd_sc_hd__a21oi_1 _26288_ (.A1(_21406_),
    .A2(_21443_),
    .B1(_22915_),
    .Y(_22917_));
 sky130_fd_sc_hd__nor2_1 _26289_ (.A(_22916_),
    .B(_22917_),
    .Y(_22918_));
 sky130_fd_sc_hd__o21a_1 _26290_ (.A1(_21649_),
    .A2(net113),
    .B1(_22918_),
    .X(_22920_));
 sky130_fd_sc_hd__nor3_1 _26291_ (.A(_21649_),
    .B(net113),
    .C(_22918_),
    .Y(_22921_));
 sky130_fd_sc_hd__nor2_1 _26292_ (.A(_22920_),
    .B(_22921_),
    .Y(_22922_));
 sky130_fd_sc_hd__nand2_1 _26293_ (.A(_21445_),
    .B(_21551_),
    .Y(_22923_));
 sky130_fd_sc_hd__nand2_2 _26294_ (.A(_21550_),
    .B(_22923_),
    .Y(_22924_));
 sky130_fd_sc_hd__clkbuf_2 _26295_ (.A(\delay_line[18][8] ),
    .X(_22925_));
 sky130_fd_sc_hd__nor2_1 _26296_ (.A(\delay_line[18][4] ),
    .B(_22925_),
    .Y(_22926_));
 sky130_fd_sc_hd__and2_1 _26297_ (.A(\delay_line[18][4] ),
    .B(_22925_),
    .X(_22927_));
 sky130_fd_sc_hd__o21ai_2 _26298_ (.A1(_22926_),
    .A2(_22927_),
    .B1(_21364_),
    .Y(_22928_));
 sky130_fd_sc_hd__xnor2_1 _26299_ (.A(_23852_),
    .B(_01666_),
    .Y(_22929_));
 sky130_fd_sc_hd__clkbuf_2 _26300_ (.A(\delay_line[18][8] ),
    .X(_22931_));
 sky130_fd_sc_hd__nand2_1 _26301_ (.A(_18384_),
    .B(_22931_),
    .Y(_22932_));
 sky130_fd_sc_hd__nand3b_2 _26302_ (.A_N(_22926_),
    .B(_22932_),
    .C(_21359_),
    .Y(_22933_));
 sky130_fd_sc_hd__nand3_2 _26303_ (.A(_22928_),
    .B(_22929_),
    .C(_22933_),
    .Y(_22934_));
 sky130_fd_sc_hd__a21o_1 _26304_ (.A1(_22933_),
    .A2(_22928_),
    .B1(_22929_),
    .X(_22935_));
 sky130_fd_sc_hd__and4_1 _26305_ (.A(_21365_),
    .B(_21366_),
    .C(_22934_),
    .D(_22935_),
    .X(_22936_));
 sky130_fd_sc_hd__a22oi_4 _26306_ (.A1(_21365_),
    .A2(_21367_),
    .B1(_22934_),
    .B2(_22935_),
    .Y(_22937_));
 sky130_fd_sc_hd__nor2_1 _26307_ (.A(_22936_),
    .B(_22937_),
    .Y(_22938_));
 sky130_fd_sc_hd__a41o_1 _26308_ (.A1(_19397_),
    .A2(_20544_),
    .A3(_21367_),
    .A4(_21368_),
    .B1(_21371_),
    .X(_22939_));
 sky130_fd_sc_hd__xnor2_1 _26309_ (.A(_22938_),
    .B(_22939_),
    .Y(_22940_));
 sky130_fd_sc_hd__buf_1 _26310_ (.A(_21384_),
    .X(_22942_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26311_ (.A(_21394_),
    .X(_22943_));
 sky130_fd_sc_hd__clkbuf_2 _26312_ (.A(_21378_),
    .X(_22944_));
 sky130_fd_sc_hd__a22oi_2 _26313_ (.A1(_22944_),
    .A2(_20548_),
    .B1(_21377_),
    .B2(_07393_),
    .Y(_22945_));
 sky130_fd_sc_hd__clkbuf_2 _26314_ (.A(\delay_line[19][8] ),
    .X(_22946_));
 sky130_fd_sc_hd__nor2_1 _26315_ (.A(_21381_),
    .B(_22946_),
    .Y(_22947_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26316_ (.A(\delay_line[19][8] ),
    .X(_22948_));
 sky130_fd_sc_hd__and2_1 _26317_ (.A(_21381_),
    .B(_22948_),
    .X(_22949_));
 sky130_fd_sc_hd__nand2_1 _26318_ (.A(_20560_),
    .B(_21381_),
    .Y(_22950_));
 sky130_fd_sc_hd__o21ai_2 _26319_ (.A1(_22947_),
    .A2(_22949_),
    .B1(_22950_),
    .Y(_22951_));
 sky130_fd_sc_hd__buf_1 _26320_ (.A(_21375_),
    .X(_22953_));
 sky130_fd_sc_hd__inv_2 _26321_ (.A(_22948_),
    .Y(_22954_));
 sky130_fd_sc_hd__nand2_1 _26322_ (.A(_22953_),
    .B(_22954_),
    .Y(_22955_));
 sky130_fd_sc_hd__buf_1 _26323_ (.A(_18367_),
    .X(_22956_));
 sky130_fd_sc_hd__a21o_1 _26324_ (.A1(_22951_),
    .A2(_22955_),
    .B1(_22956_),
    .X(_22957_));
 sky130_fd_sc_hd__o211ai_1 _26325_ (.A1(_22946_),
    .A2(_22950_),
    .B1(_22956_),
    .C1(_22951_),
    .Y(_22958_));
 sky130_fd_sc_hd__nand3b_2 _26326_ (.A_N(_22945_),
    .B(_22957_),
    .C(_22958_),
    .Y(_22959_));
 sky130_fd_sc_hd__a21oi_1 _26327_ (.A1(_22951_),
    .A2(_22955_),
    .B1(_18368_),
    .Y(_22960_));
 sky130_fd_sc_hd__and3_1 _26328_ (.A(_22951_),
    .B(_22955_),
    .C(_22956_),
    .X(_22961_));
 sky130_fd_sc_hd__o21ai_2 _26329_ (.A1(_22960_),
    .A2(_22961_),
    .B1(_22945_),
    .Y(_22962_));
 sky130_fd_sc_hd__nand2_1 _26330_ (.A(_23874_),
    .B(_07448_),
    .Y(_22964_));
 sky130_fd_sc_hd__o21ai_1 _26331_ (.A1(_23885_),
    .A2(_07404_),
    .B1(_22964_),
    .Y(_22965_));
 sky130_fd_sc_hd__nand3_2 _26332_ (.A(_22959_),
    .B(_22962_),
    .C(_22965_),
    .Y(_22966_));
 sky130_fd_sc_hd__a21o_1 _26333_ (.A1(_22959_),
    .A2(_22962_),
    .B1(_22965_),
    .X(_22967_));
 sky130_fd_sc_hd__nand4_1 _26334_ (.A(_22942_),
    .B(_22943_),
    .C(_22966_),
    .D(_22967_),
    .Y(_22968_));
 sky130_fd_sc_hd__a22o_1 _26335_ (.A1(_22942_),
    .A2(_22943_),
    .B1(_22966_),
    .B2(_22967_),
    .X(_22969_));
 sky130_fd_sc_hd__nand3_1 _26336_ (.A(_20566_),
    .B(_20567_),
    .C(_20565_),
    .Y(_22970_));
 sky130_fd_sc_hd__a21oi_1 _26337_ (.A1(_22943_),
    .A2(_21395_),
    .B1(_21393_),
    .Y(_22971_));
 sky130_fd_sc_hd__o21ai_1 _26338_ (.A1(_22970_),
    .A2(_22971_),
    .B1(_21396_),
    .Y(_22972_));
 sky130_fd_sc_hd__nand3_1 _26339_ (.A(_22968_),
    .B(_22969_),
    .C(_22972_),
    .Y(_22973_));
 sky130_fd_sc_hd__a22oi_2 _26340_ (.A1(_22942_),
    .A2(_22943_),
    .B1(_22966_),
    .B2(_22967_),
    .Y(_22975_));
 sky130_fd_sc_hd__and4_1 _26341_ (.A(_22942_),
    .B(_21394_),
    .C(_22966_),
    .D(_22967_),
    .X(_22976_));
 sky130_fd_sc_hd__o221ai_2 _26342_ (.A1(_22971_),
    .A2(_22970_),
    .B1(_22975_),
    .B2(_22976_),
    .C1(_21396_),
    .Y(_22977_));
 sky130_fd_sc_hd__o21ai_1 _26343_ (.A1(_20573_),
    .A2(_21403_),
    .B1(_21401_),
    .Y(_22978_));
 sky130_fd_sc_hd__and3_1 _26344_ (.A(_22973_),
    .B(_22977_),
    .C(_22978_),
    .X(_22979_));
 sky130_fd_sc_hd__a21oi_1 _26345_ (.A1(_22973_),
    .A2(_22977_),
    .B1(_22978_),
    .Y(_22980_));
 sky130_fd_sc_hd__nor3_1 _26346_ (.A(_22940_),
    .B(_22979_),
    .C(_22980_),
    .Y(_22981_));
 sky130_fd_sc_hd__o21ai_4 _26347_ (.A1(_01622_),
    .A2(_21433_),
    .B1(_21422_),
    .Y(_22982_));
 sky130_fd_sc_hd__a2bb2o_1 _26348_ (.A1_N(_21418_),
    .A2_N(_21413_),
    .B1(_21419_),
    .B2(_21414_),
    .X(_22983_));
 sky130_fd_sc_hd__buf_1 _26349_ (.A(net359),
    .X(_22984_));
 sky130_fd_sc_hd__nor2_1 _26350_ (.A(_21415_),
    .B(_22984_),
    .Y(_22986_));
 sky130_fd_sc_hd__and2_1 _26351_ (.A(\delay_line[21][7] ),
    .B(net359),
    .X(_22987_));
 sky130_fd_sc_hd__nand2_1 _26352_ (.A(_20521_),
    .B(_21415_),
    .Y(_22988_));
 sky130_fd_sc_hd__o21ai_1 _26353_ (.A1(_22986_),
    .A2(_22987_),
    .B1(_22988_),
    .Y(_22989_));
 sky130_fd_sc_hd__or2_1 _26354_ (.A(_22984_),
    .B(_22988_),
    .X(_22990_));
 sky130_fd_sc_hd__a21o_1 _26355_ (.A1(_22989_),
    .A2(_22990_),
    .B1(_18352_),
    .X(_22991_));
 sky130_fd_sc_hd__clkbuf_2 _26356_ (.A(_22984_),
    .X(_22992_));
 sky130_fd_sc_hd__o211ai_2 _26357_ (.A1(_22992_),
    .A2(_22988_),
    .B1(_18352_),
    .C1(_22989_),
    .Y(_22993_));
 sky130_fd_sc_hd__and3_1 _26358_ (.A(_22983_),
    .B(_22991_),
    .C(_22993_),
    .X(_22994_));
 sky130_fd_sc_hd__a21o_1 _26359_ (.A1(_22991_),
    .A2(_22993_),
    .B1(_22983_),
    .X(_22995_));
 sky130_fd_sc_hd__nand2_1 _26360_ (.A(_23984_),
    .B(_07316_),
    .Y(_22997_));
 sky130_fd_sc_hd__o211ai_4 _26361_ (.A1(_07338_),
    .A2(_07327_),
    .B1(_22995_),
    .C1(_22997_),
    .Y(_22998_));
 sky130_fd_sc_hd__nand3_2 _26362_ (.A(_22983_),
    .B(_22991_),
    .C(_22993_),
    .Y(_22999_));
 sky130_fd_sc_hd__o21a_1 _26363_ (.A1(_23995_),
    .A2(_07327_),
    .B1(_22997_),
    .X(_23000_));
 sky130_fd_sc_hd__a21o_1 _26364_ (.A1(_22999_),
    .A2(_22995_),
    .B1(_23000_),
    .X(_23001_));
 sky130_fd_sc_hd__o21ai_4 _26365_ (.A1(_22994_),
    .A2(_22998_),
    .B1(_23001_),
    .Y(_23002_));
 sky130_fd_sc_hd__xor2_4 _26366_ (.A(_22982_),
    .B(_23002_),
    .X(_23003_));
 sky130_fd_sc_hd__a21o_1 _26367_ (.A1(_21435_),
    .A2(_21436_),
    .B1(_23003_),
    .X(_23004_));
 sky130_fd_sc_hd__nand3_1 _26368_ (.A(_21435_),
    .B(_21436_),
    .C(_23003_),
    .Y(_23005_));
 sky130_fd_sc_hd__nand2_2 _26369_ (.A(_23004_),
    .B(_23005_),
    .Y(_23006_));
 sky130_fd_sc_hd__a21boi_4 _26370_ (.A1(_21440_),
    .A2(_20538_),
    .B1_N(_21439_),
    .Y(_23008_));
 sky130_fd_sc_hd__xnor2_2 _26371_ (.A(_23006_),
    .B(_23008_),
    .Y(_23009_));
 sky130_fd_sc_hd__o21ai_1 _26372_ (.A1(_22979_),
    .A2(_22980_),
    .B1(_22940_),
    .Y(_23010_));
 sky130_fd_sc_hd__inv_2 _26373_ (.A(_23010_),
    .Y(_23011_));
 sky130_fd_sc_hd__nor3_4 _26374_ (.A(_22981_),
    .B(_23009_),
    .C(_23011_),
    .Y(_23012_));
 sky130_fd_sc_hd__o21a_1 _26375_ (.A1(_23011_),
    .A2(net117),
    .B1(_23009_),
    .X(_23013_));
 sky130_fd_sc_hd__nor2_2 _26376_ (.A(_23012_),
    .B(_23013_),
    .Y(_23014_));
 sky130_fd_sc_hd__nand2_1 _26377_ (.A(_21531_),
    .B(_21532_),
    .Y(_23015_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26378_ (.A(\delay_line[16][5] ),
    .X(_23016_));
 sky130_fd_sc_hd__o21ai_2 _26379_ (.A1(_21514_),
    .A2(_23016_),
    .B1(_16656_),
    .Y(_23017_));
 sky130_fd_sc_hd__a21o_1 _26380_ (.A1(_18399_),
    .A2(_19435_),
    .B1(_23017_),
    .X(_23019_));
 sky130_fd_sc_hd__and2_1 _26381_ (.A(_21514_),
    .B(_23016_),
    .X(_23020_));
 sky130_fd_sc_hd__nor2_1 _26382_ (.A(_18399_),
    .B(_19435_),
    .Y(_23021_));
 sky130_fd_sc_hd__o21ai_2 _26383_ (.A1(_23020_),
    .A2(_23021_),
    .B1(_16667_),
    .Y(_23022_));
 sky130_fd_sc_hd__clkbuf_2 _26384_ (.A(net383),
    .X(_23023_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26385_ (.A(_23023_),
    .X(_23024_));
 sky130_fd_sc_hd__a21oi_1 _26386_ (.A1(_23019_),
    .A2(_23022_),
    .B1(_23024_),
    .Y(_23025_));
 sky130_fd_sc_hd__clkbuf_2 _26387_ (.A(_23024_),
    .X(_23026_));
 sky130_fd_sc_hd__o211ai_2 _26388_ (.A1(_23020_),
    .A2(_23017_),
    .B1(_23026_),
    .C1(_23022_),
    .Y(_23027_));
 sky130_fd_sc_hd__nand3b_1 _26389_ (.A_N(_23025_),
    .B(_21525_),
    .C(_23027_),
    .Y(_23028_));
 sky130_fd_sc_hd__and3_1 _26390_ (.A(_23022_),
    .B(_23024_),
    .C(_23019_),
    .X(_23030_));
 sky130_fd_sc_hd__o21ai_2 _26391_ (.A1(_23030_),
    .A2(_23025_),
    .B1(_21521_),
    .Y(_23031_));
 sky130_fd_sc_hd__o21a_1 _26392_ (.A1(_21509_),
    .A2(_21513_),
    .B1(_21515_),
    .X(_23032_));
 sky130_fd_sc_hd__a21o_1 _26393_ (.A1(_23028_),
    .A2(_23031_),
    .B1(_23032_),
    .X(_23033_));
 sky130_fd_sc_hd__o2111ai_2 _26394_ (.A1(_21536_),
    .A2(_21513_),
    .B1(_21515_),
    .C1(_23028_),
    .D1(_23031_),
    .Y(_23034_));
 sky130_fd_sc_hd__nand3_1 _26395_ (.A(_23015_),
    .B(_23033_),
    .C(_23034_),
    .Y(_23035_));
 sky130_fd_sc_hd__a21o_1 _26396_ (.A1(_23033_),
    .A2(_23034_),
    .B1(_23015_),
    .X(_23036_));
 sky130_fd_sc_hd__a21oi_1 _26397_ (.A1(_23035_),
    .A2(_23036_),
    .B1(_21511_),
    .Y(_23037_));
 sky130_fd_sc_hd__and3_1 _26398_ (.A(_23036_),
    .B(_21511_),
    .C(_23035_),
    .X(_23038_));
 sky130_fd_sc_hd__o31a_1 _26399_ (.A1(_16645_),
    .A2(_19437_),
    .A3(_21535_),
    .B1(_21538_),
    .X(_23039_));
 sky130_fd_sc_hd__o21ai_2 _26400_ (.A1(_23037_),
    .A2(_23038_),
    .B1(_23039_),
    .Y(_23041_));
 sky130_fd_sc_hd__o21ai_2 _26401_ (.A1(_21508_),
    .A2(_21544_),
    .B1(_21542_),
    .Y(_23042_));
 sky130_fd_sc_hd__a21o_1 _26402_ (.A1(_23035_),
    .A2(_23036_),
    .B1(_21511_),
    .X(_23043_));
 sky130_fd_sc_hd__a21oi_2 _26403_ (.A1(_21538_),
    .A2(_21539_),
    .B1(_23038_),
    .Y(_23044_));
 sky130_fd_sc_hd__a21boi_1 _26404_ (.A1(_23043_),
    .A2(_23044_),
    .B1_N(_23041_),
    .Y(_23045_));
 sky130_fd_sc_hd__nor2_1 _26405_ (.A(_23042_),
    .B(_23045_),
    .Y(_23046_));
 sky130_fd_sc_hd__a21oi_1 _26406_ (.A1(_23041_),
    .A2(_23042_),
    .B1(_23046_),
    .Y(_23047_));
 sky130_fd_sc_hd__a21oi_1 _26407_ (.A1(_21491_),
    .A2(_07173_),
    .B1(net394),
    .Y(_23048_));
 sky130_fd_sc_hd__and3_1 _26408_ (.A(net394),
    .B(_16821_),
    .C(_20584_),
    .X(_23049_));
 sky130_fd_sc_hd__and2_1 _26409_ (.A(net392),
    .B(_18405_),
    .X(_23050_));
 sky130_fd_sc_hd__buf_1 _26410_ (.A(\delay_line[14][4] ),
    .X(_23052_));
 sky130_fd_sc_hd__nor2_1 _26411_ (.A(_16821_),
    .B(_23052_),
    .Y(_23053_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26412_ (.A(net390),
    .X(_23054_));
 sky130_fd_sc_hd__o21bai_1 _26413_ (.A1(_23050_),
    .A2(_23053_),
    .B1_N(_23054_),
    .Y(_23055_));
 sky130_fd_sc_hd__o21ai_1 _26414_ (.A1(net392),
    .A2(_18405_),
    .B1(_23054_),
    .Y(_23056_));
 sky130_fd_sc_hd__a21o_1 _26415_ (.A1(_16821_),
    .A2(_23052_),
    .B1(_23056_),
    .X(_23057_));
 sky130_fd_sc_hd__and3_1 _26416_ (.A(_23055_),
    .B(_21494_),
    .C(_23057_),
    .X(_23058_));
 sky130_fd_sc_hd__a21oi_1 _26417_ (.A1(_23057_),
    .A2(_23055_),
    .B1(_21494_),
    .Y(_23059_));
 sky130_fd_sc_hd__nor4_1 _26418_ (.A(_23048_),
    .B(_23049_),
    .C(_23058_),
    .D(_23059_),
    .Y(_23060_));
 sky130_fd_sc_hd__or2_1 _26419_ (.A(_23048_),
    .B(_23049_),
    .X(_23061_));
 sky130_fd_sc_hd__o21ai_1 _26420_ (.A1(_23058_),
    .A2(_23059_),
    .B1(_23061_),
    .Y(_23063_));
 sky130_fd_sc_hd__or2b_2 _26421_ (.A(_23060_),
    .B_N(_23063_),
    .X(_23064_));
 sky130_fd_sc_hd__o211ai_2 _26422_ (.A1(_21501_),
    .A2(_21489_),
    .B1(_21499_),
    .C1(_23064_),
    .Y(_23065_));
 sky130_fd_sc_hd__o21ai_1 _26423_ (.A1(_21501_),
    .A2(_21489_),
    .B1(_21499_),
    .Y(_23066_));
 sky130_fd_sc_hd__nand3b_1 _26424_ (.A_N(_23060_),
    .B(_23063_),
    .C(_23066_),
    .Y(_23067_));
 sky130_fd_sc_hd__nand4_2 _26425_ (.A(_23065_),
    .B(_21502_),
    .C(_20593_),
    .D(_23067_),
    .Y(_23068_));
 sky130_fd_sc_hd__a22o_1 _26426_ (.A1(_20593_),
    .A2(_21502_),
    .B1(_23067_),
    .B2(_23065_),
    .X(_23069_));
 sky130_fd_sc_hd__nand2_2 _26427_ (.A(_23068_),
    .B(_23069_),
    .Y(_23070_));
 sky130_fd_sc_hd__nor2_1 _26428_ (.A(_21467_),
    .B(_21468_),
    .Y(_23071_));
 sky130_fd_sc_hd__o21a_1 _26429_ (.A1(_21463_),
    .A2(_21464_),
    .B1(_21465_),
    .X(_23072_));
 sky130_fd_sc_hd__o21ai_1 _26430_ (.A1(_23071_),
    .A2(_23072_),
    .B1(_21462_),
    .Y(_23074_));
 sky130_fd_sc_hd__and2_2 _26431_ (.A(_20599_),
    .B(net386),
    .X(_23075_));
 sky130_fd_sc_hd__clkbuf_2 _26432_ (.A(net386),
    .X(_23076_));
 sky130_fd_sc_hd__o21ai_2 _26433_ (.A1(_20600_),
    .A2(_23076_),
    .B1(_21450_),
    .Y(_23077_));
 sky130_fd_sc_hd__buf_2 _26434_ (.A(net386),
    .X(_23078_));
 sky130_fd_sc_hd__nor2_1 _26435_ (.A(_20599_),
    .B(_23078_),
    .Y(_23079_));
 sky130_fd_sc_hd__o21bai_2 _26436_ (.A1(_23075_),
    .A2(_23079_),
    .B1_N(_21450_),
    .Y(_23080_));
 sky130_fd_sc_hd__o211ai_1 _26437_ (.A1(_23075_),
    .A2(_23077_),
    .B1(_18411_),
    .C1(_23080_),
    .Y(_23081_));
 sky130_fd_sc_hd__nand2_1 _26438_ (.A(_20600_),
    .B(_23076_),
    .Y(_23082_));
 sky130_fd_sc_hd__nand3b_1 _26439_ (.A_N(_23079_),
    .B(_21451_),
    .C(_23082_),
    .Y(_23083_));
 sky130_fd_sc_hd__a21o_1 _26440_ (.A1(_23083_),
    .A2(_23080_),
    .B1(_18411_),
    .X(_23085_));
 sky130_fd_sc_hd__o2bb2ai_1 _26441_ (.A1_N(_07074_),
    .A2_N(_21456_),
    .B1(_21453_),
    .B2(_21451_),
    .Y(_23086_));
 sky130_fd_sc_hd__nand3_2 _26442_ (.A(_23081_),
    .B(_23085_),
    .C(_23086_),
    .Y(_23087_));
 sky130_fd_sc_hd__o211a_1 _26443_ (.A1(_23075_),
    .A2(_23077_),
    .B1(_16733_),
    .C1(_23080_),
    .X(_23088_));
 sky130_fd_sc_hd__a21oi_1 _26444_ (.A1(_23083_),
    .A2(_23080_),
    .B1(_18411_),
    .Y(_23089_));
 sky130_fd_sc_hd__o21bai_2 _26445_ (.A1(_23088_),
    .A2(_23089_),
    .B1_N(_23086_),
    .Y(_23090_));
 sky130_fd_sc_hd__o21a_1 _26446_ (.A1(\delay_line[15][0] ),
    .A2(_07063_),
    .B1(_16722_),
    .X(_23091_));
 sky130_fd_sc_hd__and3b_1 _26447_ (.A_N(_22391_),
    .B(\delay_line[15][1] ),
    .C(_20606_),
    .X(_23092_));
 sky130_fd_sc_hd__nor2_1 _26448_ (.A(_23091_),
    .B(_23092_),
    .Y(_23093_));
 sky130_fd_sc_hd__a21bo_1 _26449_ (.A1(_23087_),
    .A2(_23090_),
    .B1_N(_23093_),
    .X(_23094_));
 sky130_fd_sc_hd__o211ai_1 _26450_ (.A1(_23091_),
    .A2(_23092_),
    .B1(_23087_),
    .C1(_23090_),
    .Y(_23096_));
 sky130_fd_sc_hd__nand3b_2 _26451_ (.A_N(_23074_),
    .B(_23094_),
    .C(_23096_),
    .Y(_23097_));
 sky130_fd_sc_hd__nand3_1 _26452_ (.A(_23087_),
    .B(_23090_),
    .C(_23093_),
    .Y(_23098_));
 sky130_fd_sc_hd__a21o_1 _26453_ (.A1(_23087_),
    .A2(_23090_),
    .B1(_23093_),
    .X(_23099_));
 sky130_fd_sc_hd__nand3_2 _26454_ (.A(_23074_),
    .B(_23098_),
    .C(_23099_),
    .Y(_23100_));
 sky130_fd_sc_hd__nand3_2 _26455_ (.A(_23097_),
    .B(_23100_),
    .C(_22413_),
    .Y(_23101_));
 sky130_fd_sc_hd__a21o_1 _26456_ (.A1(_23097_),
    .A2(_23100_),
    .B1(_22413_),
    .X(_23102_));
 sky130_fd_sc_hd__o2111ai_4 _26457_ (.A1(_21448_),
    .A2(_21478_),
    .B1(_21476_),
    .C1(_23101_),
    .D1(_23102_),
    .Y(_23103_));
 sky130_fd_sc_hd__a22o_1 _26458_ (.A1(_21476_),
    .A2(_21477_),
    .B1(_23101_),
    .B2(_23102_),
    .X(_23104_));
 sky130_fd_sc_hd__a22oi_2 _26459_ (.A1(_21483_),
    .A2(_21487_),
    .B1(_23103_),
    .B2(_23104_),
    .Y(_23105_));
 sky130_fd_sc_hd__and4_1 _26460_ (.A(_21483_),
    .B(_21487_),
    .C(_23103_),
    .D(_23104_),
    .X(_23107_));
 sky130_fd_sc_hd__or3_1 _26461_ (.A(_23070_),
    .B(_23105_),
    .C(_23107_),
    .X(_23108_));
 sky130_fd_sc_hd__o21ai_1 _26462_ (.A1(_23105_),
    .A2(_23107_),
    .B1(_23070_),
    .Y(_23109_));
 sky130_fd_sc_hd__and2_1 _26463_ (.A(_23108_),
    .B(_23109_),
    .X(_23110_));
 sky130_fd_sc_hd__or2_1 _26464_ (.A(_23047_),
    .B(_23110_),
    .X(_23111_));
 sky130_fd_sc_hd__nand2_2 _26465_ (.A(_23047_),
    .B(_23110_),
    .Y(_23112_));
 sky130_fd_sc_hd__a311oi_4 _26466_ (.A1(_20617_),
    .A2(_21481_),
    .A3(_21486_),
    .B1(_21505_),
    .C1(_21484_),
    .Y(_23113_));
 sky130_fd_sc_hd__a221oi_1 _26467_ (.A1(_21506_),
    .A2(_21546_),
    .B1(_23111_),
    .B2(_23112_),
    .C1(_23113_),
    .Y(_23114_));
 sky130_fd_sc_hd__o211ai_4 _26468_ (.A1(_23113_),
    .A2(_21547_),
    .B1(_23112_),
    .C1(_23111_),
    .Y(_23115_));
 sky130_fd_sc_hd__and2b_4 _26469_ (.A_N(_23114_),
    .B(_23115_),
    .X(_23116_));
 sky130_fd_sc_hd__xnor2_4 _26470_ (.A(_23014_),
    .B(_23116_),
    .Y(_23118_));
 sky130_fd_sc_hd__xnor2_4 _26471_ (.A(_22924_),
    .B(_23118_),
    .Y(_23119_));
 sky130_fd_sc_hd__xor2_1 _26472_ (.A(_22922_),
    .B(_23119_),
    .X(_23120_));
 sky130_fd_sc_hd__o21ai_1 _26473_ (.A1(_21554_),
    .A2(_21658_),
    .B1(_23120_),
    .Y(_23121_));
 sky130_fd_sc_hd__a211o_1 _26474_ (.A1(_21555_),
    .A2(_21657_),
    .B1(_23120_),
    .C1(_21554_),
    .X(_23122_));
 sky130_fd_sc_hd__nand2_1 _26475_ (.A(_23121_),
    .B(_23122_),
    .Y(_23123_));
 sky130_fd_sc_hd__a211o_1 _26476_ (.A1(_21202_),
    .A2(_21217_),
    .B1(_21220_),
    .C1(_21255_),
    .X(_23124_));
 sky130_fd_sc_hd__nor2_1 _26477_ (.A(\delay_line[26][3] ),
    .B(_18488_),
    .Y(_23125_));
 sky130_fd_sc_hd__and2_1 _26478_ (.A(_16009_),
    .B(_18488_),
    .X(_23126_));
 sky130_fd_sc_hd__o21ai_2 _26479_ (.A1(_23125_),
    .A2(_23126_),
    .B1(_24347_),
    .Y(_23127_));
 sky130_fd_sc_hd__nand2_1 _26480_ (.A(_16009_),
    .B(_18486_),
    .Y(_23129_));
 sky130_fd_sc_hd__nand3b_2 _26481_ (.A_N(_23125_),
    .B(_23129_),
    .C(_18485_),
    .Y(_23130_));
 sky130_fd_sc_hd__o2bb2ai_1 _26482_ (.A1_N(_23127_),
    .A2_N(_23130_),
    .B1(_21223_),
    .B2(_06480_),
    .Y(_23131_));
 sky130_fd_sc_hd__o211ai_4 _26483_ (.A1(_18487_),
    .A2(_18489_),
    .B1(_16020_),
    .C1(_06590_),
    .Y(_23132_));
 sky130_fd_sc_hd__a22oi_1 _26484_ (.A1(_01172_),
    .A2(_21225_),
    .B1(_23131_),
    .B2(_23132_),
    .Y(_23133_));
 sky130_fd_sc_hd__or3b_2 _26485_ (.A(_16020_),
    .B(_06469_),
    .C_N(_19266_),
    .X(_23134_));
 sky130_fd_sc_hd__a22oi_4 _26486_ (.A1(_16020_),
    .A2(_06590_),
    .B1(_23127_),
    .B2(_23130_),
    .Y(_23135_));
 sky130_fd_sc_hd__nor2_1 _26487_ (.A(_23134_),
    .B(_23135_),
    .Y(_23136_));
 sky130_fd_sc_hd__o2bb2ai_1 _26488_ (.A1_N(_19263_),
    .A2_N(_21224_),
    .B1(_23133_),
    .B2(_23136_),
    .Y(_23137_));
 sky130_fd_sc_hd__nand4_2 _26489_ (.A(_06480_),
    .B(_23131_),
    .C(_19263_),
    .D(_16031_),
    .Y(_23138_));
 sky130_fd_sc_hd__clkbuf_2 _26490_ (.A(\delay_line[26][8] ),
    .X(_23140_));
 sky130_fd_sc_hd__inv_2 _26491_ (.A(_23140_),
    .Y(_23141_));
 sky130_fd_sc_hd__a21oi_2 _26492_ (.A1(_23137_),
    .A2(_23138_),
    .B1(_23141_),
    .Y(_23142_));
 sky130_fd_sc_hd__and3_1 _26493_ (.A(_23141_),
    .B(_23137_),
    .C(_23138_),
    .X(_23143_));
 sky130_fd_sc_hd__or4_1 _26494_ (.A(_21229_),
    .B(_21231_),
    .C(_23142_),
    .D(_23143_),
    .X(_23144_));
 sky130_fd_sc_hd__o22ai_4 _26495_ (.A1(_21229_),
    .A2(_21231_),
    .B1(_23142_),
    .B2(_23143_),
    .Y(_23145_));
 sky130_fd_sc_hd__nand2_1 _26496_ (.A(_23144_),
    .B(_23145_),
    .Y(_23146_));
 sky130_fd_sc_hd__clkbuf_2 _26497_ (.A(_20379_),
    .X(_23147_));
 sky130_fd_sc_hd__nor2_1 _26498_ (.A(_21235_),
    .B(_23147_),
    .Y(_23148_));
 sky130_fd_sc_hd__a21boi_1 _26499_ (.A1(_21236_),
    .A2(_21242_),
    .B1_N(_01205_),
    .Y(_23149_));
 sky130_fd_sc_hd__buf_1 _26500_ (.A(_21239_),
    .X(_23151_));
 sky130_fd_sc_hd__nor2_1 _26501_ (.A(\delay_line[27][7] ),
    .B(net331),
    .Y(_23152_));
 sky130_fd_sc_hd__nand2_1 _26502_ (.A(_20373_),
    .B(net331),
    .Y(_23153_));
 sky130_fd_sc_hd__nand3b_1 _26503_ (.A_N(_23152_),
    .B(_23153_),
    .C(_21240_),
    .Y(_23154_));
 sky130_fd_sc_hd__and2_2 _26504_ (.A(\delay_line[27][7] ),
    .B(net331),
    .X(_23155_));
 sky130_fd_sc_hd__o21ai_1 _26505_ (.A1(_23152_),
    .A2(_23155_),
    .B1(_21238_),
    .Y(_23156_));
 sky130_fd_sc_hd__nand2_1 _26506_ (.A(_23154_),
    .B(_23156_),
    .Y(_23157_));
 sky130_fd_sc_hd__clkbuf_2 _26507_ (.A(net331),
    .X(_23158_));
 sky130_fd_sc_hd__nor2_1 _26508_ (.A(_23158_),
    .B(_23151_),
    .Y(_23159_));
 sky130_fd_sc_hd__a211o_1 _26509_ (.A1(_23151_),
    .A2(_23157_),
    .B1(_23159_),
    .C1(_16206_),
    .X(_23160_));
 sky130_fd_sc_hd__clkbuf_2 _26510_ (.A(_23154_),
    .X(_23162_));
 sky130_fd_sc_hd__a21boi_1 _26511_ (.A1(_23162_),
    .A2(_23156_),
    .B1_N(_23151_),
    .Y(_23163_));
 sky130_fd_sc_hd__o21ai_1 _26512_ (.A1(_23163_),
    .A2(_23159_),
    .B1(_16206_),
    .Y(_23164_));
 sky130_fd_sc_hd__o211ai_2 _26513_ (.A1(_23148_),
    .A2(_23149_),
    .B1(_23160_),
    .C1(_23164_),
    .Y(_23165_));
 sky130_fd_sc_hd__a211o_1 _26514_ (.A1(_23160_),
    .A2(_23164_),
    .B1(_23148_),
    .C1(_23149_),
    .X(_23166_));
 sky130_fd_sc_hd__nand2_1 _26515_ (.A(_23165_),
    .B(_23166_),
    .Y(_23167_));
 sky130_fd_sc_hd__o211ai_2 _26516_ (.A1(_20374_),
    .A2(_20382_),
    .B1(_21243_),
    .C1(_21244_),
    .Y(_23168_));
 sky130_fd_sc_hd__o21ai_1 _26517_ (.A1(_21246_),
    .A2(_20389_),
    .B1(_23168_),
    .Y(_23169_));
 sky130_fd_sc_hd__xnor2_1 _26518_ (.A(_23167_),
    .B(_23169_),
    .Y(_23170_));
 sky130_fd_sc_hd__o32ai_4 _26519_ (.A1(_20390_),
    .A2(_21245_),
    .A3(_21246_),
    .B1(_21250_),
    .B2(_20394_),
    .Y(_23171_));
 sky130_fd_sc_hd__xnor2_2 _26520_ (.A(_23170_),
    .B(_23171_),
    .Y(_23173_));
 sky130_fd_sc_hd__xor2_1 _26521_ (.A(_23146_),
    .B(_23173_),
    .X(_23174_));
 sky130_fd_sc_hd__and3b_1 _26522_ (.A_N(_21204_),
    .B(_20410_),
    .C(_19304_),
    .X(_23175_));
 sky130_fd_sc_hd__a31o_1 _26523_ (.A1(_21203_),
    .A2(_21205_),
    .A3(_06414_),
    .B1(_23175_),
    .X(_23176_));
 sky130_fd_sc_hd__clkbuf_2 _26524_ (.A(\delay_line[28][8] ),
    .X(_23177_));
 sky130_fd_sc_hd__clkbuf_2 _26525_ (.A(\delay_line[28][9] ),
    .X(_23178_));
 sky130_fd_sc_hd__inv_2 _26526_ (.A(\delay_line[28][9] ),
    .Y(_23179_));
 sky130_fd_sc_hd__nand3_1 _26527_ (.A(_23179_),
    .B(\delay_line[28][8] ),
    .C(_20410_),
    .Y(_23180_));
 sky130_fd_sc_hd__nand3b_1 _26528_ (.A_N(_20410_),
    .B(_21204_),
    .C(\delay_line[28][9] ),
    .Y(_23181_));
 sky130_fd_sc_hd__o2111ai_2 _26529_ (.A1(_23177_),
    .A2(_23178_),
    .B1(_15965_),
    .C1(_23180_),
    .D1(_23181_),
    .Y(_23182_));
 sky130_fd_sc_hd__o211ai_1 _26530_ (.A1(_23177_),
    .A2(_23178_),
    .B1(_23180_),
    .C1(_23181_),
    .Y(_23184_));
 sky130_fd_sc_hd__nand2_1 _26531_ (.A(_20428_),
    .B(_23184_),
    .Y(_23185_));
 sky130_fd_sc_hd__nand3_1 _26532_ (.A(_23176_),
    .B(_23182_),
    .C(_23185_),
    .Y(_23186_));
 sky130_fd_sc_hd__a21o_1 _26533_ (.A1(_23182_),
    .A2(_23185_),
    .B1(_23176_),
    .X(_23187_));
 sky130_fd_sc_hd__a21oi_1 _26534_ (.A1(_23186_),
    .A2(_23187_),
    .B1(_06425_),
    .Y(_23188_));
 sky130_fd_sc_hd__and3_1 _26535_ (.A(_23187_),
    .B(_06425_),
    .C(_23186_),
    .X(_23189_));
 sky130_fd_sc_hd__nand3_1 _26536_ (.A(_21209_),
    .B(_21210_),
    .C(_01128_),
    .Y(_23190_));
 sky130_fd_sc_hd__o211ai_1 _26537_ (.A1(_23188_),
    .A2(_23189_),
    .B1(_21210_),
    .C1(_23190_),
    .Y(_23191_));
 sky130_fd_sc_hd__a211o_1 _26538_ (.A1(_21210_),
    .A2(_23190_),
    .B1(_23188_),
    .C1(_23189_),
    .X(_23192_));
 sky130_fd_sc_hd__nand2_2 _26539_ (.A(_23191_),
    .B(_23192_),
    .Y(_23193_));
 sky130_fd_sc_hd__xor2_4 _26540_ (.A(net171),
    .B(_23193_),
    .X(_23195_));
 sky130_fd_sc_hd__a21oi_4 _26541_ (.A1(_21202_),
    .A2(_21217_),
    .B1(_21218_),
    .Y(_23196_));
 sky130_fd_sc_hd__xor2_4 _26542_ (.A(_23195_),
    .B(_23196_),
    .X(_23197_));
 sky130_fd_sc_hd__or2_1 _26543_ (.A(_23174_),
    .B(_23197_),
    .X(_23198_));
 sky130_fd_sc_hd__nand2_1 _26544_ (.A(_23174_),
    .B(_23197_),
    .Y(_23199_));
 sky130_fd_sc_hd__nand2_1 _26545_ (.A(_23198_),
    .B(_23199_),
    .Y(_23200_));
 sky130_fd_sc_hd__and3_1 _26546_ (.A(_21254_),
    .B(_23124_),
    .C(_23200_),
    .X(_23201_));
 sky130_fd_sc_hd__inv_2 _26547_ (.A(_23201_),
    .Y(_23202_));
 sky130_fd_sc_hd__a21o_2 _26548_ (.A1(_21254_),
    .A2(_23124_),
    .B1(_23200_),
    .X(_23203_));
 sky130_fd_sc_hd__nand3_2 _26549_ (.A(_22226_),
    .B(_21287_),
    .C(_21286_),
    .Y(_23204_));
 sky130_fd_sc_hd__buf_1 _26550_ (.A(\delay_line[31][9] ),
    .X(_23206_));
 sky130_fd_sc_hd__inv_2 _26551_ (.A(_23206_),
    .Y(_23207_));
 sky130_fd_sc_hd__nor2_1 _26552_ (.A(_21264_),
    .B(_23206_),
    .Y(_23208_));
 sky130_fd_sc_hd__nand2_1 _26553_ (.A(_21264_),
    .B(_23206_),
    .Y(_23209_));
 sky130_fd_sc_hd__nand3b_2 _26554_ (.A_N(_23208_),
    .B(_23209_),
    .C(_20313_),
    .Y(_23210_));
 sky130_fd_sc_hd__o2111ai_4 _26555_ (.A1(_20313_),
    .A2(_23207_),
    .B1(_21269_),
    .C1(_21274_),
    .D1(_23210_),
    .Y(_23211_));
 sky130_fd_sc_hd__clkbuf_2 _26556_ (.A(_20308_),
    .X(_23212_));
 sky130_fd_sc_hd__clkbuf_2 _26557_ (.A(\delay_line[31][9] ),
    .X(_23213_));
 sky130_fd_sc_hd__nand2_1 _26558_ (.A(_23212_),
    .B(_23213_),
    .Y(_23214_));
 sky130_fd_sc_hd__a22o_1 _26559_ (.A1(_21269_),
    .A2(_21274_),
    .B1(_23210_),
    .B2(_23214_),
    .X(_23215_));
 sky130_fd_sc_hd__xor2_1 _26560_ (.A(_20317_),
    .B(_06216_),
    .X(_23217_));
 sky130_fd_sc_hd__a21o_1 _26561_ (.A1(_23211_),
    .A2(_23215_),
    .B1(_23217_),
    .X(_23218_));
 sky130_fd_sc_hd__nand3_1 _26562_ (.A(_23217_),
    .B(_23211_),
    .C(_23215_),
    .Y(_23219_));
 sky130_fd_sc_hd__nand4_1 _26563_ (.A(_21276_),
    .B(_21281_),
    .C(_23218_),
    .D(_23219_),
    .Y(_23220_));
 sky130_fd_sc_hd__a22o_2 _26564_ (.A1(_21276_),
    .A2(_21281_),
    .B1(_23218_),
    .B2(_23219_),
    .X(_23221_));
 sky130_fd_sc_hd__nand3b_2 _26565_ (.A_N(_21283_),
    .B(_23220_),
    .C(_23221_),
    .Y(_23222_));
 sky130_fd_sc_hd__nand2_1 _26566_ (.A(_23220_),
    .B(_23221_),
    .Y(_23223_));
 sky130_fd_sc_hd__nand2_1 _26567_ (.A(_21283_),
    .B(_23223_),
    .Y(_23224_));
 sky130_fd_sc_hd__nand2_1 _26568_ (.A(_23222_),
    .B(_23224_),
    .Y(_23225_));
 sky130_fd_sc_hd__a21o_1 _26569_ (.A1(_21288_),
    .A2(_23204_),
    .B1(_23225_),
    .X(_23226_));
 sky130_fd_sc_hd__nand3_1 _26570_ (.A(_21288_),
    .B(_23204_),
    .C(_23225_),
    .Y(_23228_));
 sky130_fd_sc_hd__a31o_1 _26571_ (.A1(_21292_),
    .A2(_21294_),
    .A3(_23204_),
    .B1(_21296_),
    .X(_23229_));
 sky130_fd_sc_hd__and3_2 _26572_ (.A(_23226_),
    .B(_23228_),
    .C(_23229_),
    .X(_23230_));
 sky130_fd_sc_hd__a21oi_2 _26573_ (.A1(_23226_),
    .A2(_23228_),
    .B1(_23229_),
    .Y(_23231_));
 sky130_fd_sc_hd__and2b_1 _26574_ (.A_N(_15646_),
    .B(_21300_),
    .X(_23232_));
 sky130_fd_sc_hd__nand2_1 _26575_ (.A(_18450_),
    .B(\delay_line[29][7] ),
    .Y(_23233_));
 sky130_fd_sc_hd__or2_1 _26576_ (.A(\delay_line[29][7] ),
    .B(_18450_),
    .X(_23234_));
 sky130_fd_sc_hd__nand2_1 _26577_ (.A(_23233_),
    .B(_23234_),
    .Y(_23235_));
 sky130_fd_sc_hd__o21a_1 _26578_ (.A1(_23232_),
    .A2(_21303_),
    .B1(_23235_),
    .X(_23236_));
 sky130_fd_sc_hd__and4bb_1 _26579_ (.A_N(_23232_),
    .B_N(_21303_),
    .C(_23233_),
    .D(_23234_),
    .X(_23237_));
 sky130_fd_sc_hd__nor3_1 _26580_ (.A(net235),
    .B(_23236_),
    .C(_23237_),
    .Y(_23239_));
 sky130_fd_sc_hd__o21a_1 _26581_ (.A1(_23236_),
    .A2(_23237_),
    .B1(_21304_),
    .X(_23240_));
 sky130_fd_sc_hd__nand2_1 _26582_ (.A(_21331_),
    .B(_21335_),
    .Y(_23241_));
 sky130_fd_sc_hd__a31o_1 _26583_ (.A1(_21322_),
    .A2(_21317_),
    .A3(_21320_),
    .B1(_21325_),
    .X(_23242_));
 sky130_fd_sc_hd__or3b_1 _26584_ (.A(_06315_),
    .B(_20343_),
    .C_N(_01018_),
    .X(_23243_));
 sky130_fd_sc_hd__inv_2 _26585_ (.A(_21312_),
    .Y(_23244_));
 sky130_fd_sc_hd__o211a_1 _26586_ (.A1(_21318_),
    .A2(_21319_),
    .B1(_21312_),
    .C1(_21314_),
    .X(_23245_));
 sky130_fd_sc_hd__clkbuf_2 _26587_ (.A(_21308_),
    .X(_23246_));
 sky130_fd_sc_hd__or2_1 _26588_ (.A(\delay_line[30][8] ),
    .B(\delay_line[30][9] ),
    .X(_23247_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26589_ (.A(\delay_line[30][9] ),
    .X(_23248_));
 sky130_fd_sc_hd__nand2_2 _26590_ (.A(\delay_line[30][8] ),
    .B(_23248_),
    .Y(_23250_));
 sky130_fd_sc_hd__nand2_1 _26591_ (.A(\delay_line[30][4] ),
    .B(\delay_line[30][6] ),
    .Y(_23251_));
 sky130_fd_sc_hd__nand2_1 _26592_ (.A(_20342_),
    .B(_19328_),
    .Y(_23252_));
 sky130_fd_sc_hd__nand4_1 _26593_ (.A(_23247_),
    .B(_23250_),
    .C(_23251_),
    .D(_23252_),
    .Y(_23253_));
 sky130_fd_sc_hd__clkbuf_2 _26594_ (.A(_23253_),
    .X(_23254_));
 sky130_fd_sc_hd__nor2_1 _26595_ (.A(_21307_),
    .B(_23248_),
    .Y(_23255_));
 sky130_fd_sc_hd__and2_1 _26596_ (.A(\delay_line[30][8] ),
    .B(_23248_),
    .X(_23256_));
 sky130_fd_sc_hd__and2_1 _26597_ (.A(_20340_),
    .B(\delay_line[30][6] ),
    .X(_23257_));
 sky130_fd_sc_hd__nor2_1 _26598_ (.A(_15569_),
    .B(_19335_),
    .Y(_23258_));
 sky130_fd_sc_hd__o22ai_2 _26599_ (.A1(_23255_),
    .A2(_23256_),
    .B1(_23257_),
    .B2(_23258_),
    .Y(_23259_));
 sky130_fd_sc_hd__a22o_1 _26600_ (.A1(_18452_),
    .A2(_23246_),
    .B1(_23254_),
    .B2(_23259_),
    .X(_23261_));
 sky130_fd_sc_hd__o2bb2a_1 _26601_ (.A1_N(_01007_),
    .A2_N(_06293_),
    .B1(_19332_),
    .B2(_19333_),
    .X(_23262_));
 sky130_fd_sc_hd__and3_2 _26602_ (.A(_24611_),
    .B(_01007_),
    .C(_06293_),
    .X(_23263_));
 sky130_fd_sc_hd__nor2_1 _26603_ (.A(_23262_),
    .B(_23263_),
    .Y(_23264_));
 sky130_fd_sc_hd__nand4_1 _26604_ (.A(_23246_),
    .B(_23254_),
    .C(_23259_),
    .D(_18452_),
    .Y(_23265_));
 sky130_fd_sc_hd__nand3_1 _26605_ (.A(_23261_),
    .B(_23264_),
    .C(_23265_),
    .Y(_23266_));
 sky130_fd_sc_hd__and3b_1 _26606_ (.A_N(_21309_),
    .B(_23253_),
    .C(_23259_),
    .X(_23267_));
 sky130_fd_sc_hd__clkbuf_2 _26607_ (.A(_21310_),
    .X(_23268_));
 sky130_fd_sc_hd__clkbuf_2 _26608_ (.A(_21307_),
    .X(_23269_));
 sky130_fd_sc_hd__o2bb2a_1 _26609_ (.A1_N(_23254_),
    .A2_N(_23259_),
    .B1(_23268_),
    .B2(_23269_),
    .X(_23270_));
 sky130_fd_sc_hd__o22ai_2 _26610_ (.A1(_23262_),
    .A2(_23263_),
    .B1(_23267_),
    .B2(_23270_),
    .Y(_23272_));
 sky130_fd_sc_hd__o211a_2 _26611_ (.A1(_23244_),
    .A2(_23245_),
    .B1(_23266_),
    .C1(_23272_),
    .X(_23273_));
 sky130_fd_sc_hd__nand2_1 _26612_ (.A(_21312_),
    .B(_21320_),
    .Y(_23274_));
 sky130_fd_sc_hd__a21oi_1 _26613_ (.A1(_23266_),
    .A2(_23272_),
    .B1(_23274_),
    .Y(_23275_));
 sky130_fd_sc_hd__nor3_2 _26614_ (.A(_23243_),
    .B(_23273_),
    .C(_23275_),
    .Y(_23276_));
 sky130_fd_sc_hd__o21a_1 _26615_ (.A1(_23273_),
    .A2(_23275_),
    .B1(_23243_),
    .X(_23277_));
 sky130_fd_sc_hd__nor2_1 _26616_ (.A(_23276_),
    .B(_23277_),
    .Y(_23278_));
 sky130_fd_sc_hd__xor2_1 _26617_ (.A(_23242_),
    .B(_23278_),
    .X(_23279_));
 sky130_fd_sc_hd__or2_1 _26618_ (.A(_23241_),
    .B(_23279_),
    .X(_23280_));
 sky130_fd_sc_hd__nand2_1 _26619_ (.A(_23279_),
    .B(_23241_),
    .Y(_23281_));
 sky130_fd_sc_hd__nand2_1 _26620_ (.A(_23280_),
    .B(_23281_),
    .Y(_23283_));
 sky130_fd_sc_hd__a311o_1 _26621_ (.A1(_22292_),
    .A2(_01040_),
    .A3(_20357_),
    .B1(_20359_),
    .C1(_19345_),
    .X(_23284_));
 sky130_fd_sc_hd__o21ai_1 _26622_ (.A1(_23284_),
    .A2(_21337_),
    .B1(_21340_),
    .Y(_23285_));
 sky130_fd_sc_hd__xor2_1 _26623_ (.A(_23283_),
    .B(_23285_),
    .X(_23286_));
 sky130_fd_sc_hd__o21ai_1 _26624_ (.A1(_23239_),
    .A2(_23240_),
    .B1(_23286_),
    .Y(_23287_));
 sky130_fd_sc_hd__or3_1 _26625_ (.A(_23239_),
    .B(_23240_),
    .C(_23286_),
    .X(_23288_));
 sky130_fd_sc_hd__nand2_1 _26626_ (.A(_23287_),
    .B(_23288_),
    .Y(_23289_));
 sky130_fd_sc_hd__or3_4 _26627_ (.A(_23230_),
    .B(_23231_),
    .C(_23289_),
    .X(_23290_));
 sky130_fd_sc_hd__o21ai_4 _26628_ (.A1(_23230_),
    .A2(_23231_),
    .B1(_23289_),
    .Y(_23291_));
 sky130_fd_sc_hd__a22oi_4 _26629_ (.A1(_23202_),
    .A2(_23203_),
    .B1(_23290_),
    .B2(_23291_),
    .Y(_23292_));
 sky130_fd_sc_hd__nand4_4 _26630_ (.A(_23202_),
    .B(_23203_),
    .C(_23290_),
    .D(_23291_),
    .Y(_23294_));
 sky130_fd_sc_hd__inv_2 _26631_ (.A(_23294_),
    .Y(_23295_));
 sky130_fd_sc_hd__o21a_1 _26632_ (.A1(_21557_),
    .A2(_21654_),
    .B1(_21655_),
    .X(_23296_));
 sky130_fd_sc_hd__o21ai_1 _26633_ (.A1(_23292_),
    .A2(_23295_),
    .B1(_23296_),
    .Y(_23297_));
 sky130_fd_sc_hd__or3_1 _26634_ (.A(_23296_),
    .B(_23292_),
    .C(_23295_),
    .X(_23298_));
 sky130_fd_sc_hd__nand2_1 _26635_ (.A(_23297_),
    .B(_23298_),
    .Y(_23299_));
 sky130_fd_sc_hd__a21oi_4 _26636_ (.A1(_21348_),
    .A2(_21258_),
    .B1(_21257_),
    .Y(_23300_));
 sky130_fd_sc_hd__xnor2_1 _26637_ (.A(_23299_),
    .B(_23300_),
    .Y(_23301_));
 sky130_fd_sc_hd__or2_1 _26638_ (.A(_23123_),
    .B(_23301_),
    .X(_23302_));
 sky130_fd_sc_hd__nand2_1 _26639_ (.A(_23123_),
    .B(_23301_),
    .Y(_23303_));
 sky130_fd_sc_hd__and2_1 _26640_ (.A(_23302_),
    .B(_23303_),
    .X(_23305_));
 sky130_fd_sc_hd__xnor2_1 _26641_ (.A(_22810_),
    .B(_23305_),
    .Y(_23306_));
 sky130_fd_sc_hd__a21o_1 _26642_ (.A1(_21352_),
    .A2(_21201_),
    .B1(_21350_),
    .X(_23307_));
 sky130_fd_sc_hd__a21o_1 _26643_ (.A1(_21187_),
    .A2(_21188_),
    .B1(_21186_),
    .X(_23308_));
 sky130_fd_sc_hd__nand2_1 _26644_ (.A(_21108_),
    .B(_21109_),
    .Y(_23309_));
 sky130_fd_sc_hd__a21boi_2 _26645_ (.A1(_20749_),
    .A2(_21104_),
    .B1_N(_21105_),
    .Y(_23310_));
 sky130_fd_sc_hd__nor2_1 _26646_ (.A(\delay_line[34][7] ),
    .B(\delay_line[34][9] ),
    .Y(_23311_));
 sky130_fd_sc_hd__buf_1 _26647_ (.A(\delay_line[34][9] ),
    .X(_23312_));
 sky130_fd_sc_hd__nand2_1 _26648_ (.A(_20743_),
    .B(_23312_),
    .Y(_23313_));
 sky130_fd_sc_hd__nand3b_1 _26649_ (.A_N(_23311_),
    .B(_21084_),
    .C(_23313_),
    .Y(_23314_));
 sky130_fd_sc_hd__buf_1 _26650_ (.A(_23314_),
    .X(_23316_));
 sky130_fd_sc_hd__and2_1 _26651_ (.A(_20743_),
    .B(_23312_),
    .X(_23317_));
 sky130_fd_sc_hd__o21ai_2 _26652_ (.A1(_23317_),
    .A2(_23311_),
    .B1(_21090_),
    .Y(_23318_));
 sky130_fd_sc_hd__nor2_1 _26653_ (.A(_18633_),
    .B(_19553_),
    .Y(_23319_));
 sky130_fd_sc_hd__and2_1 _26654_ (.A(_18631_),
    .B(_19549_),
    .X(_23320_));
 sky130_fd_sc_hd__nor2_1 _26655_ (.A(_23319_),
    .B(_23320_),
    .Y(_23321_));
 sky130_fd_sc_hd__a21boi_1 _26656_ (.A1(_23316_),
    .A2(_23318_),
    .B1_N(_23321_),
    .Y(_23322_));
 sky130_fd_sc_hd__o211ai_1 _26657_ (.A1(_23319_),
    .A2(_23320_),
    .B1(_23316_),
    .C1(_23318_),
    .Y(_23323_));
 sky130_fd_sc_hd__a21boi_1 _26658_ (.A1(_21088_),
    .A2(_21089_),
    .B1_N(_21091_),
    .Y(_23324_));
 sky130_fd_sc_hd__nand3b_1 _26659_ (.A_N(_23322_),
    .B(_23323_),
    .C(_23324_),
    .Y(_23325_));
 sky130_fd_sc_hd__nand3_1 _26660_ (.A(_23318_),
    .B(_23321_),
    .C(_23316_),
    .Y(_23327_));
 sky130_fd_sc_hd__a21o_1 _26661_ (.A1(_23314_),
    .A2(_23318_),
    .B1(_23321_),
    .X(_23328_));
 sky130_fd_sc_hd__nand3b_1 _26662_ (.A_N(_23324_),
    .B(_23327_),
    .C(_23328_),
    .Y(_23329_));
 sky130_fd_sc_hd__xor2_1 _26663_ (.A(_02249_),
    .B(_21097_),
    .X(_23330_));
 sky130_fd_sc_hd__a21o_1 _26664_ (.A1(_23325_),
    .A2(_23329_),
    .B1(_23330_),
    .X(_23331_));
 sky130_fd_sc_hd__nand3_1 _26665_ (.A(_23325_),
    .B(_23329_),
    .C(_23330_),
    .Y(_23332_));
 sky130_fd_sc_hd__a21oi_1 _26666_ (.A1(_21092_),
    .A2(_21093_),
    .B1(_21094_),
    .Y(_23333_));
 sky130_fd_sc_hd__o21ai_1 _26667_ (.A1(_21100_),
    .A2(_23333_),
    .B1(_21096_),
    .Y(_23334_));
 sky130_fd_sc_hd__a21o_1 _26668_ (.A1(_23331_),
    .A2(_23332_),
    .B1(_23334_),
    .X(_23335_));
 sky130_fd_sc_hd__nand3_1 _26669_ (.A(_23334_),
    .B(_23331_),
    .C(_23332_),
    .Y(_23336_));
 sky130_fd_sc_hd__and3_1 _26670_ (.A(_23335_),
    .B(_23336_),
    .C(_21098_),
    .X(_23338_));
 sky130_fd_sc_hd__a21oi_1 _26671_ (.A1(_23335_),
    .A2(_23336_),
    .B1(_21098_),
    .Y(_23339_));
 sky130_fd_sc_hd__or2_1 _26672_ (.A(_23338_),
    .B(_23339_),
    .X(_23340_));
 sky130_fd_sc_hd__xor2_1 _26673_ (.A(_23310_),
    .B(_23340_),
    .X(_23341_));
 sky130_fd_sc_hd__xor2_1 _26674_ (.A(_23309_),
    .B(_23341_),
    .X(_23342_));
 sky130_fd_sc_hd__and3_1 _26675_ (.A(_21169_),
    .B(_21170_),
    .C(_21171_),
    .X(_23343_));
 sky130_fd_sc_hd__a21oi_2 _26676_ (.A1(_21169_),
    .A2(_21170_),
    .B1(_21171_),
    .Y(_23344_));
 sky130_fd_sc_hd__nor2_1 _26677_ (.A(_22523_),
    .B(_23344_),
    .Y(_23345_));
 sky130_fd_sc_hd__nand2_1 _26678_ (.A(_21166_),
    .B(_21169_),
    .Y(_23346_));
 sky130_fd_sc_hd__nor2_1 _26679_ (.A(\delay_line[33][8] ),
    .B(\delay_line[33][9] ),
    .Y(_23347_));
 sky130_fd_sc_hd__nand2_1 _26680_ (.A(_21161_),
    .B(\delay_line[33][9] ),
    .Y(_23349_));
 sky130_fd_sc_hd__inv_2 _26681_ (.A(\delay_line[33][4] ),
    .Y(_23350_));
 sky130_fd_sc_hd__nand2_1 _26682_ (.A(_23350_),
    .B(_18650_),
    .Y(_23351_));
 sky130_fd_sc_hd__buf_1 _26683_ (.A(net312),
    .X(_23352_));
 sky130_fd_sc_hd__nand2_1 _26684_ (.A(_17822_),
    .B(_23352_),
    .Y(_23353_));
 sky130_fd_sc_hd__nand4b_1 _26685_ (.A_N(_23347_),
    .B(_23349_),
    .C(_23351_),
    .D(_23353_),
    .Y(_23354_));
 sky130_fd_sc_hd__clkbuf_2 _26686_ (.A(_23354_),
    .X(_23355_));
 sky130_fd_sc_hd__inv_2 _26687_ (.A(_21161_),
    .Y(_23356_));
 sky130_fd_sc_hd__clkbuf_2 _26688_ (.A(_23356_),
    .X(_23357_));
 sky130_fd_sc_hd__and2_1 _26689_ (.A(_21161_),
    .B(\delay_line[33][9] ),
    .X(_23358_));
 sky130_fd_sc_hd__nor2_1 _26690_ (.A(_17822_),
    .B(_23352_),
    .Y(_23360_));
 sky130_fd_sc_hd__nor2_1 _26691_ (.A(_23350_),
    .B(_18650_),
    .Y(_23361_));
 sky130_fd_sc_hd__o22ai_2 _26692_ (.A1(_23347_),
    .A2(_23358_),
    .B1(_23360_),
    .B2(_23361_),
    .Y(_23362_));
 sky130_fd_sc_hd__nand4_2 _26693_ (.A(_23355_),
    .B(_17823_),
    .C(_23357_),
    .D(_23362_),
    .Y(_23363_));
 sky130_fd_sc_hd__clkbuf_2 _26694_ (.A(_23356_),
    .X(_23364_));
 sky130_fd_sc_hd__a22o_1 _26695_ (.A1(_17823_),
    .A2(_23364_),
    .B1(_23354_),
    .B2(_23362_),
    .X(_23365_));
 sky130_fd_sc_hd__inv_2 _26696_ (.A(net313),
    .Y(_23366_));
 sky130_fd_sc_hd__buf_2 _26697_ (.A(_23366_),
    .X(_23367_));
 sky130_fd_sc_hd__o21a_1 _26698_ (.A1(_19571_),
    .A2(_19572_),
    .B1(_05337_),
    .X(_23368_));
 sky130_fd_sc_hd__a21oi_1 _26699_ (.A1(_00568_),
    .A2(_23367_),
    .B1(_23368_),
    .Y(_23369_));
 sky130_fd_sc_hd__a21o_1 _26700_ (.A1(_23363_),
    .A2(_23365_),
    .B1(_23369_),
    .X(_23371_));
 sky130_fd_sc_hd__nand3_1 _26701_ (.A(_23363_),
    .B(_23365_),
    .C(_23369_),
    .Y(_23372_));
 sky130_fd_sc_hd__nand3_1 _26702_ (.A(_23371_),
    .B(_21164_),
    .C(_23372_),
    .Y(_23373_));
 sky130_fd_sc_hd__a21o_1 _26703_ (.A1(_23372_),
    .A2(_23371_),
    .B1(_21164_),
    .X(_23374_));
 sky130_fd_sc_hd__and3_1 _26704_ (.A(_23346_),
    .B(_23373_),
    .C(_23374_),
    .X(_23375_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26705_ (.A(_23373_),
    .X(_23376_));
 sky130_fd_sc_hd__a21oi_2 _26706_ (.A1(_23376_),
    .A2(_23374_),
    .B1(_23346_),
    .Y(_23377_));
 sky130_fd_sc_hd__nor2_1 _26707_ (.A(_23375_),
    .B(_23377_),
    .Y(_23378_));
 sky130_fd_sc_hd__o21ai_1 _26708_ (.A1(_23343_),
    .A2(_23345_),
    .B1(_23378_),
    .Y(_23379_));
 sky130_fd_sc_hd__o221ai_4 _26709_ (.A1(_22523_),
    .A2(_23344_),
    .B1(_23375_),
    .B2(_23377_),
    .C1(_21172_),
    .Y(_23380_));
 sky130_fd_sc_hd__o2bb2a_1 _26710_ (.A1_N(_23379_),
    .A2_N(_23380_),
    .B1(_20684_),
    .B2(_21176_),
    .X(_23382_));
 sky130_fd_sc_hd__o31a_1 _26711_ (.A1(_23343_),
    .A2(_23378_),
    .A3(_23345_),
    .B1(_21175_),
    .X(_23383_));
 sky130_fd_sc_hd__o2bb2ai_2 _26712_ (.A1_N(_24512_),
    .A2_N(_21144_),
    .B1(_21147_),
    .B2(_21146_),
    .Y(_23384_));
 sky130_fd_sc_hd__nand2_1 _26713_ (.A(_24523_),
    .B(_05304_),
    .Y(_23385_));
 sky130_fd_sc_hd__nand2_1 _26714_ (.A(_05249_),
    .B(_24457_),
    .Y(_23386_));
 sky130_fd_sc_hd__and3_1 _26715_ (.A(_23385_),
    .B(_23386_),
    .C(_19587_),
    .X(_23387_));
 sky130_fd_sc_hd__a21oi_1 _26716_ (.A1(_23385_),
    .A2(_23386_),
    .B1(_19587_),
    .Y(_23388_));
 sky130_fd_sc_hd__clkbuf_2 _26717_ (.A(\delay_line[32][9] ),
    .X(_23389_));
 sky130_fd_sc_hd__a21boi_1 _26718_ (.A1(_21115_),
    .A2(_23389_),
    .B1_N(_20686_),
    .Y(_23390_));
 sky130_fd_sc_hd__o21ai_1 _26719_ (.A1(_21116_),
    .A2(_23389_),
    .B1(_23390_),
    .Y(_23391_));
 sky130_fd_sc_hd__nand2_1 _26720_ (.A(_20690_),
    .B(_23389_),
    .Y(_23393_));
 sky130_fd_sc_hd__a21oi_2 _26721_ (.A1(_23391_),
    .A2(_23393_),
    .B1(_21112_),
    .Y(_23394_));
 sky130_fd_sc_hd__and3_1 _26722_ (.A(_21112_),
    .B(_23391_),
    .C(_23393_),
    .X(_23395_));
 sky130_fd_sc_hd__a21boi_1 _26723_ (.A1(_21118_),
    .A2(_21122_),
    .B1_N(_21121_),
    .Y(_23396_));
 sky130_fd_sc_hd__o21a_1 _26724_ (.A1(_23394_),
    .A2(_23395_),
    .B1(_23396_),
    .X(_23397_));
 sky130_fd_sc_hd__nor3_2 _26725_ (.A(_23394_),
    .B(_23395_),
    .C(_23396_),
    .Y(_23398_));
 sky130_fd_sc_hd__o22a_1 _26726_ (.A1(_23387_),
    .A2(_23388_),
    .B1(_23397_),
    .B2(_23398_),
    .X(_23399_));
 sky130_fd_sc_hd__or2_1 _26727_ (.A(_23387_),
    .B(_23388_),
    .X(_23400_));
 sky130_fd_sc_hd__nor3_2 _26728_ (.A(_23400_),
    .B(_23397_),
    .C(_23398_),
    .Y(_23401_));
 sky130_fd_sc_hd__a21oi_1 _26729_ (.A1(_20706_),
    .A2(_20710_),
    .B1(_21132_),
    .Y(_23402_));
 sky130_fd_sc_hd__a21oi_1 _26730_ (.A1(_02117_),
    .A2(_21133_),
    .B1(_23402_),
    .Y(_23404_));
 sky130_fd_sc_hd__nor3_1 _26731_ (.A(_23399_),
    .B(_23401_),
    .C(_23404_),
    .Y(_23405_));
 sky130_fd_sc_hd__o211a_1 _26732_ (.A1(_23399_),
    .A2(_23401_),
    .B1(_21130_),
    .C1(_21139_),
    .X(_23406_));
 sky130_fd_sc_hd__nor2_1 _26733_ (.A(_23405_),
    .B(_23406_),
    .Y(_23407_));
 sky130_fd_sc_hd__xnor2_1 _26734_ (.A(_21141_),
    .B(_23407_),
    .Y(_23408_));
 sky130_fd_sc_hd__xor2_1 _26735_ (.A(_23384_),
    .B(_23408_),
    .X(_23409_));
 sky130_fd_sc_hd__o21a_1 _26736_ (.A1(_21156_),
    .A2(_21157_),
    .B1(_23409_),
    .X(_23410_));
 sky130_fd_sc_hd__nand2_1 _26737_ (.A(_21145_),
    .B(_21151_),
    .Y(_23411_));
 sky130_fd_sc_hd__and3_1 _26738_ (.A(_24512_),
    .B(_21142_),
    .C(_21144_),
    .X(_23412_));
 sky130_fd_sc_hd__o22ai_2 _26739_ (.A1(_23411_),
    .A2(_23412_),
    .B1(_21152_),
    .B2(_21155_),
    .Y(_23413_));
 sky130_fd_sc_hd__nor2_1 _26740_ (.A(_23409_),
    .B(_23413_),
    .Y(_23415_));
 sky130_fd_sc_hd__or4_2 _26741_ (.A(_23382_),
    .B(_23383_),
    .C(_23410_),
    .D(_23415_),
    .X(_23416_));
 sky130_fd_sc_hd__o22a_1 _26742_ (.A1(_23382_),
    .A2(_23383_),
    .B1(_23410_),
    .B2(_23415_),
    .X(_23417_));
 sky130_fd_sc_hd__inv_2 _26743_ (.A(_23417_),
    .Y(_23418_));
 sky130_fd_sc_hd__nand2_1 _26744_ (.A(_23416_),
    .B(_23418_),
    .Y(_23419_));
 sky130_fd_sc_hd__xnor2_1 _26745_ (.A(_23342_),
    .B(_23419_),
    .Y(_23420_));
 sky130_fd_sc_hd__nand3_1 _26746_ (.A(_21344_),
    .B(_21346_),
    .C(_23420_),
    .Y(_23421_));
 sky130_fd_sc_hd__a21o_1 _26747_ (.A1(_21344_),
    .A2(_21346_),
    .B1(_23420_),
    .X(_23422_));
 sky130_fd_sc_hd__nand2_1 _26748_ (.A(_23421_),
    .B(_23422_),
    .Y(_23423_));
 sky130_fd_sc_hd__a21o_1 _26749_ (.A1(_21180_),
    .A2(_21182_),
    .B1(_23423_),
    .X(_23424_));
 sky130_fd_sc_hd__nand3_1 _26750_ (.A(_21180_),
    .B(_21182_),
    .C(_23423_),
    .Y(_23426_));
 sky130_fd_sc_hd__and2_1 _26751_ (.A(_23424_),
    .B(_23426_),
    .X(_23427_));
 sky130_fd_sc_hd__xnor2_1 _26752_ (.A(_23308_),
    .B(_23427_),
    .Y(_23428_));
 sky130_fd_sc_hd__clkbuf_2 _26753_ (.A(_20787_),
    .X(_23429_));
 sky130_fd_sc_hd__nand4_1 _26754_ (.A(_05568_),
    .B(_23429_),
    .C(_20786_),
    .D(_21006_),
    .Y(_23430_));
 sky130_fd_sc_hd__nor2_1 _26755_ (.A(_20787_),
    .B(net286),
    .Y(_23431_));
 sky130_fd_sc_hd__nand2_1 _26756_ (.A(_20787_),
    .B(net286),
    .Y(_23432_));
 sky130_fd_sc_hd__and2b_1 _26757_ (.A_N(_23431_),
    .B(_23432_),
    .X(_23433_));
 sky130_fd_sc_hd__buf_1 _26758_ (.A(\delay_line[38][7] ),
    .X(_23434_));
 sky130_fd_sc_hd__o211a_1 _26759_ (.A1(_21003_),
    .A2(net287),
    .B1(_23434_),
    .C1(_19649_),
    .X(_23435_));
 sky130_fd_sc_hd__a211oi_1 _26760_ (.A1(_21003_),
    .A2(net287),
    .B1(_23433_),
    .C1(_23435_),
    .Y(_23437_));
 sky130_fd_sc_hd__o21a_1 _26761_ (.A1(_21005_),
    .A2(_23435_),
    .B1(_23433_),
    .X(_23438_));
 sky130_fd_sc_hd__a211oi_2 _26762_ (.A1(_21012_),
    .A2(_23430_),
    .B1(_23437_),
    .C1(_23438_),
    .Y(_23439_));
 sky130_fd_sc_hd__o211a_1 _26763_ (.A1(_23438_),
    .A2(_23437_),
    .B1(_23430_),
    .C1(_21012_),
    .X(_23440_));
 sky130_fd_sc_hd__o21ba_1 _26764_ (.A1(_20801_),
    .A2(_20807_),
    .B1_N(_20996_),
    .X(_23441_));
 sky130_fd_sc_hd__nand2_1 _26765_ (.A(net282),
    .B(net281),
    .Y(_23442_));
 sky130_fd_sc_hd__buf_1 _26766_ (.A(\delay_line[39][9] ),
    .X(_23443_));
 sky130_fd_sc_hd__nor2_1 _26767_ (.A(net281),
    .B(_23443_),
    .Y(_23444_));
 sky130_fd_sc_hd__clkbuf_2 _26768_ (.A(_20987_),
    .X(_23445_));
 sky130_fd_sc_hd__inv_2 _26769_ (.A(\delay_line[39][9] ),
    .Y(_23446_));
 sky130_fd_sc_hd__nor2_1 _26770_ (.A(_23445_),
    .B(_23446_),
    .Y(_23448_));
 sky130_fd_sc_hd__or3_2 _26771_ (.A(_20986_),
    .B(_23444_),
    .C(_23448_),
    .X(_23449_));
 sky130_fd_sc_hd__o21ai_1 _26772_ (.A1(_23444_),
    .A2(_23448_),
    .B1(_20986_),
    .Y(_23450_));
 sky130_fd_sc_hd__nand2_2 _26773_ (.A(_23449_),
    .B(_23450_),
    .Y(_23451_));
 sky130_fd_sc_hd__a21oi_2 _26774_ (.A1(_23442_),
    .A2(_20989_),
    .B1(_23451_),
    .Y(_23452_));
 sky130_fd_sc_hd__a311oi_4 _26775_ (.A1(_20985_),
    .A2(_23442_),
    .A3(_23451_),
    .B1(_19662_),
    .C1(_23452_),
    .Y(_23453_));
 sky130_fd_sc_hd__and3_1 _26776_ (.A(_23442_),
    .B(_20989_),
    .C(_23451_),
    .X(_23454_));
 sky130_fd_sc_hd__o21a_1 _26777_ (.A1(_23452_),
    .A2(_23454_),
    .B1(_19662_),
    .X(_23455_));
 sky130_fd_sc_hd__nor2_1 _26778_ (.A(_23453_),
    .B(_23455_),
    .Y(_23456_));
 sky130_fd_sc_hd__or2_1 _26779_ (.A(_20992_),
    .B(_23456_),
    .X(_23457_));
 sky130_fd_sc_hd__o21a_1 _26780_ (.A1(_20992_),
    .A2(_20993_),
    .B1(_23456_),
    .X(_23459_));
 sky130_fd_sc_hd__o21ba_1 _26781_ (.A1(_20993_),
    .A2(_23457_),
    .B1_N(_23459_),
    .X(_23460_));
 sky130_fd_sc_hd__nor3_1 _26782_ (.A(_23441_),
    .B(_20999_),
    .C(_23460_),
    .Y(_23461_));
 sky130_fd_sc_hd__o21a_1 _26783_ (.A1(_23441_),
    .A2(_20999_),
    .B1(_23460_),
    .X(_23462_));
 sky130_fd_sc_hd__or4_1 _26784_ (.A(_23439_),
    .B(_23440_),
    .C(_23461_),
    .D(_23462_),
    .X(_23463_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26785_ (.A(_21019_),
    .X(_23464_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26786_ (.A(\delay_line[40][9] ),
    .X(_23465_));
 sky130_fd_sc_hd__a21oi_1 _26787_ (.A1(_21017_),
    .A2(_23464_),
    .B1(_23465_),
    .Y(_23466_));
 sky130_fd_sc_hd__and3_1 _26788_ (.A(_21017_),
    .B(_23464_),
    .C(\delay_line[40][9] ),
    .X(_23467_));
 sky130_fd_sc_hd__nor3_1 _26789_ (.A(_19633_),
    .B(_23466_),
    .C(_23467_),
    .Y(_23468_));
 sky130_fd_sc_hd__o21a_1 _26790_ (.A1(_23466_),
    .A2(_23467_),
    .B1(_19633_),
    .X(_23470_));
 sky130_fd_sc_hd__o211a_1 _26791_ (.A1(net272),
    .A2(_23470_),
    .B1(_21020_),
    .C1(_21023_),
    .X(_23471_));
 sky130_fd_sc_hd__a211oi_1 _26792_ (.A1(_21020_),
    .A2(_21023_),
    .B1(net272),
    .C1(_23470_),
    .Y(_23472_));
 sky130_fd_sc_hd__o21bai_1 _26793_ (.A1(_21026_),
    .A2(_21027_),
    .B1_N(_21025_),
    .Y(_23473_));
 sky130_fd_sc_hd__or3b_1 _26794_ (.A(_23471_),
    .B(_23472_),
    .C_N(_23473_),
    .X(_23474_));
 sky130_fd_sc_hd__o21bai_1 _26795_ (.A1(_23471_),
    .A2(_23472_),
    .B1_N(_23473_),
    .Y(_23475_));
 sky130_fd_sc_hd__and2_1 _26796_ (.A(_23474_),
    .B(_23475_),
    .X(_23476_));
 sky130_fd_sc_hd__o22ai_2 _26797_ (.A1(_23439_),
    .A2(_23440_),
    .B1(_23461_),
    .B2(_23462_),
    .Y(_23477_));
 sky130_fd_sc_hd__and3_1 _26798_ (.A(_23463_),
    .B(_23476_),
    .C(_23477_),
    .X(_23478_));
 sky130_fd_sc_hd__a21oi_1 _26799_ (.A1(_23477_),
    .A2(_23463_),
    .B1(_23476_),
    .Y(_23479_));
 sky130_fd_sc_hd__nor2_4 _26800_ (.A(_23478_),
    .B(_23479_),
    .Y(_23481_));
 sky130_fd_sc_hd__or2_1 _26801_ (.A(_21056_),
    .B(_21075_),
    .X(_23482_));
 sky130_fd_sc_hd__nand4b_2 _26802_ (.A_N(net298),
    .B(_19715_),
    .C(_21049_),
    .D(_20827_),
    .Y(_23483_));
 sky130_fd_sc_hd__and2b_1 _26803_ (.A_N(\delay_line[36][4] ),
    .B(\delay_line[36][6] ),
    .X(_23484_));
 sky130_fd_sc_hd__and2b_1 _26804_ (.A_N(\delay_line[36][6] ),
    .B(_21046_),
    .X(_23485_));
 sky130_fd_sc_hd__nor2_1 _26805_ (.A(_23484_),
    .B(_23485_),
    .Y(_23486_));
 sky130_fd_sc_hd__a211oi_2 _26806_ (.A1(_20825_),
    .A2(_21051_),
    .B1(_23486_),
    .C1(_21048_),
    .Y(_23487_));
 sky130_fd_sc_hd__and3b_1 _26807_ (.A_N(_18545_),
    .B(_21046_),
    .C(_21051_),
    .X(_23488_));
 sky130_fd_sc_hd__o21a_1 _26808_ (.A1(_21048_),
    .A2(_23488_),
    .B1(_23486_),
    .X(_23489_));
 sky130_fd_sc_hd__a211oi_4 _26809_ (.A1(_21054_),
    .A2(_23483_),
    .B1(_23487_),
    .C1(_23489_),
    .Y(_23490_));
 sky130_fd_sc_hd__o211a_1 _26810_ (.A1(_23489_),
    .A2(_23487_),
    .B1(_23483_),
    .C1(_21054_),
    .X(_23492_));
 sky130_fd_sc_hd__o21ba_1 _26811_ (.A1(_04338_),
    .A2(_21068_),
    .B1_N(_21066_),
    .X(_23493_));
 sky130_fd_sc_hd__and3b_1 _26812_ (.A_N(_21057_),
    .B(_21058_),
    .C(_20837_),
    .X(_23494_));
 sky130_fd_sc_hd__buf_1 _26813_ (.A(\delay_line[35][8] ),
    .X(_23495_));
 sky130_fd_sc_hd__buf_1 _26814_ (.A(\delay_line[35][9] ),
    .X(_23496_));
 sky130_fd_sc_hd__nor2_1 _26815_ (.A(_23495_),
    .B(_23496_),
    .Y(_23497_));
 sky130_fd_sc_hd__and2_1 _26816_ (.A(_23495_),
    .B(\delay_line[35][9] ),
    .X(_23498_));
 sky130_fd_sc_hd__or3b_1 _26817_ (.A(_23497_),
    .B(_23498_),
    .C_N(_20838_),
    .X(_23499_));
 sky130_fd_sc_hd__o21bai_1 _26818_ (.A1(_23497_),
    .A2(_23498_),
    .B1_N(_20838_),
    .Y(_23500_));
 sky130_fd_sc_hd__o211a_1 _26819_ (.A1(_21060_),
    .A2(_23494_),
    .B1(_23499_),
    .C1(_23500_),
    .X(_23501_));
 sky130_fd_sc_hd__clkbuf_2 _26820_ (.A(_23495_),
    .X(_23503_));
 sky130_fd_sc_hd__a221oi_2 _26821_ (.A1(_20842_),
    .A2(_23503_),
    .B1(_23499_),
    .B2(_23500_),
    .C1(_23494_),
    .Y(_23504_));
 sky130_fd_sc_hd__nor3_1 _26822_ (.A(_21065_),
    .B(_23501_),
    .C(_23504_),
    .Y(_23505_));
 sky130_fd_sc_hd__o21ai_1 _26823_ (.A1(_23501_),
    .A2(_23504_),
    .B1(_21065_),
    .Y(_23506_));
 sky130_fd_sc_hd__or2b_1 _26824_ (.A(_23505_),
    .B_N(_23506_),
    .X(_23507_));
 sky130_fd_sc_hd__xor2_1 _26825_ (.A(_05909_),
    .B(_23507_),
    .X(_23508_));
 sky130_fd_sc_hd__and2b_1 _26826_ (.A_N(_23493_),
    .B(_23508_),
    .X(_23509_));
 sky130_fd_sc_hd__and2b_1 _26827_ (.A_N(_23508_),
    .B(_23493_),
    .X(_23510_));
 sky130_fd_sc_hd__nor2_1 _26828_ (.A(_23509_),
    .B(_23510_),
    .Y(_23511_));
 sky130_fd_sc_hd__a21o_1 _26829_ (.A1(_21074_),
    .A2(_21073_),
    .B1(_21071_),
    .X(_23512_));
 sky130_fd_sc_hd__nor2_1 _26830_ (.A(_23511_),
    .B(_23512_),
    .Y(_23514_));
 sky130_fd_sc_hd__and2_1 _26831_ (.A(_23512_),
    .B(_23511_),
    .X(_23515_));
 sky130_fd_sc_hd__nor4_1 _26832_ (.A(_23490_),
    .B(_23492_),
    .C(_23514_),
    .D(_23515_),
    .Y(_23516_));
 sky130_fd_sc_hd__inv_2 _26833_ (.A(_23516_),
    .Y(_23517_));
 sky130_fd_sc_hd__o22ai_4 _26834_ (.A1(_23490_),
    .A2(_23492_),
    .B1(_23514_),
    .B2(_23515_),
    .Y(_23518_));
 sky130_fd_sc_hd__nand2_1 _26835_ (.A(_21036_),
    .B(_21038_),
    .Y(_23519_));
 sky130_fd_sc_hd__and2b_1 _26836_ (.A_N(net292),
    .B(\delay_line[37][9] ),
    .X(_23520_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26837_ (.A(\delay_line[37][9] ),
    .X(_23521_));
 sky130_fd_sc_hd__and2b_1 _26838_ (.A_N(_23521_),
    .B(net292),
    .X(_23522_));
 sky130_fd_sc_hd__nor2_1 _26839_ (.A(_23520_),
    .B(_23522_),
    .Y(_23523_));
 sky130_fd_sc_hd__a21bo_1 _26840_ (.A1(_20817_),
    .A2(_21037_),
    .B1_N(_21035_),
    .X(_23525_));
 sky130_fd_sc_hd__xnor2_1 _26841_ (.A(_23523_),
    .B(_23525_),
    .Y(_23526_));
 sky130_fd_sc_hd__a21oi_1 _26842_ (.A1(_21044_),
    .A2(_23519_),
    .B1(_23526_),
    .Y(_23527_));
 sky130_fd_sc_hd__and3_1 _26843_ (.A(_21044_),
    .B(_23526_),
    .C(_23519_),
    .X(_23528_));
 sky130_fd_sc_hd__nor2_2 _26844_ (.A(_23527_),
    .B(_23528_),
    .Y(_23529_));
 sky130_fd_sc_hd__and3_2 _26845_ (.A(_23517_),
    .B(_23518_),
    .C(_23529_),
    .X(_23530_));
 sky130_fd_sc_hd__a21oi_2 _26846_ (.A1(_23517_),
    .A2(_23518_),
    .B1(_23529_),
    .Y(_23531_));
 sky130_fd_sc_hd__a211oi_4 _26847_ (.A1(_23482_),
    .A2(_21077_),
    .B1(_23530_),
    .C1(_23531_),
    .Y(_23532_));
 sky130_fd_sc_hd__o221ai_4 _26848_ (.A1(_21056_),
    .A2(_21075_),
    .B1(_23530_),
    .B2(_23531_),
    .C1(_21077_),
    .Y(_23533_));
 sky130_fd_sc_hd__and2b_1 _26849_ (.A_N(_23532_),
    .B(_23533_),
    .X(_23534_));
 sky130_fd_sc_hd__xnor2_2 _26850_ (.A(_23481_),
    .B(_23534_),
    .Y(_23536_));
 sky130_fd_sc_hd__nand2_1 _26851_ (.A(_23428_),
    .B(_23536_),
    .Y(_23537_));
 sky130_fd_sc_hd__or2_1 _26852_ (.A(_23428_),
    .B(_23536_),
    .X(_23538_));
 sky130_fd_sc_hd__and3_2 _26853_ (.A(_23307_),
    .B(_23537_),
    .C(_23538_),
    .X(_23539_));
 sky130_fd_sc_hd__a21oi_1 _26854_ (.A1(_23537_),
    .A2(_23538_),
    .B1(_23307_),
    .Y(_23540_));
 sky130_fd_sc_hd__or2_1 _26855_ (.A(_23539_),
    .B(_23540_),
    .X(_23541_));
 sky130_fd_sc_hd__a21o_1 _26856_ (.A1(_21192_),
    .A2(_21193_),
    .B1(_23541_),
    .X(_23542_));
 sky130_fd_sc_hd__o211ai_1 _26857_ (.A1(_21083_),
    .A2(_21194_),
    .B1(_23541_),
    .C1(_21192_),
    .Y(_23543_));
 sky130_fd_sc_hd__nand2_1 _26858_ (.A(_23542_),
    .B(_23543_),
    .Y(_23544_));
 sky130_fd_sc_hd__xnor2_1 _26859_ (.A(_23306_),
    .B(_23544_),
    .Y(_23545_));
 sky130_fd_sc_hd__a21oi_2 _26860_ (.A1(_21665_),
    .A2(_21670_),
    .B1(_23545_),
    .Y(_23547_));
 sky130_fd_sc_hd__o211a_1 _26861_ (.A1(_21666_),
    .A2(_21664_),
    .B1(_21670_),
    .C1(_23545_),
    .X(_23548_));
 sky130_fd_sc_hd__nor2_1 _26862_ (.A(_23547_),
    .B(_23548_),
    .Y(_23549_));
 sky130_fd_sc_hd__o21bai_2 _26863_ (.A1(_22805_),
    .A2(_22808_),
    .B1_N(_23549_),
    .Y(_23550_));
 sky130_fd_sc_hd__o211ai_2 _26864_ (.A1(_22126_),
    .A2(_22806_),
    .B1(_22807_),
    .C1(_22803_),
    .Y(_23551_));
 sky130_fd_sc_hd__nand3b_1 _26865_ (.A_N(_22805_),
    .B(_23551_),
    .C(_23549_),
    .Y(_23552_));
 sky130_fd_sc_hd__and3_1 _26866_ (.A(_22213_),
    .B(_23550_),
    .C(_23552_),
    .X(_23553_));
 sky130_fd_sc_hd__o21ai_1 _26867_ (.A1(_20871_),
    .A2(_22149_),
    .B1(_22141_),
    .Y(_23554_));
 sky130_fd_sc_hd__nor2_1 _26868_ (.A(_20929_),
    .B(_20931_),
    .Y(_23555_));
 sky130_fd_sc_hd__and3_1 _26869_ (.A(_19790_),
    .B(_19795_),
    .C(_23555_),
    .X(_23556_));
 sky130_fd_sc_hd__clkbuf_2 _26870_ (.A(\delay_line[20][9] ),
    .X(_23558_));
 sky130_fd_sc_hd__nor2_1 _26871_ (.A(_20930_),
    .B(_23558_),
    .Y(_23559_));
 sky130_fd_sc_hd__and2_1 _26872_ (.A(_20930_),
    .B(\delay_line[20][9] ),
    .X(_23560_));
 sky130_fd_sc_hd__nor2_1 _26873_ (.A(_23559_),
    .B(_23560_),
    .Y(_23561_));
 sky130_fd_sc_hd__and3_1 _26874_ (.A(_19792_),
    .B(_20930_),
    .C(_23561_),
    .X(_23562_));
 sky130_fd_sc_hd__buf_1 _26875_ (.A(_20930_),
    .X(_23563_));
 sky130_fd_sc_hd__o2bb2a_1 _26876_ (.A1_N(_19792_),
    .A2_N(_23563_),
    .B1(_23559_),
    .B2(_23560_),
    .X(_23564_));
 sky130_fd_sc_hd__nor2_1 _26877_ (.A(_19791_),
    .B(_19793_),
    .Y(_23565_));
 sky130_fd_sc_hd__xnor2_1 _26878_ (.A(_18740_),
    .B(_23565_),
    .Y(_23566_));
 sky130_fd_sc_hd__or3_2 _26879_ (.A(_23562_),
    .B(_23564_),
    .C(_23566_),
    .X(_23567_));
 sky130_fd_sc_hd__clkbuf_2 _26880_ (.A(_23566_),
    .X(_23569_));
 sky130_fd_sc_hd__o21ai_1 _26881_ (.A1(_23562_),
    .A2(_23564_),
    .B1(_23569_),
    .Y(_23570_));
 sky130_fd_sc_hd__o211a_1 _26882_ (.A1(_23556_),
    .A2(_20934_),
    .B1(_23567_),
    .C1(_23570_),
    .X(_23571_));
 sky130_fd_sc_hd__a221oi_1 _26883_ (.A1(_19791_),
    .A2(_23555_),
    .B1(_23567_),
    .B2(_23570_),
    .C1(_20934_),
    .Y(_23572_));
 sky130_fd_sc_hd__or4b_1 _26884_ (.A(_15394_),
    .B(_22127_),
    .C(_22128_),
    .D_N(_19216_),
    .X(_23573_));
 sky130_fd_sc_hd__o21a_1 _26885_ (.A1(_23571_),
    .A2(_23572_),
    .B1(_23573_),
    .X(_23574_));
 sky130_fd_sc_hd__or3_1 _26886_ (.A(_23573_),
    .B(_23571_),
    .C(_23572_),
    .X(_23575_));
 sky130_fd_sc_hd__or2b_1 _26887_ (.A(_23574_),
    .B_N(_23575_),
    .X(_23576_));
 sky130_fd_sc_hd__xor2_1 _26888_ (.A(_20940_),
    .B(_23576_),
    .X(_23577_));
 sky130_fd_sc_hd__o311a_1 _26889_ (.A1(_20291_),
    .A2(_20940_),
    .A3(_20937_),
    .B1(_20942_),
    .C1(_23577_),
    .X(_23578_));
 sky130_fd_sc_hd__o31a_1 _26890_ (.A1(_20291_),
    .A2(_20940_),
    .A3(_20937_),
    .B1(_20942_),
    .X(_23579_));
 sky130_fd_sc_hd__nor2_1 _26891_ (.A(_23577_),
    .B(_23579_),
    .Y(_23580_));
 sky130_fd_sc_hd__nor2_1 _26892_ (.A(_23578_),
    .B(_23580_),
    .Y(_23581_));
 sky130_fd_sc_hd__and3_1 _26893_ (.A(_20956_),
    .B(_20960_),
    .C(_20953_),
    .X(_23582_));
 sky130_fd_sc_hd__a21boi_1 _26894_ (.A1(_11449_),
    .A2(_18800_),
    .B1_N(_19796_),
    .Y(_23583_));
 sky130_fd_sc_hd__nor2_1 _26895_ (.A(_23583_),
    .B(_18798_),
    .Y(_23584_));
 sky130_fd_sc_hd__and2_1 _26896_ (.A(_18798_),
    .B(_23583_),
    .X(_23585_));
 sky130_fd_sc_hd__nor3_1 _26897_ (.A(_18814_),
    .B(_23584_),
    .C(_23585_),
    .Y(_23586_));
 sky130_fd_sc_hd__o21a_1 _26898_ (.A1(_23584_),
    .A2(_23585_),
    .B1(_18814_),
    .X(_23587_));
 sky130_fd_sc_hd__nor2_1 _26899_ (.A(_20948_),
    .B(_20950_),
    .Y(_23588_));
 sky130_fd_sc_hd__o21ai_1 _26900_ (.A1(net234),
    .A2(_23587_),
    .B1(_23588_),
    .Y(_23590_));
 sky130_fd_sc_hd__or3_1 _26901_ (.A(_23588_),
    .B(net234),
    .C(_23587_),
    .X(_23591_));
 sky130_fd_sc_hd__inv_2 _26902_ (.A(\delay_line[17][9] ),
    .Y(_23592_));
 sky130_fd_sc_hd__and2_1 _26903_ (.A(_23592_),
    .B(net377),
    .X(_23593_));
 sky130_fd_sc_hd__nor2_1 _26904_ (.A(net377),
    .B(_23592_),
    .Y(_23594_));
 sky130_fd_sc_hd__or2_2 _26905_ (.A(_23593_),
    .B(_23594_),
    .X(_23595_));
 sky130_fd_sc_hd__xnor2_1 _26906_ (.A(_11020_),
    .B(_23595_),
    .Y(_23596_));
 sky130_fd_sc_hd__and3_1 _26907_ (.A(_23590_),
    .B(_23591_),
    .C(_23596_),
    .X(_23597_));
 sky130_fd_sc_hd__a21oi_1 _26908_ (.A1(_23590_),
    .A2(_23591_),
    .B1(_23596_),
    .Y(_23598_));
 sky130_fd_sc_hd__or4_2 _26909_ (.A(_20955_),
    .B(_23582_),
    .C(_23597_),
    .D(_23598_),
    .X(_23599_));
 sky130_fd_sc_hd__o22ai_4 _26910_ (.A1(_20955_),
    .A2(_23582_),
    .B1(_23597_),
    .B2(_23598_),
    .Y(_23601_));
 sky130_fd_sc_hd__buf_1 _26911_ (.A(\delay_line[17][8] ),
    .X(_23602_));
 sky130_fd_sc_hd__or3b_1 _26912_ (.A(_22183_),
    .B(_23602_),
    .C_N(_19809_),
    .X(_23603_));
 sky130_fd_sc_hd__clkbuf_2 _26913_ (.A(_19810_),
    .X(_23604_));
 sky130_fd_sc_hd__nand3b_1 _26914_ (.A_N(_20964_),
    .B(_23602_),
    .C(_22183_),
    .Y(_23605_));
 sky130_fd_sc_hd__and3_1 _26915_ (.A(_23603_),
    .B(_23604_),
    .C(_23605_),
    .X(_23606_));
 sky130_fd_sc_hd__a21oi_2 _26916_ (.A1(_23605_),
    .A2(_23603_),
    .B1(_23604_),
    .Y(_23607_));
 sky130_fd_sc_hd__a211o_1 _26917_ (.A1(_23599_),
    .A2(_23601_),
    .B1(_23606_),
    .C1(_23607_),
    .X(_23608_));
 sky130_fd_sc_hd__o211ai_4 _26918_ (.A1(_23606_),
    .A2(_23607_),
    .B1(_23599_),
    .C1(_23601_),
    .Y(_23609_));
 sky130_fd_sc_hd__and3_1 _26919_ (.A(_23581_),
    .B(_23608_),
    .C(_23609_),
    .X(_23610_));
 sky130_fd_sc_hd__a21oi_1 _26920_ (.A1(_23608_),
    .A2(_23609_),
    .B1(_23581_),
    .Y(_23612_));
 sky130_fd_sc_hd__or2_1 _26921_ (.A(_23610_),
    .B(_23612_),
    .X(_23613_));
 sky130_fd_sc_hd__a21o_1 _26922_ (.A1(_22146_),
    .A2(_23554_),
    .B1(_23613_),
    .X(_23614_));
 sky130_fd_sc_hd__nand3_1 _26923_ (.A(_22146_),
    .B(_23554_),
    .C(_23613_),
    .Y(_23615_));
 sky130_fd_sc_hd__nand2_1 _26924_ (.A(_23614_),
    .B(_23615_),
    .Y(_23616_));
 sky130_fd_sc_hd__and2b_1 _26925_ (.A_N(_20945_),
    .B(_20974_),
    .X(_23617_));
 sky130_fd_sc_hd__a21o_1 _26926_ (.A1(_20927_),
    .A2(_20944_),
    .B1(_23617_),
    .X(_23618_));
 sky130_fd_sc_hd__and2_1 _26927_ (.A(_23616_),
    .B(_23618_),
    .X(_23619_));
 sky130_fd_sc_hd__nor2_1 _26928_ (.A(_23616_),
    .B(_23618_),
    .Y(_23620_));
 sky130_fd_sc_hd__a21o_1 _26929_ (.A1(_23550_),
    .A2(_23552_),
    .B1(_22213_),
    .X(_23621_));
 sky130_fd_sc_hd__o21ai_1 _26930_ (.A1(_23619_),
    .A2(_23620_),
    .B1(_23621_),
    .Y(_23623_));
 sky130_fd_sc_hd__a21oi_1 _26931_ (.A1(_23550_),
    .A2(_23552_),
    .B1(_22213_),
    .Y(_23624_));
 sky130_fd_sc_hd__nor2_1 _26932_ (.A(_23619_),
    .B(_23620_),
    .Y(_23625_));
 sky130_fd_sc_hd__o21ai_1 _26933_ (.A1(_23624_),
    .A2(_23553_),
    .B1(_23625_),
    .Y(_23626_));
 sky130_fd_sc_hd__o221ai_2 _26934_ (.A1(_22160_),
    .A2(_22212_),
    .B1(_23553_),
    .B2(_23623_),
    .C1(_23626_),
    .Y(_23627_));
 sky130_fd_sc_hd__buf_1 _26935_ (.A(_23627_),
    .X(_23628_));
 sky130_fd_sc_hd__o21bai_1 _26936_ (.A1(_23624_),
    .A2(_23553_),
    .B1_N(_23625_),
    .Y(_23629_));
 sky130_fd_sc_hd__o31a_1 _26937_ (.A1(_20980_),
    .A2(_20981_),
    .A3(_22158_),
    .B1(_22167_),
    .X(_23630_));
 sky130_fd_sc_hd__nand2_1 _26938_ (.A(_23551_),
    .B(_23549_),
    .Y(_23631_));
 sky130_fd_sc_hd__o211ai_1 _26939_ (.A1(_23631_),
    .A2(_22805_),
    .B1(_22213_),
    .C1(_23550_),
    .Y(_23632_));
 sky130_fd_sc_hd__nand3_1 _26940_ (.A(_23621_),
    .B(_23632_),
    .C(_23625_),
    .Y(_23634_));
 sky130_fd_sc_hd__nand3_2 _26941_ (.A(_23629_),
    .B(_23630_),
    .C(_23634_),
    .Y(_23635_));
 sky130_fd_sc_hd__a21boi_2 _26942_ (.A1(_20977_),
    .A2(_20979_),
    .B1_N(_20976_),
    .Y(_23636_));
 sky130_fd_sc_hd__and3_1 _26943_ (.A(_20898_),
    .B(_18780_),
    .C(_18823_),
    .X(_23637_));
 sky130_fd_sc_hd__nor2_1 _26944_ (.A(_05161_),
    .B(_22177_),
    .Y(_23638_));
 sky130_fd_sc_hd__nor2_1 _26945_ (.A(_22139_),
    .B(_19757_),
    .Y(_23639_));
 sky130_fd_sc_hd__nor4_1 _26946_ (.A(_20965_),
    .B(_20966_),
    .C(_23638_),
    .D(_23639_),
    .Y(_23640_));
 sky130_fd_sc_hd__o22a_1 _26947_ (.A1(_20965_),
    .A2(_20966_),
    .B1(_23638_),
    .B2(_23639_),
    .X(_23641_));
 sky130_fd_sc_hd__o211ai_1 _26948_ (.A1(_23640_),
    .A2(_23641_),
    .B1(_20971_),
    .C1(_20972_),
    .Y(_23642_));
 sky130_fd_sc_hd__a211o_2 _26949_ (.A1(_20971_),
    .A2(_20972_),
    .B1(_23640_),
    .C1(_23641_),
    .X(_23643_));
 sky130_fd_sc_hd__or4bb_4 _26950_ (.A(_18824_),
    .B(_19826_),
    .C_N(_23642_),
    .D_N(_23643_),
    .X(_23645_));
 sky130_fd_sc_hd__a32o_1 _26951_ (.A1(_22177_),
    .A2(_18780_),
    .A3(_22178_),
    .B1(_23642_),
    .B2(_23643_),
    .X(_23646_));
 sky130_fd_sc_hd__o211a_2 _26952_ (.A1(_23637_),
    .A2(_22182_),
    .B1(_23645_),
    .C1(_23646_),
    .X(_23647_));
 sky130_fd_sc_hd__a211oi_1 _26953_ (.A1(_23645_),
    .A2(_23646_),
    .B1(_23637_),
    .C1(_22182_),
    .Y(_23648_));
 sky130_fd_sc_hd__nor2_1 _26954_ (.A(_23647_),
    .B(_23648_),
    .Y(_23649_));
 sky130_fd_sc_hd__xor2_2 _26955_ (.A(_23636_),
    .B(_23649_),
    .X(_23650_));
 sky130_fd_sc_hd__xor2_2 _26956_ (.A(_22187_),
    .B(_23650_),
    .X(_23651_));
 sky130_fd_sc_hd__a21oi_1 _26957_ (.A1(_23628_),
    .A2(_23635_),
    .B1(_23651_),
    .Y(_23652_));
 sky130_fd_sc_hd__and3_1 _26958_ (.A(_23627_),
    .B(_23635_),
    .C(_23651_),
    .X(_23653_));
 sky130_fd_sc_hd__a31oi_1 _26959_ (.A1(_22173_),
    .A2(_22170_),
    .A3(_22171_),
    .B1(_22195_),
    .Y(_23654_));
 sky130_fd_sc_hd__a31o_1 _26960_ (.A1(_20925_),
    .A2(_22162_),
    .A3(_22168_),
    .B1(_23654_),
    .X(_23656_));
 sky130_fd_sc_hd__o21bai_4 _26961_ (.A1(_23652_),
    .A2(_23653_),
    .B1_N(_23656_),
    .Y(_23657_));
 sky130_fd_sc_hd__a21o_1 _26962_ (.A1(_23628_),
    .A2(_23635_),
    .B1(_23651_),
    .X(_23658_));
 sky130_fd_sc_hd__nand3_1 _26963_ (.A(_23628_),
    .B(_23635_),
    .C(_23651_),
    .Y(_23659_));
 sky130_fd_sc_hd__nand3_2 _26964_ (.A(_23656_),
    .B(_23658_),
    .C(_23659_),
    .Y(_23660_));
 sky130_fd_sc_hd__nand2_1 _26965_ (.A(_22189_),
    .B(_22190_),
    .Y(_23661_));
 sky130_fd_sc_hd__a21boi_1 _26966_ (.A1(_19839_),
    .A2(_22176_),
    .B1_N(_22188_),
    .Y(_23662_));
 sky130_fd_sc_hd__a31o_2 _26967_ (.A1(_23661_),
    .A2(_22192_),
    .A3(_20895_),
    .B1(_23662_),
    .X(_23663_));
 sky130_fd_sc_hd__a21oi_2 _26968_ (.A1(_23657_),
    .A2(_23660_),
    .B1(_23663_),
    .Y(_23664_));
 sky130_fd_sc_hd__a21boi_1 _26969_ (.A1(_22199_),
    .A2(_22203_),
    .B1_N(_22200_),
    .Y(_23665_));
 sky130_fd_sc_hd__a31o_1 _26970_ (.A1(_23663_),
    .A2(_23657_),
    .A3(_23660_),
    .B1(_23665_),
    .X(_23667_));
 sky130_fd_sc_hd__a21o_1 _26971_ (.A1(_23657_),
    .A2(_23660_),
    .B1(_23663_),
    .X(_23668_));
 sky130_fd_sc_hd__nand3_1 _26972_ (.A(_23663_),
    .B(_23657_),
    .C(_23660_),
    .Y(_23669_));
 sky130_fd_sc_hd__a21boi_2 _26973_ (.A1(_23668_),
    .A2(_23669_),
    .B1_N(_23665_),
    .Y(_23670_));
 sky130_fd_sc_hd__o21ba_1 _26974_ (.A1(_23664_),
    .A2(_23667_),
    .B1_N(_23670_),
    .X(_23671_));
 sky130_fd_sc_hd__xnor2_2 _26975_ (.A(_22211_),
    .B(_23671_),
    .Y(_00040_));
 sky130_fd_sc_hd__o22ai_4 _26976_ (.A1(_23664_),
    .A2(_23667_),
    .B1(_23670_),
    .B2(_22211_),
    .Y(_23672_));
 sky130_fd_sc_hd__nand2_1 _26977_ (.A(_23635_),
    .B(_23651_),
    .Y(_23673_));
 sky130_fd_sc_hd__nand2_1 _26978_ (.A(_23628_),
    .B(_23673_),
    .Y(_23674_));
 sky130_fd_sc_hd__o21ai_1 _26979_ (.A1(_23625_),
    .A2(_23624_),
    .B1(_23632_),
    .Y(_23675_));
 sky130_fd_sc_hd__a31o_1 _26980_ (.A1(_23581_),
    .A2(_23608_),
    .A3(_23609_),
    .B1(_23580_),
    .X(_23677_));
 sky130_fd_sc_hd__or4_1 _26981_ (.A(_20934_),
    .B(_20935_),
    .C(_20936_),
    .D(_23576_),
    .X(_23678_));
 sky130_fd_sc_hd__a21boi_1 _26982_ (.A1(_23513_),
    .A2(_22783_),
    .B1_N(_22780_),
    .Y(_23679_));
 sky130_fd_sc_hd__or3b_1 _26983_ (.A(_23559_),
    .B(_23560_),
    .C_N(_20929_),
    .X(_23680_));
 sky130_fd_sc_hd__buf_1 _26984_ (.A(_23558_),
    .X(_23681_));
 sky130_fd_sc_hd__clkbuf_2 _26985_ (.A(\delay_line[20][10] ),
    .X(_23682_));
 sky130_fd_sc_hd__nor2_1 _26986_ (.A(_23558_),
    .B(_23682_),
    .Y(_23683_));
 sky130_fd_sc_hd__and2_1 _26987_ (.A(_23558_),
    .B(\delay_line[20][10] ),
    .X(_23684_));
 sky130_fd_sc_hd__nor2_1 _26988_ (.A(_23683_),
    .B(_23684_),
    .Y(_23685_));
 sky130_fd_sc_hd__and3_1 _26989_ (.A(_23563_),
    .B(_23681_),
    .C(_23685_),
    .X(_23686_));
 sky130_fd_sc_hd__o2bb2a_1 _26990_ (.A1_N(_23563_),
    .A2_N(_23681_),
    .B1(_23683_),
    .B2(_23684_),
    .X(_23688_));
 sky130_fd_sc_hd__xnor2_1 _26991_ (.A(_19790_),
    .B(_23555_),
    .Y(_23689_));
 sky130_fd_sc_hd__or3_1 _26992_ (.A(_23686_),
    .B(_23688_),
    .C(_23689_),
    .X(_23690_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26993_ (.A(_23689_),
    .X(_23691_));
 sky130_fd_sc_hd__o21ai_1 _26994_ (.A1(_23686_),
    .A2(_23688_),
    .B1(_23691_),
    .Y(_23692_));
 sky130_fd_sc_hd__nand2_1 _26995_ (.A(_23690_),
    .B(_23692_),
    .Y(_23693_));
 sky130_fd_sc_hd__a21oi_2 _26996_ (.A1(_23680_),
    .A2(_23567_),
    .B1(_23693_),
    .Y(_23694_));
 sky130_fd_sc_hd__and3_1 _26997_ (.A(_23680_),
    .B(_23567_),
    .C(_23693_),
    .X(_23695_));
 sky130_fd_sc_hd__or3_1 _26998_ (.A(_23679_),
    .B(_23694_),
    .C(_23695_),
    .X(_23696_));
 sky130_fd_sc_hd__o21ai_1 _26999_ (.A1(_23694_),
    .A2(_23695_),
    .B1(_23679_),
    .Y(_23697_));
 sky130_fd_sc_hd__and3_1 _27000_ (.A(_23696_),
    .B(_23697_),
    .C(_23571_),
    .X(_23699_));
 sky130_fd_sc_hd__a21oi_1 _27001_ (.A1(_23696_),
    .A2(_23697_),
    .B1(_23571_),
    .Y(_23700_));
 sky130_fd_sc_hd__a211oi_1 _27002_ (.A1(_23575_),
    .A2(_23678_),
    .B1(_23699_),
    .C1(_23700_),
    .Y(_23701_));
 sky130_fd_sc_hd__o221a_1 _27003_ (.A1(_23574_),
    .A2(_20938_),
    .B1(_23700_),
    .B2(_23699_),
    .C1(_23575_),
    .X(_23702_));
 sky130_fd_sc_hd__nor2_1 _27004_ (.A(_23701_),
    .B(_23702_),
    .Y(_23703_));
 sky130_fd_sc_hd__mux2_1 _27005_ (.A0(_23593_),
    .A1(_23594_),
    .S(_20946_),
    .X(_23704_));
 sky130_fd_sc_hd__xor2_2 _27006_ (.A(_20958_),
    .B(_23704_),
    .X(_23705_));
 sky130_fd_sc_hd__inv_2 _27007_ (.A(_23590_),
    .Y(_23706_));
 sky130_fd_sc_hd__a21oi_1 _27008_ (.A1(_18740_),
    .A2(_23565_),
    .B1(_19791_),
    .Y(_23707_));
 sky130_fd_sc_hd__nor2_1 _27009_ (.A(_23707_),
    .B(_19799_),
    .Y(_23708_));
 sky130_fd_sc_hd__and2_1 _27010_ (.A(_19799_),
    .B(_23707_),
    .X(_23710_));
 sky130_fd_sc_hd__nor3_1 _27011_ (.A(_19814_),
    .B(_23708_),
    .C(_23710_),
    .Y(_23711_));
 sky130_fd_sc_hd__o21a_1 _27012_ (.A1(_23708_),
    .A2(_23710_),
    .B1(_19814_),
    .X(_23712_));
 sky130_fd_sc_hd__nor2_1 _27013_ (.A(_23711_),
    .B(_23712_),
    .Y(_23713_));
 sky130_fd_sc_hd__or2_1 _27014_ (.A(_23584_),
    .B(_23586_),
    .X(_23714_));
 sky130_fd_sc_hd__nor2_1 _27015_ (.A(_23713_),
    .B(_23714_),
    .Y(_23715_));
 sky130_fd_sc_hd__o21a_1 _27016_ (.A1(_23584_),
    .A2(_23586_),
    .B1(_23713_),
    .X(_23716_));
 sky130_fd_sc_hd__or2_1 _27017_ (.A(_23715_),
    .B(_23716_),
    .X(_23717_));
 sky130_fd_sc_hd__nor2_1 _27018_ (.A(net376),
    .B(\delay_line[17][10] ),
    .Y(_23718_));
 sky130_fd_sc_hd__buf_1 _27019_ (.A(\delay_line[17][10] ),
    .X(_23719_));
 sky130_fd_sc_hd__nand2_1 _27020_ (.A(net376),
    .B(_23719_),
    .Y(_23721_));
 sky130_fd_sc_hd__mux2_1 _27021_ (.A0(_18729_),
    .A1(_10767_),
    .S(_19819_),
    .X(_23722_));
 sky130_fd_sc_hd__and3b_1 _27022_ (.A_N(_23718_),
    .B(_23721_),
    .C(_23722_),
    .X(_23723_));
 sky130_fd_sc_hd__and2_1 _27023_ (.A(net376),
    .B(\delay_line[17][10] ),
    .X(_23724_));
 sky130_fd_sc_hd__nor2_1 _27024_ (.A(_23718_),
    .B(_23724_),
    .Y(_23725_));
 sky130_fd_sc_hd__nor2_1 _27025_ (.A(_23725_),
    .B(_23722_),
    .Y(_23726_));
 sky130_fd_sc_hd__nor2_1 _27026_ (.A(_23723_),
    .B(_23726_),
    .Y(_23727_));
 sky130_fd_sc_hd__and2_1 _27027_ (.A(_23717_),
    .B(_23727_),
    .X(_23728_));
 sky130_fd_sc_hd__nor2_2 _27028_ (.A(_23727_),
    .B(_23717_),
    .Y(_23729_));
 sky130_fd_sc_hd__or2_1 _27029_ (.A(_23728_),
    .B(_23729_),
    .X(_23730_));
 sky130_fd_sc_hd__o211a_1 _27030_ (.A1(_23596_),
    .A2(_23706_),
    .B1(_23591_),
    .C1(_23730_),
    .X(_23732_));
 sky130_fd_sc_hd__o32a_1 _27031_ (.A1(_23588_),
    .A2(net234),
    .A3(_23587_),
    .B1(_23596_),
    .B2(_23706_),
    .X(_23733_));
 sky130_fd_sc_hd__or2_1 _27032_ (.A(_23733_),
    .B(_23730_),
    .X(_23734_));
 sky130_fd_sc_hd__and2b_1 _27033_ (.A_N(_23732_),
    .B(_23734_),
    .X(_23735_));
 sky130_fd_sc_hd__xor2_2 _27034_ (.A(_23705_),
    .B(_23735_),
    .X(_23736_));
 sky130_fd_sc_hd__xor2_1 _27035_ (.A(_23703_),
    .B(_23736_),
    .X(_23737_));
 sky130_fd_sc_hd__a31o_1 _27036_ (.A1(_22801_),
    .A2(_22794_),
    .A3(_22802_),
    .B1(_22804_),
    .X(_23738_));
 sky130_fd_sc_hd__and3_1 _27037_ (.A(_22807_),
    .B(_23737_),
    .C(_23738_),
    .X(_23739_));
 sky130_fd_sc_hd__a21oi_1 _27038_ (.A1(_22807_),
    .A2(_23738_),
    .B1(_23737_),
    .Y(_23740_));
 sky130_fd_sc_hd__nor2_1 _27039_ (.A(_23739_),
    .B(_23740_),
    .Y(_23741_));
 sky130_fd_sc_hd__nor2_1 _27040_ (.A(_23677_),
    .B(_23741_),
    .Y(_23743_));
 sky130_fd_sc_hd__and2_1 _27041_ (.A(_23741_),
    .B(_23677_),
    .X(_23744_));
 sky130_fd_sc_hd__nand2_1 _27042_ (.A(_22738_),
    .B(_22740_),
    .Y(_23745_));
 sky130_fd_sc_hd__nand2_1 _27043_ (.A(_22221_),
    .B(_22736_),
    .Y(_23746_));
 sky130_fd_sc_hd__nor2_1 _27044_ (.A(_22222_),
    .B(_22266_),
    .Y(_23747_));
 sky130_fd_sc_hd__a31oi_1 _27045_ (.A1(_22417_),
    .A2(_22421_),
    .A3(_22406_),
    .B1(_22416_),
    .Y(_23748_));
 sky130_fd_sc_hd__a21boi_1 _27046_ (.A1(_23748_),
    .A2(_22428_),
    .B1_N(_22495_),
    .Y(_23749_));
 sky130_fd_sc_hd__o21a_1 _27047_ (.A1(_22476_),
    .A2(_22475_),
    .B1(_22472_),
    .X(_23750_));
 sky130_fd_sc_hd__a211o_1 _27048_ (.A1(_13042_),
    .A2(_08701_),
    .B1(_19957_),
    .C1(_19961_),
    .X(_23751_));
 sky130_fd_sc_hd__nand2_1 _27049_ (.A(_08712_),
    .B(_19961_),
    .Y(_23752_));
 sky130_fd_sc_hd__nand3b_1 _27050_ (.A_N(_22434_),
    .B(_23751_),
    .C(_23752_),
    .Y(_23754_));
 sky130_fd_sc_hd__buf_2 _27051_ (.A(_22436_),
    .X(_23755_));
 sky130_fd_sc_hd__a2bb2o_1 _27052_ (.A1_N(_23755_),
    .A2_N(_25051_),
    .B1(_23752_),
    .B2(_23751_),
    .X(_23756_));
 sky130_fd_sc_hd__nand2_1 _27053_ (.A(_23754_),
    .B(_23756_),
    .Y(_23757_));
 sky130_fd_sc_hd__inv_2 _27054_ (.A(\delay_line[10][10] ),
    .Y(_23758_));
 sky130_fd_sc_hd__nor2_1 _27055_ (.A(_17918_),
    .B(net412),
    .Y(_23759_));
 sky130_fd_sc_hd__and2_1 _27056_ (.A(\delay_line[10][5] ),
    .B(net412),
    .X(_23760_));
 sky130_fd_sc_hd__or3_1 _27057_ (.A(_23758_),
    .B(_23759_),
    .C(_23760_),
    .X(_23761_));
 sky130_fd_sc_hd__clkbuf_2 _27058_ (.A(_23758_),
    .X(_23762_));
 sky130_fd_sc_hd__o21ai_1 _27059_ (.A1(_23759_),
    .A2(_23760_),
    .B1(_23762_),
    .Y(_23763_));
 sky130_fd_sc_hd__nand3b_1 _27060_ (.A_N(_22450_),
    .B(_23761_),
    .C(_23763_),
    .Y(_23765_));
 sky130_fd_sc_hd__a32o_1 _27061_ (.A1(_22448_),
    .A2(_22444_),
    .A3(_22445_),
    .B1(_23761_),
    .B2(_23763_),
    .X(_23766_));
 sky130_fd_sc_hd__nand2_1 _27062_ (.A(_23765_),
    .B(_23766_),
    .Y(_23767_));
 sky130_fd_sc_hd__xnor2_2 _27063_ (.A(_23757_),
    .B(_23767_),
    .Y(_23768_));
 sky130_fd_sc_hd__and2b_2 _27064_ (.A_N(_17993_),
    .B(_17994_),
    .X(_23769_));
 sky130_fd_sc_hd__nand2_1 _27065_ (.A(_23769_),
    .B(_22460_),
    .Y(_23770_));
 sky130_fd_sc_hd__buf_2 _27066_ (.A(\delay_line[10][9] ),
    .X(_23771_));
 sky130_fd_sc_hd__a21o_1 _27067_ (.A1(_12152_),
    .A2(_23771_),
    .B1(_23769_),
    .X(_23772_));
 sky130_fd_sc_hd__and3b_1 _27068_ (.A_N(net403),
    .B(_21679_),
    .C(_20060_),
    .X(_23773_));
 sky130_fd_sc_hd__a211oi_1 _27069_ (.A1(_23770_),
    .A2(_23772_),
    .B1(_23773_),
    .C1(_22397_),
    .Y(_23774_));
 sky130_fd_sc_hd__o211a_1 _27070_ (.A1(_23773_),
    .A2(_22396_),
    .B1(_23770_),
    .C1(_23772_),
    .X(_23776_));
 sky130_fd_sc_hd__nor3_2 _27071_ (.A(_22461_),
    .B(_23774_),
    .C(_23776_),
    .Y(_23777_));
 sky130_fd_sc_hd__o21a_1 _27072_ (.A1(_23774_),
    .A2(_23776_),
    .B1(_22461_),
    .X(_23778_));
 sky130_fd_sc_hd__o211ai_1 _27073_ (.A1(_23777_),
    .A2(_23778_),
    .B1(_22464_),
    .C1(_22471_),
    .Y(_23779_));
 sky130_fd_sc_hd__a211o_1 _27074_ (.A1(_22464_),
    .A2(_22470_),
    .B1(_23777_),
    .C1(_23778_),
    .X(_23780_));
 sky130_fd_sc_hd__nand2_1 _27075_ (.A(_23779_),
    .B(_23780_),
    .Y(_23781_));
 sky130_fd_sc_hd__xor2_1 _27076_ (.A(_23768_),
    .B(_23781_),
    .X(_23782_));
 sky130_fd_sc_hd__o21ai_2 _27077_ (.A1(_21686_),
    .A2(_22403_),
    .B1(_22400_),
    .Y(_23783_));
 sky130_fd_sc_hd__xnor2_1 _27078_ (.A(_23782_),
    .B(_23783_),
    .Y(_23784_));
 sky130_fd_sc_hd__or2_1 _27079_ (.A(_23750_),
    .B(_23784_),
    .X(_23785_));
 sky130_fd_sc_hd__inv_2 _27080_ (.A(_23785_),
    .Y(_23787_));
 sky130_fd_sc_hd__o211a_1 _27081_ (.A1(_22475_),
    .A2(_22476_),
    .B1(_22472_),
    .C1(_23784_),
    .X(_23788_));
 sky130_fd_sc_hd__or2_1 _27082_ (.A(_23787_),
    .B(_23788_),
    .X(_23789_));
 sky130_fd_sc_hd__inv_2 _27083_ (.A(_23789_),
    .Y(_23790_));
 sky130_fd_sc_hd__a21oi_1 _27084_ (.A1(_22421_),
    .A2(_22407_),
    .B1(_22414_),
    .Y(_23791_));
 sky130_fd_sc_hd__nor2_1 _27085_ (.A(_22394_),
    .B(_22397_),
    .Y(_23792_));
 sky130_fd_sc_hd__nor2_1 _27086_ (.A(_12746_),
    .B(_18915_),
    .Y(_23793_));
 sky130_fd_sc_hd__and2_1 _27087_ (.A(_02480_),
    .B(_18915_),
    .X(_23794_));
 sky130_fd_sc_hd__clkbuf_4 _27088_ (.A(\delay_line[12][10] ),
    .X(_23795_));
 sky130_fd_sc_hd__nor2_1 _27089_ (.A(_23795_),
    .B(_22393_),
    .Y(_23796_));
 sky130_fd_sc_hd__clkbuf_2 _27090_ (.A(\delay_line[12][9] ),
    .X(_23798_));
 sky130_fd_sc_hd__clkbuf_2 _27091_ (.A(_23798_),
    .X(_23799_));
 sky130_fd_sc_hd__buf_1 _27092_ (.A(\delay_line[12][10] ),
    .X(_23800_));
 sky130_fd_sc_hd__and3b_1 _27093_ (.A_N(_22465_),
    .B(_23799_),
    .C(_23800_),
    .X(_23801_));
 sky130_fd_sc_hd__o22ai_1 _27094_ (.A1(_23793_),
    .A2(_23794_),
    .B1(_23796_),
    .B2(_23801_),
    .Y(_23802_));
 sky130_fd_sc_hd__or4_2 _27095_ (.A(_23793_),
    .B(_23794_),
    .C(_23796_),
    .D(_23801_),
    .X(_23803_));
 sky130_fd_sc_hd__nand2_1 _27096_ (.A(_23802_),
    .B(_23803_),
    .Y(_23804_));
 sky130_fd_sc_hd__a21o_1 _27097_ (.A1(_21697_),
    .A2(_22378_),
    .B1(_22381_),
    .X(_23805_));
 sky130_fd_sc_hd__xnor2_1 _27098_ (.A(_23804_),
    .B(_23805_),
    .Y(_23806_));
 sky130_fd_sc_hd__and3_1 _27099_ (.A(_25194_),
    .B(_23792_),
    .C(_23806_),
    .X(_23807_));
 sky130_fd_sc_hd__a21oi_1 _27100_ (.A1(_25194_),
    .A2(_23792_),
    .B1(_23806_),
    .Y(_23809_));
 sky130_fd_sc_hd__a31oi_4 _27101_ (.A1(_22373_),
    .A2(_22374_),
    .A3(_22375_),
    .B1(_22383_),
    .Y(_23810_));
 sky130_fd_sc_hd__clkbuf_2 _27102_ (.A(_20046_),
    .X(_23811_));
 sky130_fd_sc_hd__buf_2 _27103_ (.A(_23811_),
    .X(_23812_));
 sky130_fd_sc_hd__xor2_1 _27104_ (.A(_22362_),
    .B(\delay_line[13][10] ),
    .X(_23813_));
 sky130_fd_sc_hd__and4b_1 _27105_ (.A_N(\delay_line[13][10] ),
    .B(_22360_),
    .C(_17956_),
    .D(net396),
    .X(_23814_));
 sky130_fd_sc_hd__o21ba_1 _27106_ (.A1(_22361_),
    .A2(_23813_),
    .B1_N(_23814_),
    .X(_23815_));
 sky130_fd_sc_hd__a21boi_2 _27107_ (.A1(_17979_),
    .A2(_23812_),
    .B1_N(_23815_),
    .Y(_23816_));
 sky130_fd_sc_hd__and3b_1 _27108_ (.A_N(_23815_),
    .B(_23812_),
    .C(_17979_),
    .X(_23817_));
 sky130_fd_sc_hd__a21oi_2 _27109_ (.A1(_22344_),
    .A2(_22350_),
    .B1(_22353_),
    .Y(_23818_));
 sky130_fd_sc_hd__o211ai_2 _27110_ (.A1(_22274_),
    .A2(_21740_),
    .B1(_22333_),
    .C1(_22339_),
    .Y(_23820_));
 sky130_fd_sc_hd__and2_1 _27111_ (.A(_22323_),
    .B(\delay_line[0][10] ),
    .X(_23821_));
 sky130_fd_sc_hd__nor2_1 _27112_ (.A(_22323_),
    .B(\delay_line[0][10] ),
    .Y(_23822_));
 sky130_fd_sc_hd__inv_2 _27113_ (.A(_22321_),
    .Y(_23823_));
 sky130_fd_sc_hd__o21ai_1 _27114_ (.A1(_22298_),
    .A2(_22334_),
    .B1(_22302_),
    .Y(_23824_));
 sky130_fd_sc_hd__a21boi_1 _27115_ (.A1(_23823_),
    .A2(_23824_),
    .B1_N(\delay_line[0][9] ),
    .Y(_23825_));
 sky130_fd_sc_hd__o2111ai_4 _27116_ (.A1(_21702_),
    .A2(_21703_),
    .B1(_17941_),
    .C1(_19994_),
    .D1(_22277_),
    .Y(_23826_));
 sky130_fd_sc_hd__clkbuf_2 _27117_ (.A(\delay_line[4][7] ),
    .X(_23827_));
 sky130_fd_sc_hd__nand2_2 _27118_ (.A(_22287_),
    .B(_23827_),
    .Y(_23828_));
 sky130_fd_sc_hd__nand2b_4 _27119_ (.A_N(_23827_),
    .B(_22280_),
    .Y(_23829_));
 sky130_fd_sc_hd__nand2_2 _27120_ (.A(_22276_),
    .B(_21706_),
    .Y(_23831_));
 sky130_fd_sc_hd__a22oi_4 _27121_ (.A1(_23828_),
    .A2(_23829_),
    .B1(_23831_),
    .B2(_22278_),
    .Y(_23832_));
 sky130_fd_sc_hd__inv_2 _27122_ (.A(_22277_),
    .Y(_23833_));
 sky130_fd_sc_hd__o2111a_2 _27123_ (.A1(_19994_),
    .A2(_23833_),
    .B1(_23828_),
    .C1(_23829_),
    .D1(_23831_),
    .X(_23834_));
 sky130_fd_sc_hd__nor2_2 _27124_ (.A(_23832_),
    .B(_23834_),
    .Y(_23835_));
 sky130_fd_sc_hd__a21oi_1 _27125_ (.A1(_22302_),
    .A2(_23826_),
    .B1(_23835_),
    .Y(_23836_));
 sky130_fd_sc_hd__nor2b_1 _27126_ (.A(_12262_),
    .B_N(_21720_),
    .Y(_23837_));
 sky130_fd_sc_hd__o21ai_2 _27127_ (.A1(_22307_),
    .A2(_22308_),
    .B1(_23837_),
    .Y(_23838_));
 sky130_fd_sc_hd__buf_2 _27128_ (.A(\delay_line[11][8] ),
    .X(_23839_));
 sky130_fd_sc_hd__nand2b_1 _27129_ (.A_N(_23839_),
    .B(_20002_),
    .Y(_23840_));
 sky130_fd_sc_hd__nand2b_1 _27130_ (.A_N(_18933_),
    .B(\delay_line[11][8] ),
    .Y(_23842_));
 sky130_fd_sc_hd__nand2_2 _27131_ (.A(_23840_),
    .B(_23842_),
    .Y(_23843_));
 sky130_fd_sc_hd__a21oi_4 _27132_ (.A1(_22309_),
    .A2(_23838_),
    .B1(_23843_),
    .Y(_23844_));
 sky130_fd_sc_hd__o311a_2 _27133_ (.A1(_12273_),
    .A2(_21718_),
    .A3(_22305_),
    .B1(_23843_),
    .C1(_22313_),
    .X(_23845_));
 sky130_fd_sc_hd__nor2_2 _27134_ (.A(_23844_),
    .B(_23845_),
    .Y(_23846_));
 sky130_fd_sc_hd__o211a_1 _27135_ (.A1(_20012_),
    .A2(_22312_),
    .B1(_22315_),
    .C1(_23846_),
    .X(_23847_));
 sky130_fd_sc_hd__o21ai_2 _27136_ (.A1(_20011_),
    .A2(_22312_),
    .B1(_22315_),
    .Y(_23848_));
 sky130_fd_sc_hd__clkbuf_2 _27137_ (.A(_23848_),
    .X(_23849_));
 sky130_fd_sc_hd__o21a_1 _27138_ (.A1(_23844_),
    .A2(_23845_),
    .B1(_23849_),
    .X(_23850_));
 sky130_fd_sc_hd__a311o_1 _27139_ (.A1(_22277_),
    .A2(_21700_),
    .A3(_22296_),
    .B1(_23832_),
    .C1(_23834_),
    .X(_23851_));
 sky130_fd_sc_hd__o22ai_1 _27140_ (.A1(_23847_),
    .A2(_23850_),
    .B1(_23851_),
    .B2(_22331_),
    .Y(_23853_));
 sky130_fd_sc_hd__nor2_1 _27141_ (.A(_23836_),
    .B(_23853_),
    .Y(_23854_));
 sky130_fd_sc_hd__and3_1 _27142_ (.A(_22277_),
    .B(_21700_),
    .C(_22296_),
    .X(_23855_));
 sky130_fd_sc_hd__o22ai_4 _27143_ (.A1(_23832_),
    .A2(_23834_),
    .B1(_23855_),
    .B2(_22331_),
    .Y(_23856_));
 sky130_fd_sc_hd__nand3_1 _27144_ (.A(_22301_),
    .B(_23835_),
    .C(_23826_),
    .Y(_23857_));
 sky130_fd_sc_hd__nand2_1 _27145_ (.A(_23848_),
    .B(_23846_),
    .Y(_23858_));
 sky130_fd_sc_hd__o21a_1 _27146_ (.A1(_20011_),
    .A2(_22312_),
    .B1(_22315_),
    .X(_23859_));
 sky130_fd_sc_hd__o21ai_1 _27147_ (.A1(_23844_),
    .A2(_23845_),
    .B1(_23859_),
    .Y(_23860_));
 sky130_fd_sc_hd__and2_1 _27148_ (.A(_23858_),
    .B(_23860_),
    .X(_23861_));
 sky130_fd_sc_hd__a21oi_2 _27149_ (.A1(_23856_),
    .A2(_23857_),
    .B1(_23861_),
    .Y(_23862_));
 sky130_fd_sc_hd__o22ai_4 _27150_ (.A1(_22335_),
    .A2(_23825_),
    .B1(_23854_),
    .B2(_23862_),
    .Y(_23864_));
 sky130_fd_sc_hd__a22o_2 _27151_ (.A1(_23858_),
    .A2(_23860_),
    .B1(_23856_),
    .B2(_23857_),
    .X(_23865_));
 sky130_fd_sc_hd__a21oi_1 _27152_ (.A1(_22332_),
    .A2(\delay_line[0][9] ),
    .B1(_22335_),
    .Y(_23866_));
 sky130_fd_sc_hd__o221ai_2 _27153_ (.A1(_23847_),
    .A2(_23850_),
    .B1(_23851_),
    .B2(_22331_),
    .C1(_23856_),
    .Y(_23867_));
 sky130_fd_sc_hd__nand3_2 _27154_ (.A(_23865_),
    .B(_23866_),
    .C(_23867_),
    .Y(_23868_));
 sky130_fd_sc_hd__o211ai_2 _27155_ (.A1(_23821_),
    .A2(_23822_),
    .B1(_23864_),
    .C1(_23868_),
    .Y(_23869_));
 sky130_fd_sc_hd__nand2_1 _27156_ (.A(_23864_),
    .B(_23868_),
    .Y(_23870_));
 sky130_fd_sc_hd__nor2_1 _27157_ (.A(_23821_),
    .B(_23822_),
    .Y(_23871_));
 sky130_fd_sc_hd__nand2_1 _27158_ (.A(_23870_),
    .B(_23871_),
    .Y(_23872_));
 sky130_fd_sc_hd__o2111ai_4 _27159_ (.A1(_22342_),
    .A2(_22348_),
    .B1(_23820_),
    .C1(_23869_),
    .D1(_23872_),
    .Y(_23873_));
 sky130_fd_sc_hd__o22ai_2 _27160_ (.A1(_22346_),
    .A2(_22345_),
    .B1(_22348_),
    .B2(_22342_),
    .Y(_23875_));
 sky130_fd_sc_hd__o2bb2ai_1 _27161_ (.A1_N(_23864_),
    .A2_N(_23868_),
    .B1(_23821_),
    .B2(_23822_),
    .Y(_23876_));
 sky130_fd_sc_hd__nand3_1 _27162_ (.A(_23864_),
    .B(_23868_),
    .C(_23871_),
    .Y(_23877_));
 sky130_fd_sc_hd__nand3_2 _27163_ (.A(_23875_),
    .B(_23876_),
    .C(_23877_),
    .Y(_23878_));
 sky130_fd_sc_hd__clkbuf_2 _27164_ (.A(\delay_line[13][9] ),
    .X(_23879_));
 sky130_fd_sc_hd__clkbuf_2 _27165_ (.A(_18947_),
    .X(_23880_));
 sky130_fd_sc_hd__a21oi_2 _27166_ (.A1(_19982_),
    .A2(\delay_line[13][9] ),
    .B1(_19983_),
    .Y(_23881_));
 sky130_fd_sc_hd__a21oi_2 _27167_ (.A1(_23879_),
    .A2(_23880_),
    .B1(_23881_),
    .Y(_23882_));
 sky130_fd_sc_hd__nand3_2 _27168_ (.A(_23873_),
    .B(_23878_),
    .C(_23882_),
    .Y(_23883_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27169_ (.A(_23879_),
    .X(_23884_));
 sky130_fd_sc_hd__and3_2 _27170_ (.A(_19982_),
    .B(_19983_),
    .C(_23884_),
    .X(_23886_));
 sky130_fd_sc_hd__nand2_1 _27171_ (.A(_23873_),
    .B(_23878_),
    .Y(_23887_));
 sky130_fd_sc_hd__o21ai_2 _27172_ (.A1(_23886_),
    .A2(_23881_),
    .B1(_23887_),
    .Y(_23888_));
 sky130_fd_sc_hd__o211ai_4 _27173_ (.A1(_23818_),
    .A2(_22370_),
    .B1(_23883_),
    .C1(_23888_),
    .Y(_23889_));
 sky130_fd_sc_hd__nor2_1 _27174_ (.A(_22361_),
    .B(_22364_),
    .Y(_23890_));
 sky130_fd_sc_hd__a21oi_1 _27175_ (.A1(_22354_),
    .A2(_23890_),
    .B1(_23818_),
    .Y(_23891_));
 sky130_fd_sc_hd__o211ai_2 _27176_ (.A1(_23886_),
    .A2(_23881_),
    .B1(_23873_),
    .C1(_23878_),
    .Y(_23892_));
 sky130_fd_sc_hd__nand2_1 _27177_ (.A(_23887_),
    .B(_23882_),
    .Y(_23893_));
 sky130_fd_sc_hd__nand3_4 _27178_ (.A(_23891_),
    .B(_23892_),
    .C(_23893_),
    .Y(_23894_));
 sky130_fd_sc_hd__o211ai_4 _27179_ (.A1(_23816_),
    .A2(_23817_),
    .B1(_23889_),
    .C1(_23894_),
    .Y(_23895_));
 sky130_fd_sc_hd__and3_2 _27180_ (.A(_17978_),
    .B(_23811_),
    .C(_23815_),
    .X(_23897_));
 sky130_fd_sc_hd__buf_2 _27181_ (.A(_23811_),
    .X(_23898_));
 sky130_fd_sc_hd__a21oi_1 _27182_ (.A1(_17979_),
    .A2(_23898_),
    .B1(_23815_),
    .Y(_23899_));
 sky130_fd_sc_hd__o2bb2ai_2 _27183_ (.A1_N(_23889_),
    .A2_N(_23894_),
    .B1(_23897_),
    .B2(_23899_),
    .Y(_23900_));
 sky130_fd_sc_hd__o211ai_4 _27184_ (.A1(_22411_),
    .A2(_23810_),
    .B1(_23895_),
    .C1(_23900_),
    .Y(_23901_));
 sky130_fd_sc_hd__a21oi_1 _27185_ (.A1(_22376_),
    .A2(_22409_),
    .B1(_22411_),
    .Y(_23902_));
 sky130_fd_sc_hd__o211ai_1 _27186_ (.A1(_23897_),
    .A2(_23899_),
    .B1(_23889_),
    .C1(_23894_),
    .Y(_23903_));
 sky130_fd_sc_hd__o2bb2ai_1 _27187_ (.A1_N(_23889_),
    .A2_N(_23894_),
    .B1(_23816_),
    .B2(_23817_),
    .Y(_23904_));
 sky130_fd_sc_hd__nand3_1 _27188_ (.A(_23902_),
    .B(_23903_),
    .C(_23904_),
    .Y(_23905_));
 sky130_fd_sc_hd__o211ai_2 _27189_ (.A1(_23807_),
    .A2(_23809_),
    .B1(_23901_),
    .C1(_23905_),
    .Y(_23906_));
 sky130_fd_sc_hd__clkbuf_2 _27190_ (.A(_23905_),
    .X(_23908_));
 sky130_fd_sc_hd__nor2_1 _27191_ (.A(_22399_),
    .B(_23806_),
    .Y(_23909_));
 sky130_fd_sc_hd__o31a_1 _27192_ (.A1(_21678_),
    .A2(_22394_),
    .A3(_22397_),
    .B1(_23806_),
    .X(_23910_));
 sky130_fd_sc_hd__o2bb2ai_1 _27193_ (.A1_N(_23901_),
    .A2_N(_23908_),
    .B1(_23909_),
    .B2(_23910_),
    .Y(_23911_));
 sky130_fd_sc_hd__nand3_2 _27194_ (.A(_23791_),
    .B(_23906_),
    .C(_23911_),
    .Y(_23912_));
 sky130_fd_sc_hd__nand2_1 _27195_ (.A(_22417_),
    .B(_22408_),
    .Y(_23913_));
 sky130_fd_sc_hd__o2bb2ai_1 _27196_ (.A1_N(_23901_),
    .A2_N(_23905_),
    .B1(_23807_),
    .B2(_23809_),
    .Y(_23914_));
 sky130_fd_sc_hd__nor2_1 _27197_ (.A(_23807_),
    .B(_23809_),
    .Y(_23915_));
 sky130_fd_sc_hd__nand3_1 _27198_ (.A(_23901_),
    .B(_23908_),
    .C(_23915_),
    .Y(_23916_));
 sky130_fd_sc_hd__nand3_2 _27199_ (.A(_23913_),
    .B(_23914_),
    .C(_23916_),
    .Y(_23917_));
 sky130_fd_sc_hd__nand3_1 _27200_ (.A(_23790_),
    .B(_23912_),
    .C(_23917_),
    .Y(_23919_));
 sky130_fd_sc_hd__nand2_1 _27201_ (.A(_23912_),
    .B(_23917_),
    .Y(_23920_));
 sky130_fd_sc_hd__o21ai_1 _27202_ (.A1(_23787_),
    .A2(_23788_),
    .B1(_23920_),
    .Y(_23921_));
 sky130_fd_sc_hd__o211ai_2 _27203_ (.A1(_22497_),
    .A2(_23749_),
    .B1(_23919_),
    .C1(_23921_),
    .Y(_23922_));
 sky130_fd_sc_hd__a21o_1 _27204_ (.A1(_23912_),
    .A2(_23917_),
    .B1(_23789_),
    .X(_23923_));
 sky130_fd_sc_hd__a21oi_1 _27205_ (.A1(_22431_),
    .A2(_22495_),
    .B1(_22497_),
    .Y(_23924_));
 sky130_fd_sc_hd__o211ai_2 _27206_ (.A1(_23787_),
    .A2(_23788_),
    .B1(_23912_),
    .C1(_23917_),
    .Y(_23925_));
 sky130_fd_sc_hd__nand3_4 _27207_ (.A(_23923_),
    .B(_23924_),
    .C(_23925_),
    .Y(_23926_));
 sky130_fd_sc_hd__o21a_1 _27208_ (.A1(_22560_),
    .A2(_22535_),
    .B1(_22559_),
    .X(_23927_));
 sky130_fd_sc_hd__inv_2 _27209_ (.A(_23927_),
    .Y(_23928_));
 sky130_fd_sc_hd__a21oi_1 _27210_ (.A1(_22483_),
    .A2(_22433_),
    .B1(_22481_),
    .Y(_23930_));
 sky130_fd_sc_hd__nor2_1 _27211_ (.A(_03183_),
    .B(_11833_),
    .Y(_23931_));
 sky130_fd_sc_hd__and2_1 _27212_ (.A(_11822_),
    .B(_03183_),
    .X(_23932_));
 sky130_fd_sc_hd__nor3_2 _27213_ (.A(_22524_),
    .B(_23931_),
    .C(_23932_),
    .Y(_23933_));
 sky130_fd_sc_hd__o21a_1 _27214_ (.A1(_23931_),
    .A2(_23932_),
    .B1(_22524_),
    .X(_23934_));
 sky130_fd_sc_hd__o211a_1 _27215_ (.A1(_23933_),
    .A2(_23934_),
    .B1(_22513_),
    .C1(_22517_),
    .X(_23935_));
 sky130_fd_sc_hd__or2_1 _27216_ (.A(_23933_),
    .B(_23934_),
    .X(_23936_));
 sky130_fd_sc_hd__a21oi_1 _27217_ (.A1(_22513_),
    .A2(_22517_),
    .B1(_23936_),
    .Y(_23937_));
 sky130_fd_sc_hd__nor3_1 _27218_ (.A(_22528_),
    .B(_23935_),
    .C(_23937_),
    .Y(_23938_));
 sky130_fd_sc_hd__o21ai_1 _27219_ (.A1(_23935_),
    .A2(_23937_),
    .B1(_22528_),
    .Y(_23939_));
 sky130_fd_sc_hd__and2b_2 _27220_ (.A_N(_23938_),
    .B(_23939_),
    .X(_23941_));
 sky130_fd_sc_hd__nand2_1 _27221_ (.A(_22509_),
    .B(_21869_),
    .Y(_23942_));
 sky130_fd_sc_hd__clkbuf_2 _27222_ (.A(\delay_line[8][10] ),
    .X(_23943_));
 sky130_fd_sc_hd__nor3_1 _27223_ (.A(_21867_),
    .B(_22503_),
    .C(_23943_),
    .Y(_23944_));
 sky130_fd_sc_hd__nand2_1 _27224_ (.A(_22503_),
    .B(\delay_line[8][10] ),
    .Y(_23945_));
 sky130_fd_sc_hd__o21ai_1 _27225_ (.A1(\delay_line[8][9] ),
    .A2(\delay_line[8][10] ),
    .B1(net424),
    .Y(_23946_));
 sky130_fd_sc_hd__nand2_2 _27226_ (.A(_23945_),
    .B(_23946_),
    .Y(_23947_));
 sky130_fd_sc_hd__nand3_2 _27227_ (.A(_21867_),
    .B(_22503_),
    .C(_23943_),
    .Y(_23948_));
 sky130_fd_sc_hd__o21a_1 _27228_ (.A1(_23944_),
    .A2(_23947_),
    .B1(_23948_),
    .X(_23949_));
 sky130_fd_sc_hd__a21o_1 _27229_ (.A1(_23942_),
    .A2(_22514_),
    .B1(_23949_),
    .X(_23950_));
 sky130_fd_sc_hd__o2111ai_2 _27230_ (.A1(_23944_),
    .A2(_23947_),
    .B1(_23942_),
    .C1(_22514_),
    .D1(_23948_),
    .Y(_23952_));
 sky130_fd_sc_hd__clkbuf_2 _27231_ (.A(_22509_),
    .X(_23953_));
 sky130_fd_sc_hd__clkbuf_2 _27232_ (.A(_23953_),
    .X(_23954_));
 sky130_fd_sc_hd__nand3_1 _27233_ (.A(_23950_),
    .B(_23952_),
    .C(_23954_),
    .Y(_23955_));
 sky130_fd_sc_hd__a21o_1 _27234_ (.A1(_23950_),
    .A2(_23952_),
    .B1(_23953_),
    .X(_23956_));
 sky130_fd_sc_hd__nor3_1 _27235_ (.A(_22500_),
    .B(_22504_),
    .C(_21868_),
    .Y(_23957_));
 sky130_fd_sc_hd__or2_1 _27236_ (.A(_22502_),
    .B(_23957_),
    .X(_23958_));
 sky130_fd_sc_hd__xor2_1 _27237_ (.A(_18058_),
    .B(_23958_),
    .X(_23959_));
 sky130_fd_sc_hd__a21o_1 _27238_ (.A1(_23955_),
    .A2(_23956_),
    .B1(_23959_),
    .X(_23960_));
 sky130_fd_sc_hd__nand3_1 _27239_ (.A(_23956_),
    .B(_23959_),
    .C(_23955_),
    .Y(_23961_));
 sky130_fd_sc_hd__and3_1 _27240_ (.A(_23960_),
    .B(_23961_),
    .C(_22519_),
    .X(_23963_));
 sky130_fd_sc_hd__a21oi_1 _27241_ (.A1(_23960_),
    .A2(_23961_),
    .B1(_22519_),
    .Y(_23964_));
 sky130_fd_sc_hd__nor2_2 _27242_ (.A(_23963_),
    .B(_23964_),
    .Y(_23965_));
 sky130_fd_sc_hd__xnor2_4 _27243_ (.A(_23941_),
    .B(_23965_),
    .Y(_23966_));
 sky130_fd_sc_hd__nand3_1 _27244_ (.A(_22549_),
    .B(_21814_),
    .C(_22546_),
    .Y(_23967_));
 sky130_fd_sc_hd__nand2_1 _27245_ (.A(_23967_),
    .B(_22553_),
    .Y(_23968_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27246_ (.A(_21843_),
    .X(_23969_));
 sky130_fd_sc_hd__buf_2 _27247_ (.A(_21812_),
    .X(_23970_));
 sky130_fd_sc_hd__buf_2 _27248_ (.A(\delay_line[9][10] ),
    .X(_23971_));
 sky130_fd_sc_hd__nor2_1 _27249_ (.A(\delay_line[9][9] ),
    .B(_23971_),
    .Y(_23972_));
 sky130_fd_sc_hd__clkbuf_2 _27250_ (.A(\delay_line[9][9] ),
    .X(_23974_));
 sky130_fd_sc_hd__and2_1 _27251_ (.A(_23974_),
    .B(_23971_),
    .X(_23975_));
 sky130_fd_sc_hd__or2_2 _27252_ (.A(_23972_),
    .B(_23975_),
    .X(_23976_));
 sky130_fd_sc_hd__o21ai_1 _27253_ (.A1(_23969_),
    .A2(_23970_),
    .B1(_23976_),
    .Y(_23977_));
 sky130_fd_sc_hd__buf_1 _27254_ (.A(_23972_),
    .X(_23978_));
 sky130_fd_sc_hd__or4_2 _27255_ (.A(_23969_),
    .B(_23970_),
    .C(_23978_),
    .D(_23975_),
    .X(_23979_));
 sky130_fd_sc_hd__nand2_1 _27256_ (.A(_22441_),
    .B(_22442_),
    .Y(_23980_));
 sky130_fd_sc_hd__a21o_1 _27257_ (.A1(_23977_),
    .A2(_23979_),
    .B1(_23980_),
    .X(_23981_));
 sky130_fd_sc_hd__nand3_1 _27258_ (.A(_23980_),
    .B(_23977_),
    .C(_23979_),
    .Y(_23982_));
 sky130_fd_sc_hd__a32o_1 _27259_ (.A1(_22542_),
    .A2(_22544_),
    .A3(_08668_),
    .B1(_23970_),
    .B2(_20129_),
    .X(_23983_));
 sky130_fd_sc_hd__a21oi_1 _27260_ (.A1(_23981_),
    .A2(_23982_),
    .B1(_23983_),
    .Y(_23985_));
 sky130_fd_sc_hd__and3_1 _27261_ (.A(_23983_),
    .B(_23981_),
    .C(_23982_),
    .X(_23986_));
 sky130_fd_sc_hd__o211ai_2 _27262_ (.A1(_23985_),
    .A2(_23986_),
    .B1(_22451_),
    .C1(_22453_),
    .Y(_23987_));
 sky130_fd_sc_hd__and2_1 _27263_ (.A(_23968_),
    .B(_23987_),
    .X(_23988_));
 sky130_fd_sc_hd__a211o_1 _27264_ (.A1(_22451_),
    .A2(_22453_),
    .B1(_23985_),
    .C1(_23986_),
    .X(_23989_));
 sky130_fd_sc_hd__a21oi_1 _27265_ (.A1(_23987_),
    .A2(_23989_),
    .B1(_23968_),
    .Y(_23990_));
 sky130_fd_sc_hd__a21o_1 _27266_ (.A1(_23988_),
    .A2(_23989_),
    .B1(_23990_),
    .X(_23991_));
 sky130_fd_sc_hd__a32oi_4 _27267_ (.A1(_22540_),
    .A2(_22552_),
    .A3(_22553_),
    .B1(_22557_),
    .B2(_22539_),
    .Y(_23992_));
 sky130_fd_sc_hd__xnor2_1 _27268_ (.A(_23991_),
    .B(_23992_),
    .Y(_23993_));
 sky130_fd_sc_hd__xor2_2 _27269_ (.A(_23966_),
    .B(_23993_),
    .X(_23994_));
 sky130_fd_sc_hd__xor2_2 _27270_ (.A(_23930_),
    .B(_23994_),
    .X(_23996_));
 sky130_fd_sc_hd__nor2_1 _27271_ (.A(_23928_),
    .B(_23996_),
    .Y(_23997_));
 sky130_fd_sc_hd__and2_1 _27272_ (.A(_23928_),
    .B(_23996_),
    .X(_23998_));
 sky130_fd_sc_hd__o2bb2ai_1 _27273_ (.A1_N(_23922_),
    .A2_N(_23926_),
    .B1(_23997_),
    .B2(_23998_),
    .Y(_23999_));
 sky130_fd_sc_hd__nand2_1 _27274_ (.A(_23749_),
    .B(_22427_),
    .Y(_24000_));
 sky130_fd_sc_hd__nor2_1 _27275_ (.A(_22575_),
    .B(_22576_),
    .Y(_24001_));
 sky130_fd_sc_hd__a32oi_1 _27276_ (.A1(_22488_),
    .A2(_22498_),
    .A3(_24000_),
    .B1(_22494_),
    .B2(_24001_),
    .Y(_24002_));
 sky130_fd_sc_hd__a21o_1 _27277_ (.A1(_22559_),
    .A2(_22568_),
    .B1(_23996_),
    .X(_24003_));
 sky130_fd_sc_hd__inv_2 _27278_ (.A(_24003_),
    .Y(_24004_));
 sky130_fd_sc_hd__and3_1 _27279_ (.A(_22559_),
    .B(_22568_),
    .C(_23996_),
    .X(_24005_));
 sky130_fd_sc_hd__clkbuf_2 _27280_ (.A(_23922_),
    .X(_24007_));
 sky130_fd_sc_hd__o211ai_1 _27281_ (.A1(_24004_),
    .A2(_24005_),
    .B1(_24007_),
    .C1(_23926_),
    .Y(_24008_));
 sky130_fd_sc_hd__nand3_1 _27282_ (.A(_23999_),
    .B(_24002_),
    .C(_24008_),
    .Y(_24009_));
 sky130_fd_sc_hd__clkbuf_2 _27283_ (.A(_24009_),
    .X(_24010_));
 sky130_fd_sc_hd__o21a_1 _27284_ (.A1(_21798_),
    .A2(_21828_),
    .B1(_21835_),
    .X(_24011_));
 sky130_fd_sc_hd__a21oi_1 _27285_ (.A1(_22563_),
    .A2(_24011_),
    .B1(_22574_),
    .Y(_24012_));
 sky130_fd_sc_hd__o21bai_2 _27286_ (.A1(_22563_),
    .A2(_24011_),
    .B1_N(_24012_),
    .Y(_24013_));
 sky130_fd_sc_hd__a41o_1 _27287_ (.A1(_03568_),
    .A2(_21971_),
    .A3(_22671_),
    .A4(_22672_),
    .B1(_22682_),
    .X(_24014_));
 sky130_fd_sc_hd__and2b_1 _27288_ (.A_N(\delay_line[3][8] ),
    .B(\delay_line[3][10] ),
    .X(_24015_));
 sky130_fd_sc_hd__clkbuf_2 _27289_ (.A(\delay_line[3][10] ),
    .X(_24016_));
 sky130_fd_sc_hd__or2b_1 _27290_ (.A(_24016_),
    .B_N(_21971_),
    .X(_24018_));
 sky130_fd_sc_hd__nand3b_2 _27291_ (.A_N(_24015_),
    .B(_24018_),
    .C(_22639_),
    .Y(_24019_));
 sky130_fd_sc_hd__and2b_1 _27292_ (.A_N(_24016_),
    .B(_21971_),
    .X(_24020_));
 sky130_fd_sc_hd__o22ai_2 _27293_ (.A1(_18098_),
    .A2(_22640_),
    .B1(_24015_),
    .B2(_24020_),
    .Y(_24021_));
 sky130_fd_sc_hd__and2b_1 _27294_ (.A_N(_19885_),
    .B(net441),
    .X(_24022_));
 sky130_fd_sc_hd__a21oi_1 _27295_ (.A1(_24019_),
    .A2(_24021_),
    .B1(_24022_),
    .Y(_24023_));
 sky130_fd_sc_hd__nand3_1 _27296_ (.A(_24019_),
    .B(_24021_),
    .C(_24022_),
    .Y(_24024_));
 sky130_fd_sc_hd__nor2_1 _27297_ (.A(_22639_),
    .B(_22641_),
    .Y(_24025_));
 sky130_fd_sc_hd__and4bb_1 _27298_ (.A_N(_24023_),
    .B_N(_22643_),
    .C(_24024_),
    .D(_24025_),
    .X(_24026_));
 sky130_fd_sc_hd__and3_1 _27299_ (.A(_24019_),
    .B(_24021_),
    .C(_24022_),
    .X(_24027_));
 sky130_fd_sc_hd__o32a_1 _27300_ (.A1(_22643_),
    .A2(_22639_),
    .A3(_22641_),
    .B1(_24027_),
    .B2(_24023_),
    .X(_24029_));
 sky130_fd_sc_hd__nor2_1 _27301_ (.A(_24026_),
    .B(_24029_),
    .Y(_24030_));
 sky130_fd_sc_hd__xnor2_1 _27302_ (.A(_24014_),
    .B(_24030_),
    .Y(_24031_));
 sky130_fd_sc_hd__o31a_1 _27303_ (.A1(_21968_),
    .A2(_22658_),
    .A3(_22659_),
    .B1(_22661_),
    .X(_24032_));
 sky130_fd_sc_hd__xnor2_1 _27304_ (.A(_24031_),
    .B(_24032_),
    .Y(_24033_));
 sky130_fd_sc_hd__a21oi_2 _27305_ (.A1(_22681_),
    .A2(_22684_),
    .B1(_24033_),
    .Y(_24034_));
 sky130_fd_sc_hd__o311a_1 _27306_ (.A1(_22679_),
    .A2(_22678_),
    .A3(_22682_),
    .B1(_22684_),
    .C1(_24033_),
    .X(_24035_));
 sky130_fd_sc_hd__nor2_2 _27307_ (.A(_24034_),
    .B(_24035_),
    .Y(_24036_));
 sky130_fd_sc_hd__a211oi_1 _27308_ (.A1(_21986_),
    .A2(_21988_),
    .B1(_22634_),
    .C1(_22635_),
    .Y(_24037_));
 sky130_fd_sc_hd__a31oi_2 _27309_ (.A1(_22661_),
    .A2(_22662_),
    .A3(_22637_),
    .B1(_24037_),
    .Y(_24038_));
 sky130_fd_sc_hd__clkbuf_2 _27310_ (.A(\delay_line[5][9] ),
    .X(_24040_));
 sky130_fd_sc_hd__nand2_1 _27311_ (.A(_21962_),
    .B(_24040_),
    .Y(_24041_));
 sky130_fd_sc_hd__or2_1 _27312_ (.A(_24040_),
    .B(_21962_),
    .X(_24042_));
 sky130_fd_sc_hd__a21oi_1 _27313_ (.A1(_24041_),
    .A2(_24042_),
    .B1(_19045_),
    .Y(_24043_));
 sky130_fd_sc_hd__and3_1 _27314_ (.A(_24042_),
    .B(_19045_),
    .C(_24041_),
    .X(_24044_));
 sky130_fd_sc_hd__nand2_1 _27315_ (.A(_09217_),
    .B(net430),
    .Y(_24045_));
 sky130_fd_sc_hd__or2_1 _27316_ (.A(net430),
    .B(_09217_),
    .X(_24046_));
 sky130_fd_sc_hd__nand2_1 _27317_ (.A(_24045_),
    .B(_24046_),
    .Y(_24047_));
 sky130_fd_sc_hd__a21o_1 _27318_ (.A1(_22648_),
    .A2(_22650_),
    .B1(_24047_),
    .X(_24048_));
 sky130_fd_sc_hd__nand3_1 _27319_ (.A(_22648_),
    .B(_22651_),
    .C(_24047_),
    .Y(_24049_));
 sky130_fd_sc_hd__and3b_1 _27320_ (.A_N(_22653_),
    .B(_24048_),
    .C(_24049_),
    .X(_24051_));
 sky130_fd_sc_hd__a32oi_4 _27321_ (.A1(_22654_),
    .A2(_22651_),
    .A3(_22652_),
    .B1(_24048_),
    .B2(_24049_),
    .Y(_24052_));
 sky130_fd_sc_hd__nor4_1 _27322_ (.A(_24043_),
    .B(_24044_),
    .C(_24051_),
    .D(_24052_),
    .Y(_24053_));
 sky130_fd_sc_hd__or2_1 _27323_ (.A(_24043_),
    .B(_24044_),
    .X(_24054_));
 sky130_fd_sc_hd__o21ai_1 _27324_ (.A1(_24051_),
    .A2(_24052_),
    .B1(_24054_),
    .Y(_24055_));
 sky130_fd_sc_hd__and2b_1 _27325_ (.A_N(_24053_),
    .B(_24055_),
    .X(_24056_));
 sky130_fd_sc_hd__a31o_1 _27326_ (.A1(_19905_),
    .A2(net273),
    .A3(_22629_),
    .B1(_22635_),
    .X(_24057_));
 sky130_fd_sc_hd__buf_2 _27327_ (.A(net428),
    .X(_24058_));
 sky130_fd_sc_hd__clkbuf_2 _27328_ (.A(_21979_),
    .X(_24059_));
 sky130_fd_sc_hd__or2_1 _27329_ (.A(_24058_),
    .B(_24059_),
    .X(_24060_));
 sky130_fd_sc_hd__clkbuf_2 _27330_ (.A(\delay_line[6][10] ),
    .X(_24062_));
 sky130_fd_sc_hd__nor2_1 _27331_ (.A(_22604_),
    .B(_24062_),
    .Y(_24063_));
 sky130_fd_sc_hd__and2_1 _27332_ (.A(_22606_),
    .B(\delay_line[6][10] ),
    .X(_24064_));
 sky130_fd_sc_hd__o21a_1 _27333_ (.A1(_24063_),
    .A2(_24064_),
    .B1(_22628_),
    .X(_24065_));
 sky130_fd_sc_hd__nor3_2 _27334_ (.A(_22628_),
    .B(_24063_),
    .C(_24064_),
    .Y(_24066_));
 sky130_fd_sc_hd__o211ai_2 _27335_ (.A1(_24065_),
    .A2(_24066_),
    .B1(_22603_),
    .C1(_22605_),
    .Y(_24067_));
 sky130_fd_sc_hd__a211o_2 _27336_ (.A1(_22603_),
    .A2(_22605_),
    .B1(_24065_),
    .C1(_24066_),
    .X(_24068_));
 sky130_fd_sc_hd__a22o_1 _27337_ (.A1(_24060_),
    .A2(_18082_),
    .B1(_24067_),
    .B2(_24068_),
    .X(_24069_));
 sky130_fd_sc_hd__o2111ai_4 _27338_ (.A1(_24058_),
    .A2(_24059_),
    .B1(_18082_),
    .C1(_24068_),
    .D1(_24067_),
    .Y(_24070_));
 sky130_fd_sc_hd__nand2_1 _27339_ (.A(_24069_),
    .B(_24070_),
    .Y(_24071_));
 sky130_fd_sc_hd__xnor2_2 _27340_ (.A(_24057_),
    .B(_24071_),
    .Y(_24073_));
 sky130_fd_sc_hd__xnor2_2 _27341_ (.A(_24056_),
    .B(_24073_),
    .Y(_24074_));
 sky130_fd_sc_hd__nor2_1 _27342_ (.A(_24038_),
    .B(_24074_),
    .Y(_24075_));
 sky130_fd_sc_hd__nand2_1 _27343_ (.A(_24074_),
    .B(_24038_),
    .Y(_24076_));
 sky130_fd_sc_hd__or2b_2 _27344_ (.A(_24075_),
    .B_N(_24076_),
    .X(_24077_));
 sky130_fd_sc_hd__xor2_4 _27345_ (.A(_24036_),
    .B(_24077_),
    .X(_24078_));
 sky130_fd_sc_hd__a31o_1 _27346_ (.A1(_21928_),
    .A2(_21929_),
    .A3(_22618_),
    .B1(_22617_),
    .X(_24079_));
 sky130_fd_sc_hd__o31ai_1 _27347_ (.A1(_21864_),
    .A2(_22608_),
    .A3(_22609_),
    .B1(_22614_),
    .Y(_24080_));
 sky130_fd_sc_hd__o21ba_1 _27348_ (.A1(_22518_),
    .A2(_22519_),
    .B1_N(_21875_),
    .X(_24081_));
 sky130_fd_sc_hd__o21a_1 _27349_ (.A1(_22531_),
    .A2(_24081_),
    .B1(_22520_),
    .X(_24082_));
 sky130_fd_sc_hd__clkbuf_2 _27350_ (.A(_22596_),
    .X(_24084_));
 sky130_fd_sc_hd__o21ai_1 _27351_ (.A1(_11965_),
    .A2(_18025_),
    .B1(_08965_),
    .Y(_24085_));
 sky130_fd_sc_hd__nor2_1 _27352_ (.A(_21906_),
    .B(_21910_),
    .Y(_24086_));
 sky130_fd_sc_hd__nor2_1 _27353_ (.A(_11965_),
    .B(_03128_),
    .Y(_24087_));
 sky130_fd_sc_hd__a211o_2 _27354_ (.A1(_22593_),
    .A2(_24085_),
    .B1(_24086_),
    .C1(_24087_),
    .X(_24088_));
 sky130_fd_sc_hd__o221ai_4 _27355_ (.A1(_22591_),
    .A2(_22592_),
    .B1(_24086_),
    .B2(_24087_),
    .C1(_22593_),
    .Y(_24089_));
 sky130_fd_sc_hd__a22o_1 _27356_ (.A1(_24084_),
    .A2(_00062_),
    .B1(_24088_),
    .B2(_24089_),
    .X(_24090_));
 sky130_fd_sc_hd__clkbuf_2 _27357_ (.A(\delay_line[7][10] ),
    .X(_24091_));
 sky130_fd_sc_hd__clkbuf_2 _27358_ (.A(\delay_line[7][6] ),
    .X(_24092_));
 sky130_fd_sc_hd__xor2_2 _27359_ (.A(_18025_),
    .B(_24092_),
    .X(_24093_));
 sky130_fd_sc_hd__xor2_1 _27360_ (.A(_24091_),
    .B(_24093_),
    .X(_24095_));
 sky130_fd_sc_hd__nand4_4 _27361_ (.A(_00073_),
    .B(_24088_),
    .C(_24084_),
    .D(_24089_),
    .Y(_24096_));
 sky130_fd_sc_hd__and3_1 _27362_ (.A(_24090_),
    .B(_24095_),
    .C(_24096_),
    .X(_24097_));
 sky130_fd_sc_hd__a21oi_1 _27363_ (.A1(_24096_),
    .A2(_24090_),
    .B1(_24095_),
    .Y(_24098_));
 sky130_fd_sc_hd__a2111o_1 _27364_ (.A1(_20105_),
    .A2(_21872_),
    .B1(_22530_),
    .C1(_24097_),
    .D1(_24098_),
    .X(_24099_));
 sky130_fd_sc_hd__o22ai_2 _27365_ (.A1(_22530_),
    .A2(_22522_),
    .B1(_24098_),
    .B2(_24097_),
    .Y(_24100_));
 sky130_fd_sc_hd__a32o_1 _27366_ (.A1(_22595_),
    .A2(_22605_),
    .A3(_22607_),
    .B1(_24099_),
    .B2(_24100_),
    .X(_24101_));
 sky130_fd_sc_hd__nand3_1 _27367_ (.A(_24099_),
    .B(_24100_),
    .C(_22608_),
    .Y(_24102_));
 sky130_fd_sc_hd__nand2_1 _27368_ (.A(_24101_),
    .B(_24102_),
    .Y(_24103_));
 sky130_fd_sc_hd__or2_1 _27369_ (.A(_24082_),
    .B(_24103_),
    .X(_24104_));
 sky130_fd_sc_hd__nand2_1 _27370_ (.A(_24103_),
    .B(_24082_),
    .Y(_24106_));
 sky130_fd_sc_hd__nand3_1 _27371_ (.A(_24080_),
    .B(_24104_),
    .C(_24106_),
    .Y(_24107_));
 sky130_fd_sc_hd__a21o_1 _27372_ (.A1(_24104_),
    .A2(_24106_),
    .B1(_24080_),
    .X(_24108_));
 sky130_fd_sc_hd__nand2_1 _27373_ (.A(_24107_),
    .B(_24108_),
    .Y(_24109_));
 sky130_fd_sc_hd__xnor2_2 _27374_ (.A(_24079_),
    .B(_24109_),
    .Y(_24110_));
 sky130_fd_sc_hd__nand2_1 _27375_ (.A(_24078_),
    .B(_24110_),
    .Y(_24111_));
 sky130_fd_sc_hd__or2_1 _27376_ (.A(_24078_),
    .B(_24110_),
    .X(_24112_));
 sky130_fd_sc_hd__nand3_2 _27377_ (.A(_24013_),
    .B(_24111_),
    .C(_24112_),
    .Y(_24113_));
 sky130_fd_sc_hd__a21oi_1 _27378_ (.A1(_24111_),
    .A2(_24112_),
    .B1(_24013_),
    .Y(_24114_));
 sky130_fd_sc_hd__a21oi_2 _27379_ (.A1(_22624_),
    .A2(_22700_),
    .B1(_24114_),
    .Y(_24115_));
 sky130_fd_sc_hd__inv_2 _27380_ (.A(_24113_),
    .Y(_24117_));
 sky130_fd_sc_hd__o221a_1 _27381_ (.A1(_22696_),
    .A2(_22626_),
    .B1(_24114_),
    .B2(_24117_),
    .C1(_22624_),
    .X(_24118_));
 sky130_fd_sc_hd__a21oi_2 _27382_ (.A1(_24113_),
    .A2(_24115_),
    .B1(_24118_),
    .Y(_24119_));
 sky130_fd_sc_hd__nand2_1 _27383_ (.A(_24010_),
    .B(_24119_),
    .Y(_24120_));
 sky130_fd_sc_hd__and3_1 _27384_ (.A(_22488_),
    .B(_22498_),
    .C(_24000_),
    .X(_24121_));
 sky130_fd_sc_hd__nand2_1 _27385_ (.A(_22427_),
    .B(_22432_),
    .Y(_24122_));
 sky130_fd_sc_hd__a21oi_1 _27386_ (.A1(_24122_),
    .A2(_22495_),
    .B1(_22488_),
    .Y(_24123_));
 sky130_fd_sc_hd__a21boi_2 _27387_ (.A1(_24123_),
    .A2(_22493_),
    .B1_N(_24001_),
    .Y(_24124_));
 sky130_fd_sc_hd__inv_2 _27388_ (.A(_24007_),
    .Y(_24125_));
 sky130_fd_sc_hd__o21ai_2 _27389_ (.A1(_23997_),
    .A2(_23998_),
    .B1(_23926_),
    .Y(_24126_));
 sky130_fd_sc_hd__o2bb2ai_2 _27390_ (.A1_N(_24007_),
    .A2_N(_23926_),
    .B1(_24004_),
    .B2(_24005_),
    .Y(_24128_));
 sky130_fd_sc_hd__o221a_2 _27391_ (.A1(_24121_),
    .A2(_24124_),
    .B1(_24125_),
    .B2(_24126_),
    .C1(_24128_),
    .X(_24129_));
 sky130_fd_sc_hd__nand2_1 _27392_ (.A(_22580_),
    .B(_22705_),
    .Y(_24130_));
 sky130_fd_sc_hd__nand2_1 _27393_ (.A(_22584_),
    .B(_24130_),
    .Y(_24131_));
 sky130_fd_sc_hd__o211ai_2 _27394_ (.A1(_23997_),
    .A2(_23998_),
    .B1(_24007_),
    .C1(_23926_),
    .Y(_24132_));
 sky130_fd_sc_hd__o211ai_4 _27395_ (.A1(_24121_),
    .A2(_24124_),
    .B1(_24132_),
    .C1(_24128_),
    .Y(_24133_));
 sky130_fd_sc_hd__a21o_1 _27396_ (.A1(_24133_),
    .A2(_24009_),
    .B1(_24119_),
    .X(_24134_));
 sky130_fd_sc_hd__o211ai_4 _27397_ (.A1(_24120_),
    .A2(_24129_),
    .B1(_24131_),
    .C1(_24134_),
    .Y(_24135_));
 sky130_fd_sc_hd__a21o_1 _27398_ (.A1(_24113_),
    .A2(_24115_),
    .B1(_24118_),
    .X(_24136_));
 sky130_fd_sc_hd__a21o_1 _27399_ (.A1(_24133_),
    .A2(_24010_),
    .B1(_24136_),
    .X(_24137_));
 sky130_fd_sc_hd__nand3_1 _27400_ (.A(_24136_),
    .B(_24133_),
    .C(_24010_),
    .Y(_24139_));
 sky130_fd_sc_hd__a32oi_4 _27401_ (.A1(_22581_),
    .A2(_22582_),
    .A3(_22583_),
    .B1(_22580_),
    .B2(_22705_),
    .Y(_24140_));
 sky130_fd_sc_hd__nand3_2 _27402_ (.A(_24137_),
    .B(_24139_),
    .C(_24140_),
    .Y(_24141_));
 sky130_fd_sc_hd__nand2_1 _27403_ (.A(_24135_),
    .B(_24141_),
    .Y(_24142_));
 sky130_fd_sc_hd__nand2_1 _27404_ (.A(_22585_),
    .B(_22702_),
    .Y(_24143_));
 sky130_fd_sc_hd__a21boi_2 _27405_ (.A1(_22228_),
    .A2(_22257_),
    .B1_N(_22261_),
    .Y(_24144_));
 sky130_fd_sc_hd__nand2_1 _27406_ (.A(_22254_),
    .B(_22258_),
    .Y(_24145_));
 sky130_fd_sc_hd__nand3_1 _27407_ (.A(_22670_),
    .B(_22691_),
    .C(_22692_),
    .Y(_24146_));
 sky130_fd_sc_hd__nor2_1 _27408_ (.A(_22231_),
    .B(_22233_),
    .Y(_24147_));
 sky130_fd_sc_hd__nor2_1 _27409_ (.A(_20193_),
    .B(net449),
    .Y(_24148_));
 sky130_fd_sc_hd__and2_1 _27410_ (.A(_20193_),
    .B(net449),
    .X(_24150_));
 sky130_fd_sc_hd__nor2_1 _27411_ (.A(_24148_),
    .B(_24150_),
    .Y(_24151_));
 sky130_fd_sc_hd__nand2_1 _27412_ (.A(net440),
    .B(_24151_),
    .Y(_24152_));
 sky130_fd_sc_hd__o21bai_1 _27413_ (.A1(_24148_),
    .A2(_24150_),
    .B1_N(net440),
    .Y(_24153_));
 sky130_fd_sc_hd__nand3b_1 _27414_ (.A_N(_22238_),
    .B(_24152_),
    .C(_24153_),
    .Y(_24154_));
 sky130_fd_sc_hd__a21bo_1 _27415_ (.A1(_24152_),
    .A2(_24153_),
    .B1_N(_22238_),
    .X(_24155_));
 sky130_fd_sc_hd__buf_1 _27416_ (.A(_22023_),
    .X(_24156_));
 sky130_fd_sc_hd__buf_1 _27417_ (.A(_22235_),
    .X(_24157_));
 sky130_fd_sc_hd__o21a_1 _27418_ (.A1(_24156_),
    .A2(_24157_),
    .B1(_22232_),
    .X(_24158_));
 sky130_fd_sc_hd__nor3_1 _27419_ (.A(_24156_),
    .B(_24157_),
    .C(_22232_),
    .Y(_24159_));
 sky130_fd_sc_hd__o2bb2ai_1 _27420_ (.A1_N(_24154_),
    .A2_N(_24155_),
    .B1(_24158_),
    .B2(_24159_),
    .Y(_24161_));
 sky130_fd_sc_hd__o21a_1 _27421_ (.A1(_24156_),
    .A2(_24157_),
    .B1(_22230_),
    .X(_24162_));
 sky130_fd_sc_hd__nor3_1 _27422_ (.A(_24156_),
    .B(_24157_),
    .C(_22230_),
    .Y(_24163_));
 sky130_fd_sc_hd__o211ai_2 _27423_ (.A1(_24162_),
    .A2(_24163_),
    .B1(_24154_),
    .C1(_24155_),
    .Y(_24164_));
 sky130_fd_sc_hd__o2111a_1 _27424_ (.A1(_22027_),
    .A2(_22021_),
    .B1(_19051_),
    .C1(_22238_),
    .D1(_22240_),
    .X(_24165_));
 sky130_fd_sc_hd__a221o_1 _27425_ (.A1(_22242_),
    .A2(_24147_),
    .B1(_24161_),
    .B2(_24164_),
    .C1(_24165_),
    .X(_24166_));
 sky130_fd_sc_hd__and3_1 _27426_ (.A(_22242_),
    .B(_24147_),
    .C(_22241_),
    .X(_24167_));
 sky130_fd_sc_hd__o211ai_2 _27427_ (.A1(_24165_),
    .A2(_24167_),
    .B1(_24164_),
    .C1(_24161_),
    .Y(_24168_));
 sky130_fd_sc_hd__nand3b_1 _27428_ (.A_N(_22231_),
    .B(_24166_),
    .C(_24168_),
    .Y(_24169_));
 sky130_fd_sc_hd__a221o_1 _27429_ (.A1(_22034_),
    .A2(_22230_),
    .B1(_24166_),
    .B2(_24168_),
    .C1(_22027_),
    .X(_24170_));
 sky130_fd_sc_hd__nand4_1 _27430_ (.A(_22692_),
    .B(_24146_),
    .C(_24169_),
    .D(_24170_),
    .Y(_24172_));
 sky130_fd_sc_hd__a22o_1 _27431_ (.A1(_22692_),
    .A2(_24146_),
    .B1(_24169_),
    .B2(_24170_),
    .X(_24173_));
 sky130_fd_sc_hd__a22oi_1 _27432_ (.A1(_22247_),
    .A2(_22249_),
    .B1(_24172_),
    .B2(_24173_),
    .Y(_24174_));
 sky130_fd_sc_hd__o31ai_1 _27433_ (.A1(_22693_),
    .A2(_22694_),
    .A3(_22669_),
    .B1(_22667_),
    .Y(_24175_));
 sky130_fd_sc_hd__and4_1 _27434_ (.A(_22247_),
    .B(_22249_),
    .C(_24172_),
    .D(_24173_),
    .X(_24176_));
 sky130_fd_sc_hd__nor3_1 _27435_ (.A(_24174_),
    .B(_24175_),
    .C(_24176_),
    .Y(_24177_));
 sky130_fd_sc_hd__o21ai_1 _27436_ (.A1(_24176_),
    .A2(_24174_),
    .B1(_24175_),
    .Y(_24178_));
 sky130_fd_sc_hd__and2b_1 _27437_ (.A_N(_24177_),
    .B(_24178_),
    .X(_24179_));
 sky130_fd_sc_hd__xnor2_1 _27438_ (.A(_24145_),
    .B(_24179_),
    .Y(_24180_));
 sky130_fd_sc_hd__xnor2_1 _27439_ (.A(_24144_),
    .B(_24180_),
    .Y(_24181_));
 sky130_fd_sc_hd__and3_2 _27440_ (.A(_22701_),
    .B(_24143_),
    .C(_24181_),
    .X(_24183_));
 sky130_fd_sc_hd__a21oi_1 _27441_ (.A1(_22701_),
    .A2(_24143_),
    .B1(_24181_),
    .Y(_24184_));
 sky130_fd_sc_hd__a21oi_2 _27442_ (.A1(_22227_),
    .A2(_22263_),
    .B1(_24184_),
    .Y(_24185_));
 sky130_fd_sc_hd__nor2_1 _27443_ (.A(_24183_),
    .B(_24185_),
    .Y(_24186_));
 sky130_fd_sc_hd__o211a_1 _27444_ (.A1(_24184_),
    .A2(_24183_),
    .B1(_22227_),
    .C1(_22263_),
    .X(_24187_));
 sky130_fd_sc_hd__o21ba_1 _27445_ (.A1(_24183_),
    .A2(_24186_),
    .B1_N(_24187_),
    .X(_24188_));
 sky130_fd_sc_hd__nand2_1 _27446_ (.A(_24142_),
    .B(_24188_),
    .Y(_24189_));
 sky130_fd_sc_hd__o21ai_1 _27447_ (.A1(_22716_),
    .A2(_22711_),
    .B1(_22717_),
    .Y(_24190_));
 sky130_fd_sc_hd__nand3b_1 _27448_ (.A_N(_24188_),
    .B(_24135_),
    .C(_24141_),
    .Y(_24191_));
 sky130_fd_sc_hd__nand3_2 _27449_ (.A(_24189_),
    .B(_24190_),
    .C(_24191_),
    .Y(_24192_));
 sky130_fd_sc_hd__clkbuf_2 _27450_ (.A(_24192_),
    .X(_24194_));
 sky130_fd_sc_hd__nand2_2 _27451_ (.A(_24135_),
    .B(_24188_),
    .Y(_24195_));
 sky130_fd_sc_hd__and3_2 _27452_ (.A(_24137_),
    .B(_24139_),
    .C(_24140_),
    .X(_24196_));
 sky130_fd_sc_hd__o21ai_1 _27453_ (.A1(_22722_),
    .A2(_22723_),
    .B1(_22717_),
    .Y(_24197_));
 sky130_fd_sc_hd__nand2_1 _27454_ (.A(_22715_),
    .B(_24197_),
    .Y(_24198_));
 sky130_fd_sc_hd__a21o_1 _27455_ (.A1(_24135_),
    .A2(_24141_),
    .B1(_24188_),
    .X(_24199_));
 sky130_fd_sc_hd__o211ai_4 _27456_ (.A1(_24195_),
    .A2(_24196_),
    .B1(_24198_),
    .C1(_24199_),
    .Y(_24200_));
 sky130_fd_sc_hd__o211a_1 _27457_ (.A1(_22720_),
    .A2(_23747_),
    .B1(_24194_),
    .C1(_24200_),
    .X(_24201_));
 sky130_fd_sc_hd__nor2_1 _27458_ (.A(_22223_),
    .B(_22720_),
    .Y(_24202_));
 sky130_fd_sc_hd__a31o_1 _27459_ (.A1(_22224_),
    .A2(_22225_),
    .A3(_22264_),
    .B1(_24202_),
    .X(_24203_));
 sky130_fd_sc_hd__a21boi_1 _27460_ (.A1(_24192_),
    .A2(_24200_),
    .B1_N(_24203_),
    .Y(_24205_));
 sky130_fd_sc_hd__clkbuf_2 _27461_ (.A(_22733_),
    .X(_24206_));
 sky130_fd_sc_hd__o21a_1 _27462_ (.A1(_22737_),
    .A2(_22719_),
    .B1(_24206_),
    .X(_24207_));
 sky130_fd_sc_hd__o21ai_2 _27463_ (.A1(_24201_),
    .A2(_24205_),
    .B1(_24207_),
    .Y(_24208_));
 sky130_fd_sc_hd__o21ai_4 _27464_ (.A1(_22737_),
    .A2(_22719_),
    .B1(_24206_),
    .Y(_24209_));
 sky130_fd_sc_hd__o211ai_4 _27465_ (.A1(_22720_),
    .A2(_23747_),
    .B1(_24192_),
    .C1(_24200_),
    .Y(_24210_));
 sky130_fd_sc_hd__nand2_1 _27466_ (.A(_24192_),
    .B(_24200_),
    .Y(_24211_));
 sky130_fd_sc_hd__nand2_1 _27467_ (.A(_24211_),
    .B(_24203_),
    .Y(_24212_));
 sky130_fd_sc_hd__nand3_4 _27468_ (.A(_24209_),
    .B(_24210_),
    .C(_24212_),
    .Y(_24213_));
 sky130_fd_sc_hd__nand2_1 _27469_ (.A(_24208_),
    .B(_24213_),
    .Y(_24214_));
 sky130_fd_sc_hd__o211ai_4 _27470_ (.A1(_23745_),
    .A2(_22729_),
    .B1(_23746_),
    .C1(_24214_),
    .Y(_24216_));
 sky130_fd_sc_hd__nand2_1 _27471_ (.A(_24210_),
    .B(_24212_),
    .Y(_24217_));
 sky130_fd_sc_hd__a31oi_1 _27472_ (.A1(_22713_),
    .A2(_22724_),
    .A3(_22725_),
    .B1(_22726_),
    .Y(_24218_));
 sky130_fd_sc_hd__a2bb2oi_1 _27473_ (.A1_N(_22730_),
    .A2_N(_22069_),
    .B1(_22739_),
    .B2(_24206_),
    .Y(_24219_));
 sky130_fd_sc_hd__a211oi_1 _27474_ (.A1(_24218_),
    .A2(_22739_),
    .B1(_22728_),
    .C1(_24219_),
    .Y(_24220_));
 sky130_fd_sc_hd__a21oi_1 _27475_ (.A1(_24217_),
    .A2(_24207_),
    .B1(_24220_),
    .Y(_24221_));
 sky130_fd_sc_hd__or3_1 _27476_ (.A(_22083_),
    .B(_22081_),
    .C(_22095_),
    .X(_24222_));
 sky130_fd_sc_hd__o211ai_2 _27477_ (.A1(_22090_),
    .A2(_22089_),
    .B1(_22741_),
    .C1(_24222_),
    .Y(_24223_));
 sky130_fd_sc_hd__nand3_4 _27478_ (.A(_24221_),
    .B(_24223_),
    .C(_24213_),
    .Y(_24224_));
 sky130_fd_sc_hd__buf_2 _27479_ (.A(net348),
    .X(_24225_));
 sky130_fd_sc_hd__a21oi_4 _27480_ (.A1(_24216_),
    .A2(_24224_),
    .B1(_24225_),
    .Y(_24227_));
 sky130_fd_sc_hd__a21oi_1 _27481_ (.A1(_22739_),
    .A2(_24206_),
    .B1(_22726_),
    .Y(_24228_));
 sky130_fd_sc_hd__o211a_1 _27482_ (.A1(_22730_),
    .A2(_22069_),
    .B1(_22739_),
    .C1(_24206_),
    .X(_24229_));
 sky130_fd_sc_hd__nor2_1 _27483_ (.A(_24228_),
    .B(_24229_),
    .Y(_24230_));
 sky130_fd_sc_hd__a21oi_4 _27484_ (.A1(_24230_),
    .A2(_22728_),
    .B1(_22221_),
    .Y(_24231_));
 sky130_fd_sc_hd__nand3_4 _27485_ (.A(_22736_),
    .B(_24208_),
    .C(_24213_),
    .Y(_24232_));
 sky130_fd_sc_hd__o211ai_4 _27486_ (.A1(_24231_),
    .A2(_24232_),
    .B1(_24225_),
    .C1(_24216_),
    .Y(_24233_));
 sky130_fd_sc_hd__buf_1 _27487_ (.A(_22749_),
    .X(_24234_));
 sky130_fd_sc_hd__nand2_1 _27488_ (.A(_24233_),
    .B(_24234_),
    .Y(_24235_));
 sky130_fd_sc_hd__nor2_2 _27489_ (.A(_24227_),
    .B(_24235_),
    .Y(_24236_));
 sky130_fd_sc_hd__inv_2 _27490_ (.A(net348),
    .Y(_24238_));
 sky130_fd_sc_hd__o21ai_2 _27491_ (.A1(_24231_),
    .A2(_24232_),
    .B1(_24216_),
    .Y(_24239_));
 sky130_fd_sc_hd__nand2_1 _27492_ (.A(_24238_),
    .B(_24239_),
    .Y(_24240_));
 sky130_fd_sc_hd__clkbuf_2 _27493_ (.A(_24234_),
    .X(_24241_));
 sky130_fd_sc_hd__a21oi_1 _27494_ (.A1(_24240_),
    .A2(_24233_),
    .B1(_24241_),
    .Y(_24242_));
 sky130_fd_sc_hd__a21bo_2 _27495_ (.A1(_23476_),
    .A2(_23477_),
    .B1_N(_23463_),
    .X(_24243_));
 sky130_fd_sc_hd__o21bai_4 _27496_ (.A1(_24236_),
    .A2(_24242_),
    .B1_N(_24243_),
    .Y(_24244_));
 sky130_fd_sc_hd__and3_2 _27497_ (.A(_24216_),
    .B(_24224_),
    .C(_24225_),
    .X(_24245_));
 sky130_fd_sc_hd__o21bai_1 _27498_ (.A1(_24227_),
    .A2(_24245_),
    .B1_N(_24234_),
    .Y(_24246_));
 sky130_fd_sc_hd__o211ai_2 _27499_ (.A1(_24235_),
    .A2(_24227_),
    .B1(_24243_),
    .C1(_24246_),
    .Y(_24247_));
 sky130_fd_sc_hd__nand2_1 _27500_ (.A(_24244_),
    .B(_24247_),
    .Y(_24249_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27501_ (.A(_22761_),
    .X(_24250_));
 sky130_fd_sc_hd__buf_2 _27502_ (.A(_24250_),
    .X(_24251_));
 sky130_fd_sc_hd__clkbuf_2 _27503_ (.A(_24234_),
    .X(_24252_));
 sky130_fd_sc_hd__o211a_2 _27504_ (.A1(_24250_),
    .A2(_24234_),
    .B1(_22742_),
    .C1(_22746_),
    .X(_24253_));
 sky130_fd_sc_hd__a21oi_2 _27505_ (.A1(_24251_),
    .A2(_24252_),
    .B1(_24253_),
    .Y(_24254_));
 sky130_fd_sc_hd__nand2_1 _27506_ (.A(_24249_),
    .B(_24254_),
    .Y(_24255_));
 sky130_fd_sc_hd__buf_2 _27507_ (.A(_22748_),
    .X(_24256_));
 sky130_fd_sc_hd__buf_2 _27508_ (.A(_24247_),
    .X(_24257_));
 sky130_fd_sc_hd__o211ai_4 _27509_ (.A1(_24256_),
    .A2(_24253_),
    .B1(_24244_),
    .C1(_24257_),
    .Y(_24258_));
 sky130_fd_sc_hd__nand2_1 _27510_ (.A(_24255_),
    .B(_24258_),
    .Y(_24260_));
 sky130_fd_sc_hd__a21o_1 _27511_ (.A1(_23481_),
    .A2(_23533_),
    .B1(_23532_),
    .X(_24261_));
 sky130_fd_sc_hd__inv_2 _27512_ (.A(_24261_),
    .Y(_24262_));
 sky130_fd_sc_hd__a32o_1 _27513_ (.A1(_22220_),
    .A2(_22751_),
    .A3(_22755_),
    .B1(_22759_),
    .B2(_22763_),
    .X(_24263_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27514_ (.A(_24263_),
    .X(_24264_));
 sky130_fd_sc_hd__a21boi_1 _27515_ (.A1(_24260_),
    .A2(_24262_),
    .B1_N(_24264_),
    .Y(_24265_));
 sky130_fd_sc_hd__and2_1 _27516_ (.A(_23481_),
    .B(_23533_),
    .X(_24266_));
 sky130_fd_sc_hd__o211ai_4 _27517_ (.A1(_23532_),
    .A2(_24266_),
    .B1(_24255_),
    .C1(_24258_),
    .Y(_24267_));
 sky130_fd_sc_hd__o32a_2 _27518_ (.A1(_22218_),
    .A2(_22764_),
    .A3(_22766_),
    .B1(_22770_),
    .B2(_22773_),
    .X(_24268_));
 sky130_fd_sc_hd__a21boi_2 _27519_ (.A1(_24244_),
    .A2(_24257_),
    .B1_N(_24254_),
    .Y(_24269_));
 sky130_fd_sc_hd__o211a_2 _27520_ (.A1(_24256_),
    .A2(_24253_),
    .B1(_24244_),
    .C1(_24247_),
    .X(_24271_));
 sky130_fd_sc_hd__o21bai_4 _27521_ (.A1(_24269_),
    .A2(_24271_),
    .B1_N(_24261_),
    .Y(_24272_));
 sky130_fd_sc_hd__a21oi_2 _27522_ (.A1(_24272_),
    .A2(_24267_),
    .B1(_24264_),
    .Y(_24273_));
 sky130_fd_sc_hd__a211oi_2 _27523_ (.A1(_24265_),
    .A2(_24267_),
    .B1(_24268_),
    .C1(_24273_),
    .Y(_24274_));
 sky130_fd_sc_hd__a21o_1 _27524_ (.A1(_24272_),
    .A2(_24267_),
    .B1(_24264_),
    .X(_24275_));
 sky130_fd_sc_hd__o2bb2ai_1 _27525_ (.A1_N(_24254_),
    .A2_N(_24249_),
    .B1(_23532_),
    .B2(_24266_),
    .Y(_24276_));
 sky130_fd_sc_hd__o211ai_2 _27526_ (.A1(_24271_),
    .A2(_24276_),
    .B1(_24272_),
    .C1(_24264_),
    .Y(_24277_));
 sky130_fd_sc_hd__o21ai_4 _27527_ (.A1(_22773_),
    .A2(_22770_),
    .B1(_22774_),
    .Y(_24278_));
 sky130_fd_sc_hd__a21oi_2 _27528_ (.A1(_24275_),
    .A2(_24277_),
    .B1(_24278_),
    .Y(_24279_));
 sky130_fd_sc_hd__nor2_1 _27529_ (.A(_00755_),
    .B(_10635_),
    .Y(_24280_));
 sky130_fd_sc_hd__nand2_1 _27530_ (.A(_17895_),
    .B(_07909_),
    .Y(_24282_));
 sky130_fd_sc_hd__and2_1 _27531_ (.A(_22129_),
    .B(_22761_),
    .X(_24283_));
 sky130_fd_sc_hd__nor2_1 _27532_ (.A(_22130_),
    .B(_24250_),
    .Y(_24284_));
 sky130_fd_sc_hd__or3b_2 _27533_ (.A(_24283_),
    .B(_24284_),
    .C_N(_22778_),
    .X(_24285_));
 sky130_fd_sc_hd__clkbuf_2 _27534_ (.A(_22760_),
    .X(_24286_));
 sky130_fd_sc_hd__a2bb2o_1 _27535_ (.A1_N(_24283_),
    .A2_N(_24284_),
    .B1(_19849_),
    .B2(_24286_),
    .X(_24287_));
 sky130_fd_sc_hd__and4b_1 _27536_ (.A_N(_24280_),
    .B(_24282_),
    .C(_24285_),
    .D(_24287_),
    .X(_24288_));
 sky130_fd_sc_hd__and2_1 _27537_ (.A(_23513_),
    .B(_07909_),
    .X(_24289_));
 sky130_fd_sc_hd__nand2_1 _27538_ (.A(_24285_),
    .B(_24287_),
    .Y(_24290_));
 sky130_fd_sc_hd__o21a_1 _27539_ (.A1(_24280_),
    .A2(_24289_),
    .B1(_24290_),
    .X(_24291_));
 sky130_fd_sc_hd__nor2_1 _27540_ (.A(_24288_),
    .B(_24291_),
    .Y(_24293_));
 sky130_fd_sc_hd__o21ai_2 _27541_ (.A1(_24274_),
    .A2(_24279_),
    .B1(_24293_),
    .Y(_24294_));
 sky130_fd_sc_hd__inv_2 _27542_ (.A(_23542_),
    .Y(_24295_));
 sky130_fd_sc_hd__nor2_1 _27543_ (.A(_23539_),
    .B(_24295_),
    .Y(_24296_));
 sky130_fd_sc_hd__nand3_2 _27544_ (.A(_24278_),
    .B(_24275_),
    .C(_24277_),
    .Y(_24297_));
 sky130_fd_sc_hd__o211a_1 _27545_ (.A1(_24276_),
    .A2(_24271_),
    .B1(_24264_),
    .C1(_24272_),
    .X(_24298_));
 sky130_fd_sc_hd__o21bai_4 _27546_ (.A1(_24273_),
    .A2(_24298_),
    .B1_N(_24278_),
    .Y(_24299_));
 sky130_fd_sc_hd__o211ai_2 _27547_ (.A1(_24288_),
    .A2(_24291_),
    .B1(_24297_),
    .C1(_24299_),
    .Y(_24300_));
 sky130_fd_sc_hd__nand3_2 _27548_ (.A(_24294_),
    .B(_24296_),
    .C(_24300_),
    .Y(_24301_));
 sky130_fd_sc_hd__nand3_1 _27549_ (.A(_24297_),
    .B(_24299_),
    .C(_24293_),
    .Y(_24302_));
 sky130_fd_sc_hd__o2bb2ai_2 _27550_ (.A1_N(_24297_),
    .A2_N(_24299_),
    .B1(_24288_),
    .B2(_24291_),
    .Y(_24304_));
 sky130_fd_sc_hd__o211ai_4 _27551_ (.A1(_23539_),
    .A2(_24295_),
    .B1(_24302_),
    .C1(_24304_),
    .Y(_24305_));
 sky130_fd_sc_hd__nand2_2 _27552_ (.A(_22792_),
    .B(_22788_),
    .Y(_24306_));
 sky130_fd_sc_hd__a21o_1 _27553_ (.A1(_24301_),
    .A2(_24305_),
    .B1(_24306_),
    .X(_24307_));
 sky130_fd_sc_hd__nand3_2 _27554_ (.A(_24301_),
    .B(_24305_),
    .C(_24306_),
    .Y(_24308_));
 sky130_fd_sc_hd__o2bb2a_2 _27555_ (.A1_N(_23305_),
    .A2_N(_22810_),
    .B1(_23544_),
    .B2(_23306_),
    .X(_24309_));
 sky130_fd_sc_hd__or2_1 _27556_ (.A(_23146_),
    .B(_23173_),
    .X(_24310_));
 sky130_fd_sc_hd__inv_2 _27557_ (.A(\delay_line[28][10] ),
    .Y(_24311_));
 sky130_fd_sc_hd__o21ai_1 _27558_ (.A1(_21204_),
    .A2(_23179_),
    .B1(_24311_),
    .Y(_24312_));
 sky130_fd_sc_hd__nand3b_1 _27559_ (.A_N(_21204_),
    .B(\delay_line[28][9] ),
    .C(\delay_line[28][10] ),
    .Y(_24313_));
 sky130_fd_sc_hd__buf_1 _27560_ (.A(_18510_),
    .X(_24315_));
 sky130_fd_sc_hd__a21o_1 _27561_ (.A1(_24312_),
    .A2(_24313_),
    .B1(_24315_),
    .X(_24316_));
 sky130_fd_sc_hd__nand3_1 _27562_ (.A(_24312_),
    .B(_24313_),
    .C(_24315_),
    .Y(_24317_));
 sky130_fd_sc_hd__o21ai_1 _27563_ (.A1(_23177_),
    .A2(_23178_),
    .B1(_23181_),
    .Y(_24318_));
 sky130_fd_sc_hd__o21ai_1 _27564_ (.A1(_18508_),
    .A2(_24318_),
    .B1(_23180_),
    .Y(_24319_));
 sky130_fd_sc_hd__a21oi_1 _27565_ (.A1(_24316_),
    .A2(_24317_),
    .B1(_24319_),
    .Y(_24320_));
 sky130_fd_sc_hd__and3_1 _27566_ (.A(_24319_),
    .B(_24316_),
    .C(_24317_),
    .X(_24321_));
 sky130_fd_sc_hd__or3_1 _27567_ (.A(_20428_),
    .B(_24320_),
    .C(_24321_),
    .X(_24322_));
 sky130_fd_sc_hd__o21ai_1 _27568_ (.A1(_24320_),
    .A2(_24321_),
    .B1(_20428_),
    .Y(_24323_));
 sky130_fd_sc_hd__and3_1 _27569_ (.A(_23176_),
    .B(_23182_),
    .C(_23185_),
    .X(_24324_));
 sky130_fd_sc_hd__a221o_1 _27570_ (.A1(_06425_),
    .A2(_23187_),
    .B1(_24322_),
    .B2(_24323_),
    .C1(_24324_),
    .X(_24326_));
 sky130_fd_sc_hd__o211ai_2 _27571_ (.A1(_24324_),
    .A2(_23189_),
    .B1(_24322_),
    .C1(_24323_),
    .Y(_24327_));
 sky130_fd_sc_hd__nand2_1 _27572_ (.A(_24326_),
    .B(_24327_),
    .Y(_24328_));
 sky130_fd_sc_hd__nor2_1 _27573_ (.A(_23192_),
    .B(_24328_),
    .Y(_24329_));
 sky130_fd_sc_hd__and2_1 _27574_ (.A(_23192_),
    .B(_24328_),
    .X(_24330_));
 sky130_fd_sc_hd__nor2_2 _27575_ (.A(_24329_),
    .B(_24330_),
    .Y(_24331_));
 sky130_fd_sc_hd__or4_1 _27576_ (.A(_21211_),
    .B(_21212_),
    .C(_21214_),
    .D(_23193_),
    .X(_24332_));
 sky130_fd_sc_hd__o21ai_4 _27577_ (.A1(_23195_),
    .A2(_23196_),
    .B1(_24332_),
    .Y(_24333_));
 sky130_fd_sc_hd__xor2_4 _27578_ (.A(_24331_),
    .B(_24333_),
    .X(_24334_));
 sky130_fd_sc_hd__a21bo_1 _27579_ (.A1(_23137_),
    .A2(_23140_),
    .B1_N(_23138_),
    .X(_24335_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27580_ (.A(net337),
    .X(_24337_));
 sky130_fd_sc_hd__buf_1 _27581_ (.A(net338),
    .X(_24338_));
 sky130_fd_sc_hd__o21ai_1 _27582_ (.A1(_18486_),
    .A2(_24338_),
    .B1(_01161_),
    .Y(_24339_));
 sky130_fd_sc_hd__and2_2 _27583_ (.A(_18488_),
    .B(net338),
    .X(_24340_));
 sky130_fd_sc_hd__o21ai_2 _27584_ (.A1(_24347_),
    .A2(_23125_),
    .B1(_23129_),
    .Y(_24341_));
 sky130_fd_sc_hd__nor2_1 _27585_ (.A(_18486_),
    .B(_24338_),
    .Y(_24342_));
 sky130_fd_sc_hd__o21bai_2 _27586_ (.A1(_24340_),
    .A2(_24342_),
    .B1_N(_19266_),
    .Y(_24343_));
 sky130_fd_sc_hd__o211ai_2 _27587_ (.A1(_24339_),
    .A2(_24340_),
    .B1(_24341_),
    .C1(_24343_),
    .Y(_24344_));
 sky130_fd_sc_hd__a21o_1 _27588_ (.A1(_19271_),
    .A2(_24338_),
    .B1(_24339_),
    .X(_24345_));
 sky130_fd_sc_hd__a21o_1 _27589_ (.A1(_24345_),
    .A2(_24343_),
    .B1(_24341_),
    .X(_24346_));
 sky130_fd_sc_hd__o2111ai_2 _27590_ (.A1(_23134_),
    .A2(_23135_),
    .B1(_23132_),
    .C1(_24344_),
    .D1(_24346_),
    .Y(_24348_));
 sky130_fd_sc_hd__o211a_1 _27591_ (.A1(_18487_),
    .A2(_18490_),
    .B1(_16031_),
    .C1(_06590_),
    .X(_24349_));
 sky130_fd_sc_hd__and3_2 _27592_ (.A(_24341_),
    .B(_24345_),
    .C(_24343_),
    .X(_24350_));
 sky130_fd_sc_hd__a21oi_2 _27593_ (.A1(_24345_),
    .A2(_24343_),
    .B1(_24341_),
    .Y(_24351_));
 sky130_fd_sc_hd__o22ai_1 _27594_ (.A1(_24349_),
    .A2(_23136_),
    .B1(_24350_),
    .B2(_24351_),
    .Y(_24352_));
 sky130_fd_sc_hd__nand3b_1 _27595_ (.A_N(_24337_),
    .B(_24348_),
    .C(_24352_),
    .Y(_24353_));
 sky130_fd_sc_hd__a21bo_1 _27596_ (.A1(_24348_),
    .A2(_24352_),
    .B1_N(_24337_),
    .X(_24354_));
 sky130_fd_sc_hd__nand2_1 _27597_ (.A(_24353_),
    .B(_24354_),
    .Y(_24355_));
 sky130_fd_sc_hd__xnor2_1 _27598_ (.A(_24335_),
    .B(_24355_),
    .Y(_24356_));
 sky130_fd_sc_hd__xor2_1 _27599_ (.A(_23145_),
    .B(_24356_),
    .X(_24357_));
 sky130_fd_sc_hd__nor2_1 _27600_ (.A(\delay_line[27][8] ),
    .B(\delay_line[27][10] ),
    .Y(_24359_));
 sky130_fd_sc_hd__buf_1 _27601_ (.A(\delay_line[27][10] ),
    .X(_24360_));
 sky130_fd_sc_hd__nand2_1 _27602_ (.A(_21235_),
    .B(_24360_),
    .Y(_24361_));
 sky130_fd_sc_hd__nand3b_2 _27603_ (.A_N(_24359_),
    .B(_24361_),
    .C(_23155_),
    .Y(_24362_));
 sky130_fd_sc_hd__and2_1 _27604_ (.A(_21235_),
    .B(_24360_),
    .X(_24363_));
 sky130_fd_sc_hd__o21ai_1 _27605_ (.A1(_24359_),
    .A2(_24363_),
    .B1(_23153_),
    .Y(_24364_));
 sky130_fd_sc_hd__nand2_1 _27606_ (.A(_24362_),
    .B(_24364_),
    .Y(_24365_));
 sky130_fd_sc_hd__clkbuf_2 _27607_ (.A(_24360_),
    .X(_24366_));
 sky130_fd_sc_hd__nor2_1 _27608_ (.A(_24366_),
    .B(_23154_),
    .Y(_24367_));
 sky130_fd_sc_hd__a21oi_1 _27609_ (.A1(_23162_),
    .A2(_24365_),
    .B1(_24367_),
    .Y(_24368_));
 sky130_fd_sc_hd__nand3_2 _27610_ (.A(_24368_),
    .B(_16119_),
    .C(_16097_),
    .Y(_24370_));
 sky130_fd_sc_hd__a21o_1 _27611_ (.A1(_16097_),
    .A2(_16119_),
    .B1(_24368_),
    .X(_24371_));
 sky130_fd_sc_hd__o21ai_1 _27612_ (.A1(_23158_),
    .A2(_23151_),
    .B1(_23160_),
    .Y(_24372_));
 sky130_fd_sc_hd__a21o_1 _27613_ (.A1(_24370_),
    .A2(_24371_),
    .B1(_24372_),
    .X(_24373_));
 sky130_fd_sc_hd__nand3_2 _27614_ (.A(_24372_),
    .B(_24370_),
    .C(_24371_),
    .Y(_24374_));
 sky130_fd_sc_hd__nand3_2 _27615_ (.A(_24373_),
    .B(_24374_),
    .C(_06524_),
    .Y(_24375_));
 sky130_fd_sc_hd__a21o_1 _27616_ (.A1(_24373_),
    .A2(_24374_),
    .B1(_06524_),
    .X(_24376_));
 sky130_fd_sc_hd__nand2_2 _27617_ (.A(_24375_),
    .B(_24376_),
    .Y(_24377_));
 sky130_fd_sc_hd__o21ai_1 _27618_ (.A1(_23168_),
    .A2(_23167_),
    .B1(_23165_),
    .Y(_24378_));
 sky130_fd_sc_hd__xnor2_2 _27619_ (.A(_24377_),
    .B(_24378_),
    .Y(_24379_));
 sky130_fd_sc_hd__or3_1 _27620_ (.A(_21245_),
    .B(_21246_),
    .C(_20389_),
    .X(_24381_));
 sky130_fd_sc_hd__a2bb2o_1 _27621_ (.A1_N(_23167_),
    .A2_N(_24381_),
    .B1(_23170_),
    .B2(_23171_),
    .X(_24382_));
 sky130_fd_sc_hd__xnor2_2 _27622_ (.A(_24379_),
    .B(_24382_),
    .Y(_24383_));
 sky130_fd_sc_hd__or2_1 _27623_ (.A(_24357_),
    .B(_24383_),
    .X(_24384_));
 sky130_fd_sc_hd__nand2_1 _27624_ (.A(_24357_),
    .B(_24383_),
    .Y(_24385_));
 sky130_fd_sc_hd__and2_1 _27625_ (.A(_24384_),
    .B(_24385_),
    .X(_24386_));
 sky130_fd_sc_hd__nand2_1 _27626_ (.A(_24334_),
    .B(_24386_),
    .Y(_24387_));
 sky130_fd_sc_hd__or2_1 _27627_ (.A(_24334_),
    .B(_24386_),
    .X(_24388_));
 sky130_fd_sc_hd__nand2_1 _27628_ (.A(_24387_),
    .B(_24388_),
    .Y(_24389_));
 sky130_fd_sc_hd__and3_1 _27629_ (.A(_24310_),
    .B(_23199_),
    .C(_24389_),
    .X(_24390_));
 sky130_fd_sc_hd__a21oi_1 _27630_ (.A1(_24310_),
    .A2(_23199_),
    .B1(_24389_),
    .Y(_24392_));
 sky130_fd_sc_hd__o211ai_2 _27631_ (.A1(_23284_),
    .A2(_21337_),
    .B1(_21340_),
    .C1(_23281_),
    .Y(_24393_));
 sky130_fd_sc_hd__nand2_2 _27632_ (.A(_21310_),
    .B(\delay_line[30][7] ),
    .Y(_24394_));
 sky130_fd_sc_hd__nand2_2 _27633_ (.A(_20339_),
    .B(\delay_line[30][5] ),
    .Y(_24395_));
 sky130_fd_sc_hd__a21boi_4 _27634_ (.A1(_24394_),
    .A2(_24395_),
    .B1_N(\delay_line[30][10] ),
    .Y(_24396_));
 sky130_fd_sc_hd__and3b_2 _27635_ (.A_N(\delay_line[30][10] ),
    .B(_24394_),
    .C(_24395_),
    .X(_24397_));
 sky130_fd_sc_hd__nor2_1 _27636_ (.A(_24396_),
    .B(_24397_),
    .Y(_24398_));
 sky130_fd_sc_hd__a31o_1 _27637_ (.A1(_23247_),
    .A2(_23251_),
    .A3(_23252_),
    .B1(_23256_),
    .X(_24399_));
 sky130_fd_sc_hd__nand2_1 _27638_ (.A(_24398_),
    .B(_24399_),
    .Y(_24400_));
 sky130_fd_sc_hd__o211ai_4 _27639_ (.A1(_24396_),
    .A2(_24397_),
    .B1(_23250_),
    .C1(_23254_),
    .Y(_24401_));
 sky130_fd_sc_hd__and3_1 _27640_ (.A(_01007_),
    .B(_20340_),
    .C(_19335_),
    .X(_24403_));
 sky130_fd_sc_hd__a211o_1 _27641_ (.A1(_21313_),
    .A2(_23251_),
    .B1(_24403_),
    .C1(_19329_),
    .X(_24404_));
 sky130_fd_sc_hd__a21oi_1 _27642_ (.A1(_20341_),
    .A2(_20344_),
    .B1(_23257_),
    .Y(_24405_));
 sky130_fd_sc_hd__o21ai_2 _27643_ (.A1(_24405_),
    .A2(_24403_),
    .B1(_19329_),
    .Y(_24406_));
 sky130_fd_sc_hd__nand2_1 _27644_ (.A(_24404_),
    .B(_24406_),
    .Y(_24407_));
 sky130_fd_sc_hd__a21o_1 _27645_ (.A1(_24400_),
    .A2(_24401_),
    .B1(_24407_),
    .X(_24408_));
 sky130_fd_sc_hd__nand3_1 _27646_ (.A(_24407_),
    .B(_24400_),
    .C(_24401_),
    .Y(_24409_));
 sky130_fd_sc_hd__nand4_1 _27647_ (.A(_23265_),
    .B(_23266_),
    .C(_24408_),
    .D(_24409_),
    .Y(_24410_));
 sky130_fd_sc_hd__a21o_1 _27648_ (.A1(_23261_),
    .A2(_23264_),
    .B1(_23267_),
    .X(_24411_));
 sky130_fd_sc_hd__nand4_1 _27649_ (.A(_24404_),
    .B(_24406_),
    .C(_24400_),
    .D(_24401_),
    .Y(_24412_));
 sky130_fd_sc_hd__a22o_1 _27650_ (.A1(_24404_),
    .A2(_24406_),
    .B1(_24400_),
    .B2(_24401_),
    .X(_24414_));
 sky130_fd_sc_hd__nand3_2 _27651_ (.A(_24411_),
    .B(_24412_),
    .C(_24414_),
    .Y(_24415_));
 sky130_fd_sc_hd__a21o_1 _27652_ (.A1(_24410_),
    .A2(_24415_),
    .B1(_23263_),
    .X(_24416_));
 sky130_fd_sc_hd__nand3_2 _27653_ (.A(_24415_),
    .B(_23263_),
    .C(_24410_),
    .Y(_24417_));
 sky130_fd_sc_hd__nand2_1 _27654_ (.A(_24416_),
    .B(_24417_),
    .Y(_24418_));
 sky130_fd_sc_hd__nor2_1 _27655_ (.A(_23273_),
    .B(_23276_),
    .Y(_24419_));
 sky130_fd_sc_hd__nand2_1 _27656_ (.A(_24418_),
    .B(_24419_),
    .Y(_24420_));
 sky130_fd_sc_hd__o211ai_4 _27657_ (.A1(_23273_),
    .A2(_23276_),
    .B1(_24416_),
    .C1(_24417_),
    .Y(_24421_));
 sky130_fd_sc_hd__nand4_2 _27658_ (.A(_23242_),
    .B(_24420_),
    .C(_23278_),
    .D(_24421_),
    .Y(_24422_));
 sky130_fd_sc_hd__inv_2 _27659_ (.A(_24422_),
    .Y(_24423_));
 sky130_fd_sc_hd__a22oi_1 _27660_ (.A1(_23278_),
    .A2(_23242_),
    .B1(_24420_),
    .B2(_24421_),
    .Y(_24425_));
 sky130_fd_sc_hd__nor2_1 _27661_ (.A(_24423_),
    .B(_24425_),
    .Y(_24426_));
 sky130_fd_sc_hd__a21o_1 _27662_ (.A1(_23280_),
    .A2(_24393_),
    .B1(_24426_),
    .X(_24427_));
 sky130_fd_sc_hd__nand3_1 _27663_ (.A(_23280_),
    .B(_24393_),
    .C(_24426_),
    .Y(_24428_));
 sky130_fd_sc_hd__and2_1 _27664_ (.A(_24427_),
    .B(_24428_),
    .X(_24429_));
 sky130_fd_sc_hd__or3b_1 _27665_ (.A(_23235_),
    .B(_15646_),
    .C_N(_21300_),
    .X(_24430_));
 sky130_fd_sc_hd__and2b_1 _27666_ (.A_N(_19322_),
    .B(net322),
    .X(_24431_));
 sky130_fd_sc_hd__and2b_1 _27667_ (.A_N(net322),
    .B(_19323_),
    .X(_24432_));
 sky130_fd_sc_hd__nor2_1 _27668_ (.A(_24431_),
    .B(_24432_),
    .Y(_24433_));
 sky130_fd_sc_hd__and3_1 _27669_ (.A(_23233_),
    .B(_24430_),
    .C(_24433_),
    .X(_24434_));
 sky130_fd_sc_hd__a21oi_1 _27670_ (.A1(_23233_),
    .A2(_24430_),
    .B1(_24433_),
    .Y(_24436_));
 sky130_fd_sc_hd__a31o_1 _27671_ (.A1(_21303_),
    .A2(_23233_),
    .A3(_23234_),
    .B1(_23240_),
    .X(_24437_));
 sky130_fd_sc_hd__o21ai_2 _27672_ (.A1(_24434_),
    .A2(_24436_),
    .B1(_24437_),
    .Y(_24438_));
 sky130_fd_sc_hd__or3_2 _27673_ (.A(_24434_),
    .B(_24436_),
    .C(_24437_),
    .X(_24439_));
 sky130_fd_sc_hd__nand3_4 _27674_ (.A(_24429_),
    .B(_24438_),
    .C(_24439_),
    .Y(_24440_));
 sky130_fd_sc_hd__a21o_1 _27675_ (.A1(_24439_),
    .A2(_24438_),
    .B1(_24429_),
    .X(_24441_));
 sky130_fd_sc_hd__nand2_1 _27676_ (.A(_24440_),
    .B(_24441_),
    .Y(_24442_));
 sky130_fd_sc_hd__inv_2 _27677_ (.A(_23211_),
    .Y(_24443_));
 sky130_fd_sc_hd__o21ai_1 _27678_ (.A1(_23217_),
    .A2(_24443_),
    .B1(_23215_),
    .Y(_24444_));
 sky130_fd_sc_hd__nor2_1 _27679_ (.A(_00952_),
    .B(_19356_),
    .Y(_24445_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27680_ (.A(_19356_),
    .X(_24447_));
 sky130_fd_sc_hd__nand2_1 _27681_ (.A(_24447_),
    .B(_00952_),
    .Y(_24448_));
 sky130_fd_sc_hd__or4b_2 _27682_ (.A(_24578_),
    .B(_06260_),
    .C(_24445_),
    .D_N(_24448_),
    .X(_24449_));
 sky130_fd_sc_hd__nand2_1 _27683_ (.A(_15712_),
    .B(_15789_),
    .Y(_24450_));
 sky130_fd_sc_hd__a2bb2o_1 _27684_ (.A1_N(_20317_),
    .A2_N(_06260_),
    .B1(_24450_),
    .B2(_24448_),
    .X(_24451_));
 sky130_fd_sc_hd__nand2_1 _27685_ (.A(_24449_),
    .B(_24451_),
    .Y(_24452_));
 sky130_fd_sc_hd__buf_1 _27686_ (.A(\delay_line[31][10] ),
    .X(_24453_));
 sky130_fd_sc_hd__nor2_1 _27687_ (.A(_23206_),
    .B(_24453_),
    .Y(_24454_));
 sky130_fd_sc_hd__nand2_1 _27688_ (.A(_23213_),
    .B(_24453_),
    .Y(_24455_));
 sky130_fd_sc_hd__nand3b_1 _27689_ (.A_N(_24454_),
    .B(_24455_),
    .C(_21264_),
    .Y(_24456_));
 sky130_fd_sc_hd__and2_1 _27690_ (.A(_23206_),
    .B(_24453_),
    .X(_24458_));
 sky130_fd_sc_hd__o21ai_1 _27691_ (.A1(_24454_),
    .A2(_24458_),
    .B1(_21262_),
    .Y(_24459_));
 sky130_fd_sc_hd__o21ai_1 _27692_ (.A1(_20308_),
    .A2(_23208_),
    .B1(_23209_),
    .Y(_24460_));
 sky130_fd_sc_hd__a21o_1 _27693_ (.A1(_24456_),
    .A2(_24459_),
    .B1(_24460_),
    .X(_24461_));
 sky130_fd_sc_hd__and3_1 _27694_ (.A(_21263_),
    .B(_23210_),
    .C(_23214_),
    .X(_24462_));
 sky130_fd_sc_hd__nand3_1 _27695_ (.A(_24460_),
    .B(_24456_),
    .C(_24459_),
    .Y(_24463_));
 sky130_fd_sc_hd__and3_1 _27696_ (.A(_24461_),
    .B(_24462_),
    .C(_24463_),
    .X(_24464_));
 sky130_fd_sc_hd__a32o_1 _27697_ (.A1(_21263_),
    .A2(_23210_),
    .A3(_23214_),
    .B1(_24463_),
    .B2(_24461_),
    .X(_24465_));
 sky130_fd_sc_hd__nor3b_1 _27698_ (.A(_24452_),
    .B(_24464_),
    .C_N(_24465_),
    .Y(_24466_));
 sky130_fd_sc_hd__nand3_1 _27699_ (.A(_24461_),
    .B(_24462_),
    .C(_24463_),
    .Y(_24467_));
 sky130_fd_sc_hd__a22oi_1 _27700_ (.A1(_24449_),
    .A2(_24451_),
    .B1(_24467_),
    .B2(_24465_),
    .Y(_24469_));
 sky130_fd_sc_hd__nor2_1 _27701_ (.A(_24466_),
    .B(_24469_),
    .Y(_24470_));
 sky130_fd_sc_hd__or2_1 _27702_ (.A(_24444_),
    .B(_24470_),
    .X(_24471_));
 sky130_fd_sc_hd__nand2_1 _27703_ (.A(_24470_),
    .B(_24444_),
    .Y(_24472_));
 sky130_fd_sc_hd__nand2_2 _27704_ (.A(_24471_),
    .B(_24472_),
    .Y(_24473_));
 sky130_fd_sc_hd__o21ai_1 _27705_ (.A1(_21283_),
    .A2(_23223_),
    .B1(_23221_),
    .Y(_24474_));
 sky130_fd_sc_hd__xnor2_1 _27706_ (.A(_24473_),
    .B(_24474_),
    .Y(_24475_));
 sky130_fd_sc_hd__nand2_1 _27707_ (.A(_23228_),
    .B(_24475_),
    .Y(_24476_));
 sky130_fd_sc_hd__a21o_1 _27708_ (.A1(_20329_),
    .A2(_19376_),
    .B1(_21260_),
    .X(_24477_));
 sky130_fd_sc_hd__nand2_1 _27709_ (.A(_21294_),
    .B(_23204_),
    .Y(_24478_));
 sky130_fd_sc_hd__o21ai_1 _27710_ (.A1(_21289_),
    .A2(_24478_),
    .B1(_23226_),
    .Y(_24480_));
 sky130_fd_sc_hd__a21oi_2 _27711_ (.A1(_24477_),
    .A2(_21295_),
    .B1(_24480_),
    .Y(_24481_));
 sky130_fd_sc_hd__nor2_1 _27712_ (.A(_24475_),
    .B(_23230_),
    .Y(_24482_));
 sky130_fd_sc_hd__a2bb2o_1 _27713_ (.A1_N(_24476_),
    .A2_N(_24481_),
    .B1(_23226_),
    .B2(_24482_),
    .X(_24483_));
 sky130_fd_sc_hd__xnor2_1 _27714_ (.A(_24442_),
    .B(_24483_),
    .Y(_24484_));
 sky130_fd_sc_hd__o21a_1 _27715_ (.A1(_24390_),
    .A2(_24392_),
    .B1(_24484_),
    .X(_24485_));
 sky130_fd_sc_hd__nor3_1 _27716_ (.A(_24390_),
    .B(_24392_),
    .C(_24484_),
    .Y(_24486_));
 sky130_fd_sc_hd__nor2_2 _27717_ (.A(_24485_),
    .B(_24486_),
    .Y(_24487_));
 sky130_fd_sc_hd__o21a_1 _27718_ (.A1(_22917_),
    .A2(_22920_),
    .B1(_24487_),
    .X(_24488_));
 sky130_fd_sc_hd__or3_1 _27719_ (.A(_22917_),
    .B(_22920_),
    .C(_24487_),
    .X(_24489_));
 sky130_fd_sc_hd__and2b_1 _27720_ (.A_N(_24488_),
    .B(_24489_),
    .X(_24491_));
 sky130_fd_sc_hd__nand2_2 _27721_ (.A(_23203_),
    .B(_23294_),
    .Y(_24492_));
 sky130_fd_sc_hd__xnor2_1 _27722_ (.A(_24491_),
    .B(_24492_),
    .Y(_24493_));
 sky130_fd_sc_hd__a21oi_2 _27723_ (.A1(_21550_),
    .A2(_22923_),
    .B1(_23118_),
    .Y(_24494_));
 sky130_fd_sc_hd__a21o_1 _27724_ (.A1(_22922_),
    .A2(_23119_),
    .B1(_24494_),
    .X(_24495_));
 sky130_fd_sc_hd__nand2_1 _27725_ (.A(_22835_),
    .B(_22840_),
    .Y(_24496_));
 sky130_fd_sc_hd__o21ai_1 _27726_ (.A1(_20501_),
    .A2(_21595_),
    .B1(_22845_),
    .Y(_24497_));
 sky130_fd_sc_hd__a2bb2oi_4 _27727_ (.A1_N(_21592_),
    .A2_N(_24496_),
    .B1(_22847_),
    .B2(_24497_),
    .Y(_24498_));
 sky130_fd_sc_hd__buf_2 _27728_ (.A(_17150_),
    .X(_24499_));
 sky130_fd_sc_hd__a21oi_1 _27729_ (.A1(_06810_),
    .A2(_17150_),
    .B1(_17182_),
    .Y(_24500_));
 sky130_fd_sc_hd__and3_1 _27730_ (.A(_06810_),
    .B(_17226_),
    .C(_06788_),
    .X(_24502_));
 sky130_fd_sc_hd__and2_1 _27731_ (.A(_21562_),
    .B(\delay_line[25][10] ),
    .X(_24503_));
 sky130_fd_sc_hd__clkbuf_2 _27732_ (.A(_24503_),
    .X(_24504_));
 sky130_fd_sc_hd__clkbuf_2 _27733_ (.A(\delay_line[25][10] ),
    .X(_24505_));
 sky130_fd_sc_hd__o211ai_4 _27734_ (.A1(_21562_),
    .A2(_24505_),
    .B1(_22819_),
    .C1(_20483_),
    .Y(_24506_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27735_ (.A(_18324_),
    .X(_24507_));
 sky130_fd_sc_hd__nor2_1 _27736_ (.A(_21563_),
    .B(_24505_),
    .Y(_24508_));
 sky130_fd_sc_hd__o21bai_2 _27737_ (.A1(_24504_),
    .A2(_24508_),
    .B1_N(_22813_),
    .Y(_24509_));
 sky130_fd_sc_hd__o211ai_2 _27738_ (.A1(_24504_),
    .A2(_24506_),
    .B1(_24507_),
    .C1(_24509_),
    .Y(_24510_));
 sky130_fd_sc_hd__buf_1 _27739_ (.A(_24505_),
    .X(_24511_));
 sky130_fd_sc_hd__a21o_1 _27740_ (.A1(_21563_),
    .A2(_24511_),
    .B1(_24506_),
    .X(_24513_));
 sky130_fd_sc_hd__a21o_1 _27741_ (.A1(_24513_),
    .A2(_24509_),
    .B1(_18324_),
    .X(_24514_));
 sky130_fd_sc_hd__o2bb2ai_2 _27742_ (.A1_N(_22822_),
    .A2_N(_22817_),
    .B1(_22815_),
    .B2(_22813_),
    .Y(_24515_));
 sky130_fd_sc_hd__nand3_2 _27743_ (.A(_24510_),
    .B(_24514_),
    .C(_24515_),
    .Y(_24516_));
 sky130_fd_sc_hd__o211a_1 _27744_ (.A1(_24504_),
    .A2(_24506_),
    .B1(_18324_),
    .C1(_24509_),
    .X(_24517_));
 sky130_fd_sc_hd__a21oi_1 _27745_ (.A1(_24513_),
    .A2(_24509_),
    .B1(_24507_),
    .Y(_24518_));
 sky130_fd_sc_hd__o21bai_2 _27746_ (.A1(_24517_),
    .A2(_24518_),
    .B1_N(_24515_),
    .Y(_24519_));
 sky130_fd_sc_hd__o211ai_1 _27747_ (.A1(_24500_),
    .A2(_24502_),
    .B1(_24516_),
    .C1(_24519_),
    .Y(_24520_));
 sky130_fd_sc_hd__a2bb2o_1 _27748_ (.A1_N(_06788_),
    .A2_N(_22836_),
    .B1(_06777_),
    .B2(_17150_),
    .X(_24521_));
 sky130_fd_sc_hd__a21o_1 _27749_ (.A1(_24516_),
    .A2(_24519_),
    .B1(_24521_),
    .X(_24522_));
 sky130_fd_sc_hd__a21boi_1 _27750_ (.A1(_22827_),
    .A2(_22829_),
    .B1_N(_22825_),
    .Y(_24524_));
 sky130_fd_sc_hd__nand3_2 _27751_ (.A(_24520_),
    .B(_24522_),
    .C(_24524_),
    .Y(_24525_));
 sky130_fd_sc_hd__o211a_1 _27752_ (.A1(_24500_),
    .A2(_24502_),
    .B1(_24516_),
    .C1(_24519_),
    .X(_24526_));
 sky130_fd_sc_hd__a21oi_1 _27753_ (.A1(_24516_),
    .A2(_24519_),
    .B1(_24521_),
    .Y(_24527_));
 sky130_fd_sc_hd__o21bai_4 _27754_ (.A1(_24526_),
    .A2(_24527_),
    .B1_N(_24524_),
    .Y(_24528_));
 sky130_fd_sc_hd__o2111ai_4 _27755_ (.A1(_24499_),
    .A2(_21577_),
    .B1(_23742_),
    .C1(_24525_),
    .D1(_24528_),
    .Y(_24529_));
 sky130_fd_sc_hd__nor2_1 _27756_ (.A(_24499_),
    .B(_21577_),
    .Y(_24530_));
 sky130_fd_sc_hd__o2bb2ai_2 _27757_ (.A1_N(_24525_),
    .A2_N(_24528_),
    .B1(_24530_),
    .B2(_06821_),
    .Y(_24531_));
 sky130_fd_sc_hd__a21o_1 _27758_ (.A1(_22834_),
    .A2(_22380_),
    .B1(_22833_),
    .X(_24532_));
 sky130_fd_sc_hd__nand3_1 _27759_ (.A(_24529_),
    .B(_24531_),
    .C(_24532_),
    .Y(_24533_));
 sky130_fd_sc_hd__a21o_1 _27760_ (.A1(_24529_),
    .A2(_24531_),
    .B1(_24532_),
    .X(_24535_));
 sky130_fd_sc_hd__o2bb2ai_1 _27761_ (.A1_N(_24533_),
    .A2_N(_24535_),
    .B1(_21591_),
    .B2(_24496_),
    .Y(_24536_));
 sky130_fd_sc_hd__and3_1 _27762_ (.A(_22835_),
    .B(_22840_),
    .C(_21584_),
    .X(_24537_));
 sky130_fd_sc_hd__nand3_2 _27763_ (.A(_24537_),
    .B(_24533_),
    .C(_24535_),
    .Y(_24538_));
 sky130_fd_sc_hd__nand2_2 _27764_ (.A(_24536_),
    .B(_24538_),
    .Y(_24539_));
 sky130_fd_sc_hd__xnor2_2 _27765_ (.A(_24498_),
    .B(_24539_),
    .Y(_24540_));
 sky130_fd_sc_hd__buf_1 _27766_ (.A(_22863_),
    .X(_24541_));
 sky130_fd_sc_hd__and3_1 _27767_ (.A(_21610_),
    .B(_24541_),
    .C(_22865_),
    .X(_24542_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27768_ (.A(\delay_line[22][9] ),
    .X(_24543_));
 sky130_fd_sc_hd__o21ai_1 _27769_ (.A1(net353),
    .A2(_24543_),
    .B1(_22857_),
    .Y(_24544_));
 sky130_fd_sc_hd__and2_1 _27770_ (.A(net353),
    .B(_24543_),
    .X(_24546_));
 sky130_fd_sc_hd__or2_1 _27771_ (.A(net355),
    .B(_22851_),
    .X(_24547_));
 sky130_fd_sc_hd__nor2_1 _27772_ (.A(net356),
    .B(net355),
    .Y(_24548_));
 sky130_fd_sc_hd__and2_1 _27773_ (.A(net356),
    .B(net355),
    .X(_24549_));
 sky130_fd_sc_hd__o21ai_2 _27774_ (.A1(_24548_),
    .A2(_24549_),
    .B1(_22852_),
    .Y(_24550_));
 sky130_fd_sc_hd__nor2_1 _27775_ (.A(net353),
    .B(_24543_),
    .Y(_24551_));
 sky130_fd_sc_hd__o21ai_2 _27776_ (.A1(_24546_),
    .A2(_24551_),
    .B1(_22855_),
    .Y(_24552_));
 sky130_fd_sc_hd__o2111a_1 _27777_ (.A1(_24544_),
    .A2(_24546_),
    .B1(_24547_),
    .C1(_24550_),
    .D1(_24552_),
    .X(_24553_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27778_ (.A(_24547_),
    .X(_24554_));
 sky130_fd_sc_hd__buf_1 _27779_ (.A(\delay_line[22][9] ),
    .X(_24555_));
 sky130_fd_sc_hd__a21o_1 _27780_ (.A1(_19501_),
    .A2(_24555_),
    .B1(_24544_),
    .X(_24557_));
 sky130_fd_sc_hd__a22oi_2 _27781_ (.A1(_24550_),
    .A2(_24554_),
    .B1(_24557_),
    .B2(_24552_),
    .Y(_24558_));
 sky130_fd_sc_hd__a211o_1 _27782_ (.A1(_22856_),
    .A2(_22861_),
    .B1(_24553_),
    .C1(_24558_),
    .X(_24559_));
 sky130_fd_sc_hd__o211ai_1 _27783_ (.A1(_24553_),
    .A2(_24558_),
    .B1(_22856_),
    .C1(_22861_),
    .Y(_24560_));
 sky130_fd_sc_hd__nand3_1 _27784_ (.A(_24559_),
    .B(_23676_),
    .C(_24560_),
    .Y(_24561_));
 sky130_fd_sc_hd__a21o_1 _27785_ (.A1(_24560_),
    .A2(_24559_),
    .B1(_23666_),
    .X(_24562_));
 sky130_fd_sc_hd__o2111ai_1 _27786_ (.A1(_21607_),
    .A2(_22866_),
    .B1(_24561_),
    .C1(_24562_),
    .D1(_24541_),
    .Y(_24563_));
 sky130_fd_sc_hd__and3_1 _27787_ (.A(_22859_),
    .B(_22861_),
    .C(_22862_),
    .X(_24564_));
 sky130_fd_sc_hd__and3_1 _27788_ (.A(_22865_),
    .B(_22849_),
    .C(_22863_),
    .X(_24565_));
 sky130_fd_sc_hd__nand2_1 _27789_ (.A(_24561_),
    .B(_24562_),
    .Y(_24566_));
 sky130_fd_sc_hd__o21ai_1 _27790_ (.A1(_24564_),
    .A2(_24565_),
    .B1(_24566_),
    .Y(_24568_));
 sky130_fd_sc_hd__nand2_1 _27791_ (.A(_24563_),
    .B(_24568_),
    .Y(_24569_));
 sky130_fd_sc_hd__xor2_1 _27792_ (.A(_24542_),
    .B(_24569_),
    .X(_24570_));
 sky130_fd_sc_hd__a21bo_1 _27793_ (.A1(_22893_),
    .A2(_22894_),
    .B1_N(_22889_),
    .X(_24571_));
 sky130_fd_sc_hd__clkbuf_2 _27794_ (.A(_22887_),
    .X(_24572_));
 sky130_fd_sc_hd__o21ai_1 _27795_ (.A1(_17018_),
    .A2(_22880_),
    .B1(_24572_),
    .Y(_24573_));
 sky130_fd_sc_hd__nor2_1 _27796_ (.A(_19512_),
    .B(\delay_line[24][6] ),
    .Y(_24574_));
 sky130_fd_sc_hd__and2_1 _27797_ (.A(\delay_line[24][5] ),
    .B(\delay_line[24][6] ),
    .X(_24575_));
 sky130_fd_sc_hd__nor3_1 _27798_ (.A(_22874_),
    .B(_24574_),
    .C(_24575_),
    .Y(_24576_));
 sky130_fd_sc_hd__o21ai_1 _27799_ (.A1(_24574_),
    .A2(_24575_),
    .B1(_22874_),
    .Y(_24577_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27800_ (.A(\delay_line[24][9] ),
    .X(_24579_));
 sky130_fd_sc_hd__nand3b_1 _27801_ (.A_N(_24576_),
    .B(_24577_),
    .C(_24579_),
    .Y(_24580_));
 sky130_fd_sc_hd__buf_1 _27802_ (.A(_24580_),
    .X(_24581_));
 sky130_fd_sc_hd__o21a_1 _27803_ (.A1(_24574_),
    .A2(_24575_),
    .B1(_22876_),
    .X(_24582_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27804_ (.A(_24579_),
    .X(_24583_));
 sky130_fd_sc_hd__o21bai_2 _27805_ (.A1(_24576_),
    .A2(_24582_),
    .B1_N(_24583_),
    .Y(_24584_));
 sky130_fd_sc_hd__a21o_1 _27806_ (.A1(_24581_),
    .A2(_24584_),
    .B1(_22888_),
    .X(_24585_));
 sky130_fd_sc_hd__buf_1 _27807_ (.A(_24580_),
    .X(_24586_));
 sky130_fd_sc_hd__nand3_1 _27808_ (.A(_22888_),
    .B(_24586_),
    .C(_24584_),
    .Y(_24587_));
 sky130_fd_sc_hd__nand3_1 _27809_ (.A(_24573_),
    .B(_24585_),
    .C(_24587_),
    .Y(_24588_));
 sky130_fd_sc_hd__nand3_1 _27810_ (.A(_22890_),
    .B(_24586_),
    .C(_24584_),
    .Y(_24590_));
 sky130_fd_sc_hd__a21o_1 _27811_ (.A1(_24581_),
    .A2(_24584_),
    .B1(_22890_),
    .X(_24591_));
 sky130_fd_sc_hd__o2111ai_2 _27812_ (.A1(_17018_),
    .A2(_22880_),
    .B1(_24572_),
    .C1(_24590_),
    .D1(_24591_),
    .Y(_24592_));
 sky130_fd_sc_hd__and3_1 _27813_ (.A(_24571_),
    .B(_24588_),
    .C(_24592_),
    .X(_24593_));
 sky130_fd_sc_hd__a21oi_1 _27814_ (.A1(_24588_),
    .A2(_24592_),
    .B1(_24571_),
    .Y(_24594_));
 sky130_fd_sc_hd__and2_1 _27815_ (.A(_18305_),
    .B(_21618_),
    .X(_24595_));
 sky130_fd_sc_hd__o211a_1 _27816_ (.A1(_17029_),
    .A2(_18310_),
    .B1(_06909_),
    .C1(_23687_),
    .X(_24596_));
 sky130_fd_sc_hd__or2_1 _27817_ (.A(_24595_),
    .B(_24596_),
    .X(_24597_));
 sky130_fd_sc_hd__o21ai_1 _27818_ (.A1(_24593_),
    .A2(_24594_),
    .B1(_24597_),
    .Y(_24598_));
 sky130_fd_sc_hd__inv_2 _27819_ (.A(_24598_),
    .Y(_24599_));
 sky130_fd_sc_hd__nand2_1 _27820_ (.A(_22898_),
    .B(_22904_),
    .Y(_24601_));
 sky130_fd_sc_hd__or4_1 _27821_ (.A(_24595_),
    .B(_24596_),
    .C(_24593_),
    .D(_24594_),
    .X(_24602_));
 sky130_fd_sc_hd__nand2_1 _27822_ (.A(_24601_),
    .B(_24602_),
    .Y(_24603_));
 sky130_fd_sc_hd__a21oi_1 _27823_ (.A1(_24602_),
    .A2(_24598_),
    .B1(_24601_),
    .Y(_24604_));
 sky130_fd_sc_hd__o21bai_1 _27824_ (.A1(_24599_),
    .A2(_24603_),
    .B1_N(_24604_),
    .Y(_24605_));
 sky130_fd_sc_hd__nand2_1 _27825_ (.A(_19523_),
    .B(_20475_),
    .Y(_24606_));
 sky130_fd_sc_hd__o21ai_1 _27826_ (.A1(_24606_),
    .A2(_21644_),
    .B1(_22869_),
    .Y(_24607_));
 sky130_fd_sc_hd__a21boi_2 _27827_ (.A1(_22905_),
    .A2(_24607_),
    .B1_N(_22907_),
    .Y(_24608_));
 sky130_fd_sc_hd__xnor2_1 _27828_ (.A(_24605_),
    .B(_24608_),
    .Y(_24609_));
 sky130_fd_sc_hd__inv_2 _27829_ (.A(_24609_),
    .Y(_24610_));
 sky130_fd_sc_hd__nand2_1 _27830_ (.A(_24570_),
    .B(_24610_),
    .Y(_24612_));
 sky130_fd_sc_hd__or2_1 _27831_ (.A(_24570_),
    .B(_24610_),
    .X(_24613_));
 sky130_fd_sc_hd__nand2_1 _27832_ (.A(_24612_),
    .B(_24613_),
    .Y(_24614_));
 sky130_fd_sc_hd__xor2_1 _27833_ (.A(_24540_),
    .B(_24614_),
    .X(_24615_));
 sky130_fd_sc_hd__nor3_1 _27834_ (.A(net117),
    .B(_23012_),
    .C(_24615_),
    .Y(_24616_));
 sky130_fd_sc_hd__o21a_1 _27835_ (.A1(net117),
    .A2(_23012_),
    .B1(_24615_),
    .X(_24617_));
 sky130_fd_sc_hd__nor2_1 _27836_ (.A(_24616_),
    .B(_24617_),
    .Y(_24618_));
 sky130_fd_sc_hd__o21a_1 _27837_ (.A1(_22912_),
    .A2(net111),
    .B1(_24618_),
    .X(_24619_));
 sky130_fd_sc_hd__nor3_1 _27838_ (.A(_22912_),
    .B(net111),
    .C(_24618_),
    .Y(_24620_));
 sky130_fd_sc_hd__nor2_1 _27839_ (.A(_24619_),
    .B(_24620_),
    .Y(_24621_));
 sky130_fd_sc_hd__nand2_1 _27840_ (.A(_23014_),
    .B(_23116_),
    .Y(_24623_));
 sky130_fd_sc_hd__a21o_1 _27841_ (.A1(_21422_),
    .A2(_21432_),
    .B1(_23002_),
    .X(_24624_));
 sky130_fd_sc_hd__o21ai_1 _27842_ (.A1(_21435_),
    .A2(_23003_),
    .B1(_24624_),
    .Y(_24625_));
 sky130_fd_sc_hd__a2bb2o_1 _27843_ (.A1_N(_22984_),
    .A2_N(_22988_),
    .B1(_16503_),
    .B2(_22989_),
    .X(_24626_));
 sky130_fd_sc_hd__and2_1 _27844_ (.A(net359),
    .B(\delay_line[21][9] ),
    .X(_24627_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27845_ (.A(\delay_line[21][9] ),
    .X(_24628_));
 sky130_fd_sc_hd__nor2_1 _27846_ (.A(_22984_),
    .B(_24628_),
    .Y(_24629_));
 sky130_fd_sc_hd__nand2_1 _27847_ (.A(_21415_),
    .B(net359),
    .Y(_24630_));
 sky130_fd_sc_hd__o21ai_2 _27848_ (.A1(_24627_),
    .A2(_24629_),
    .B1(_24630_),
    .Y(_24631_));
 sky130_fd_sc_hd__or2_1 _27849_ (.A(_24628_),
    .B(_24630_),
    .X(_24632_));
 sky130_fd_sc_hd__a21o_1 _27850_ (.A1(_24631_),
    .A2(_24632_),
    .B1(_18348_),
    .X(_24634_));
 sky130_fd_sc_hd__clkbuf_2 _27851_ (.A(_24628_),
    .X(_24635_));
 sky130_fd_sc_hd__o211ai_2 _27852_ (.A1(_24635_),
    .A2(_24630_),
    .B1(_18348_),
    .C1(_24631_),
    .Y(_24636_));
 sky130_fd_sc_hd__nand3_2 _27853_ (.A(_24626_),
    .B(_24634_),
    .C(_24636_),
    .Y(_24637_));
 sky130_fd_sc_hd__a21o_1 _27854_ (.A1(_24634_),
    .A2(_24636_),
    .B1(_24626_),
    .X(_24638_));
 sky130_fd_sc_hd__o21ba_1 _27855_ (.A1(_21419_),
    .A2(_01611_),
    .B1_N(_01589_),
    .X(_24639_));
 sky130_fd_sc_hd__xor2_1 _27856_ (.A(_18352_),
    .B(_24639_),
    .X(_24640_));
 sky130_fd_sc_hd__a21bo_1 _27857_ (.A1(_24637_),
    .A2(_24638_),
    .B1_N(_24640_),
    .X(_24641_));
 sky130_fd_sc_hd__nand3b_1 _27858_ (.A_N(_24640_),
    .B(_24637_),
    .C(_24638_),
    .Y(_24642_));
 sky130_fd_sc_hd__nand4_1 _27859_ (.A(_22999_),
    .B(_22998_),
    .C(_24641_),
    .D(_24642_),
    .Y(_24643_));
 sky130_fd_sc_hd__a22o_1 _27860_ (.A1(_22999_),
    .A2(_22998_),
    .B1(_24641_),
    .B2(_24642_),
    .X(_24645_));
 sky130_fd_sc_hd__a21boi_1 _27861_ (.A1(_07569_),
    .A2(_07591_),
    .B1_N(_24006_),
    .Y(_24646_));
 sky130_fd_sc_hd__nand3_1 _27862_ (.A(_24643_),
    .B(_24645_),
    .C(_24646_),
    .Y(_24647_));
 sky130_fd_sc_hd__a21o_1 _27863_ (.A1(_24643_),
    .A2(_24645_),
    .B1(_24646_),
    .X(_24648_));
 sky130_fd_sc_hd__nand2_1 _27864_ (.A(_24647_),
    .B(_24648_),
    .Y(_24649_));
 sky130_fd_sc_hd__xnor2_2 _27865_ (.A(_24625_),
    .B(_24649_),
    .Y(_24650_));
 sky130_fd_sc_hd__o22ai_4 _27866_ (.A1(_21436_),
    .A2(_23003_),
    .B1(_23006_),
    .B2(_23008_),
    .Y(_24651_));
 sky130_fd_sc_hd__xnor2_2 _27867_ (.A(_24650_),
    .B(_24651_),
    .Y(_24652_));
 sky130_fd_sc_hd__a21bo_1 _27868_ (.A1(_22951_),
    .A2(_22956_),
    .B1_N(_22955_),
    .X(_24653_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27869_ (.A(\delay_line[19][9] ),
    .X(_24654_));
 sky130_fd_sc_hd__and2_1 _27870_ (.A(\delay_line[19][8] ),
    .B(_24654_),
    .X(_24656_));
 sky130_fd_sc_hd__nor2_1 _27871_ (.A(_22948_),
    .B(_24654_),
    .Y(_24657_));
 sky130_fd_sc_hd__nand2_1 _27872_ (.A(net370),
    .B(_22948_),
    .Y(_24658_));
 sky130_fd_sc_hd__o21ai_2 _27873_ (.A1(_24656_),
    .A2(_24657_),
    .B1(_24658_),
    .Y(_24659_));
 sky130_fd_sc_hd__clkbuf_2 _27874_ (.A(\delay_line[19][9] ),
    .X(_24660_));
 sky130_fd_sc_hd__inv_2 _27875_ (.A(_24660_),
    .Y(_24661_));
 sky130_fd_sc_hd__nand2_1 _27876_ (.A(_22949_),
    .B(_24661_),
    .Y(_24662_));
 sky130_fd_sc_hd__a21o_1 _27877_ (.A1(_24659_),
    .A2(_24662_),
    .B1(_18375_),
    .X(_24663_));
 sky130_fd_sc_hd__o211ai_1 _27878_ (.A1(_24660_),
    .A2(_24658_),
    .B1(_18375_),
    .C1(_24659_),
    .Y(_24664_));
 sky130_fd_sc_hd__nand3_2 _27879_ (.A(_24653_),
    .B(_24663_),
    .C(_24664_),
    .Y(_24665_));
 sky130_fd_sc_hd__a21oi_1 _27880_ (.A1(_24659_),
    .A2(_24662_),
    .B1(_18376_),
    .Y(_24667_));
 sky130_fd_sc_hd__and3_1 _27881_ (.A(_24659_),
    .B(_24662_),
    .C(_18375_),
    .X(_24668_));
 sky130_fd_sc_hd__o21bai_4 _27882_ (.A1(_24667_),
    .A2(_24668_),
    .B1_N(_24653_),
    .Y(_24669_));
 sky130_fd_sc_hd__o21bai_2 _27883_ (.A1(_07393_),
    .A2(_01655_),
    .B1_N(_01633_),
    .Y(_24670_));
 sky130_fd_sc_hd__xnor2_2 _27884_ (.A(_18368_),
    .B(_24670_),
    .Y(_24671_));
 sky130_fd_sc_hd__a21bo_1 _27885_ (.A1(_24665_),
    .A2(_24669_),
    .B1_N(_24671_),
    .X(_24672_));
 sky130_fd_sc_hd__nand3b_1 _27886_ (.A_N(_24671_),
    .B(_24665_),
    .C(_24669_),
    .Y(_24673_));
 sky130_fd_sc_hd__o21a_1 _27887_ (.A1(_23885_),
    .A2(_07404_),
    .B1(_22964_),
    .X(_24674_));
 sky130_fd_sc_hd__a21boi_1 _27888_ (.A1(_22962_),
    .A2(_24674_),
    .B1_N(_22959_),
    .Y(_24675_));
 sky130_fd_sc_hd__nand3_1 _27889_ (.A(_24672_),
    .B(_24673_),
    .C(_24675_),
    .Y(_24676_));
 sky130_fd_sc_hd__nand3_1 _27890_ (.A(_24669_),
    .B(_24671_),
    .C(_24665_),
    .Y(_24678_));
 sky130_fd_sc_hd__a21o_1 _27891_ (.A1(_24665_),
    .A2(_24669_),
    .B1(_24671_),
    .X(_24679_));
 sky130_fd_sc_hd__nand3b_4 _27892_ (.A_N(_24675_),
    .B(_24678_),
    .C(_24679_),
    .Y(_24680_));
 sky130_fd_sc_hd__o2111ai_4 _27893_ (.A1(_01644_),
    .A2(_16371_),
    .B1(_23907_),
    .C1(_24676_),
    .D1(_24680_),
    .Y(_24681_));
 sky130_fd_sc_hd__a2bb2o_1 _27894_ (.A1_N(_23962_),
    .A2_N(_07481_),
    .B1(_24676_),
    .B2(_24680_),
    .X(_24682_));
 sky130_fd_sc_hd__nand2_2 _27895_ (.A(_24681_),
    .B(_24682_),
    .Y(_24683_));
 sky130_fd_sc_hd__o21ai_1 _27896_ (.A1(_21396_),
    .A2(_22976_),
    .B1(_22969_),
    .Y(_24684_));
 sky130_fd_sc_hd__xor2_2 _27897_ (.A(_24683_),
    .B(_24684_),
    .X(_24685_));
 sky130_fd_sc_hd__o31a_1 _27898_ (.A1(_21397_),
    .A2(_22976_),
    .A3(_22975_),
    .B1(_24685_),
    .X(_24686_));
 sky130_fd_sc_hd__inv_2 _27899_ (.A(_22979_),
    .Y(_24687_));
 sky130_fd_sc_hd__nand2_1 _27900_ (.A(_21371_),
    .B(_22938_),
    .Y(_24689_));
 sky130_fd_sc_hd__a22o_1 _27901_ (.A1(_21365_),
    .A2(_21367_),
    .B1(_22934_),
    .B2(_22935_),
    .X(_24690_));
 sky130_fd_sc_hd__a21oi_1 _27902_ (.A1(_23929_),
    .A2(net375),
    .B1(_21355_),
    .Y(_24691_));
 sky130_fd_sc_hd__nor3_1 _27903_ (.A(\delay_line[18][0] ),
    .B(net374),
    .C(_19393_),
    .Y(_24692_));
 sky130_fd_sc_hd__nor2_1 _27904_ (.A(_19390_),
    .B(\delay_line[18][9] ),
    .Y(_24693_));
 sky130_fd_sc_hd__clkbuf_2 _27905_ (.A(\delay_line[18][9] ),
    .X(_24694_));
 sky130_fd_sc_hd__nand2_1 _27906_ (.A(_19390_),
    .B(_24694_),
    .Y(_24695_));
 sky130_fd_sc_hd__nand3b_2 _27907_ (.A_N(_24693_),
    .B(_22927_),
    .C(_24695_),
    .Y(_24696_));
 sky130_fd_sc_hd__and2_1 _27908_ (.A(\delay_line[18][5] ),
    .B(\delay_line[18][9] ),
    .X(_24697_));
 sky130_fd_sc_hd__o21ai_2 _27909_ (.A1(_24697_),
    .A2(_24693_),
    .B1(_22932_),
    .Y(_24698_));
 sky130_fd_sc_hd__o211ai_2 _27910_ (.A1(_24691_),
    .A2(_24692_),
    .B1(_24696_),
    .C1(_24698_),
    .Y(_24700_));
 sky130_fd_sc_hd__a21oi_1 _27911_ (.A1(_23940_),
    .A2(_01666_),
    .B1(_07514_),
    .Y(_24701_));
 sky130_fd_sc_hd__and3_1 _27912_ (.A(_23940_),
    .B(_01666_),
    .C(net374),
    .X(_24702_));
 sky130_fd_sc_hd__o2bb2ai_1 _27913_ (.A1_N(_24696_),
    .A2_N(_24698_),
    .B1(_24701_),
    .B2(_24702_),
    .Y(_24703_));
 sky130_fd_sc_hd__buf_1 _27914_ (.A(_21357_),
    .X(_24704_));
 sky130_fd_sc_hd__o2bb2a_1 _27915_ (.A1_N(_24704_),
    .A2_N(_21363_),
    .B1(_22926_),
    .B2(_22927_),
    .X(_24705_));
 sky130_fd_sc_hd__o21ai_1 _27916_ (.A1(_22929_),
    .A2(_24705_),
    .B1(_22933_),
    .Y(_24706_));
 sky130_fd_sc_hd__a21oi_1 _27917_ (.A1(_24700_),
    .A2(_24703_),
    .B1(_24706_),
    .Y(_24707_));
 sky130_fd_sc_hd__nand3_1 _27918_ (.A(_24706_),
    .B(_24700_),
    .C(_24703_),
    .Y(_24708_));
 sky130_fd_sc_hd__nand3b_2 _27919_ (.A_N(_24707_),
    .B(_24708_),
    .C(_23863_),
    .Y(_24709_));
 sky130_fd_sc_hd__and3_1 _27920_ (.A(_24706_),
    .B(_24700_),
    .C(_24703_),
    .X(_24711_));
 sky130_fd_sc_hd__o21ai_2 _27921_ (.A1(_24707_),
    .A2(_24711_),
    .B1(_23951_),
    .Y(_24712_));
 sky130_fd_sc_hd__o2111ai_2 _27922_ (.A1(_21370_),
    .A2(_22936_),
    .B1(_24690_),
    .C1(_24709_),
    .D1(_24712_),
    .Y(_24713_));
 sky130_fd_sc_hd__nor3_1 _27923_ (.A(_22937_),
    .B(_21370_),
    .C(_22936_),
    .Y(_24714_));
 sky130_fd_sc_hd__nand2_1 _27924_ (.A(_24709_),
    .B(_24712_),
    .Y(_24715_));
 sky130_fd_sc_hd__o21ai_1 _27925_ (.A1(_22937_),
    .A2(_24714_),
    .B1(_24715_),
    .Y(_24716_));
 sky130_fd_sc_hd__and3_1 _27926_ (.A(_24689_),
    .B(_24713_),
    .C(_24716_),
    .X(_24717_));
 sky130_fd_sc_hd__nand2_1 _27927_ (.A(_22968_),
    .B(_22969_),
    .Y(_24718_));
 sky130_fd_sc_hd__and2_1 _27928_ (.A(_22973_),
    .B(_22977_),
    .X(_24719_));
 sky130_fd_sc_hd__a2bb2oi_1 _27929_ (.A1_N(_21397_),
    .A2_N(_24718_),
    .B1(_24719_),
    .B2(_22978_),
    .Y(_24720_));
 sky130_fd_sc_hd__nor2_1 _27930_ (.A(_24685_),
    .B(_24720_),
    .Y(_24722_));
 sky130_fd_sc_hd__a21oi_2 _27931_ (.A1(_24713_),
    .A2(_24716_),
    .B1(_24689_),
    .Y(_24723_));
 sky130_fd_sc_hd__a2111oi_2 _27932_ (.A1(_24686_),
    .A2(_24687_),
    .B1(_24717_),
    .C1(_24722_),
    .D1(_24723_),
    .Y(_24724_));
 sky130_fd_sc_hd__a21o_1 _27933_ (.A1(_24687_),
    .A2(_24686_),
    .B1(_24722_),
    .X(_24725_));
 sky130_fd_sc_hd__o21a_1 _27934_ (.A1(_24717_),
    .A2(_24723_),
    .B1(_24725_),
    .X(_24726_));
 sky130_fd_sc_hd__nor3_4 _27935_ (.A(_24652_),
    .B(net110),
    .C(_24726_),
    .Y(_24727_));
 sky130_fd_sc_hd__o21ai_1 _27936_ (.A1(net110),
    .A2(_24726_),
    .B1(_24652_),
    .Y(_24728_));
 sky130_fd_sc_hd__or2b_1 _27937_ (.A(_24727_),
    .B_N(_24728_),
    .X(_24729_));
 sky130_fd_sc_hd__a21boi_1 _27938_ (.A1(_23090_),
    .A2(_23093_),
    .B1_N(_23087_),
    .Y(_24730_));
 sky130_fd_sc_hd__a21oi_1 _27939_ (.A1(_07118_),
    .A2(_20606_),
    .B1(_16777_),
    .Y(_24731_));
 sky130_fd_sc_hd__a21o_1 _27940_ (.A1(_01798_),
    .A2(_07085_),
    .B1(_24731_),
    .X(_24733_));
 sky130_fd_sc_hd__and2_1 _27941_ (.A(\delay_line[15][8] ),
    .B(\delay_line[15][10] ),
    .X(_24734_));
 sky130_fd_sc_hd__clkbuf_2 _27942_ (.A(_24734_),
    .X(_24735_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27943_ (.A(\delay_line[15][10] ),
    .X(_24736_));
 sky130_fd_sc_hd__buf_2 _27944_ (.A(_24736_),
    .X(_24737_));
 sky130_fd_sc_hd__o211ai_4 _27945_ (.A1(_21452_),
    .A2(_24737_),
    .B1(_23078_),
    .C1(_20600_),
    .Y(_24738_));
 sky130_fd_sc_hd__inv_2 _27946_ (.A(net386),
    .Y(_24739_));
 sky130_fd_sc_hd__buf_2 _27947_ (.A(_24739_),
    .X(_24740_));
 sky130_fd_sc_hd__nor2_1 _27948_ (.A(\delay_line[15][8] ),
    .B(_24736_),
    .Y(_24741_));
 sky130_fd_sc_hd__o22ai_4 _27949_ (.A1(_20596_),
    .A2(_24740_),
    .B1(_24734_),
    .B2(_24741_),
    .Y(_24742_));
 sky130_fd_sc_hd__o211ai_4 _27950_ (.A1(_24735_),
    .A2(_24738_),
    .B1(_18416_),
    .C1(_24742_),
    .Y(_24744_));
 sky130_fd_sc_hd__buf_1 _27951_ (.A(_24737_),
    .X(_24745_));
 sky130_fd_sc_hd__a21o_1 _27952_ (.A1(_21459_),
    .A2(_24745_),
    .B1(_24738_),
    .X(_24746_));
 sky130_fd_sc_hd__a21o_1 _27953_ (.A1(_24746_),
    .A2(_24742_),
    .B1(_18422_),
    .X(_24747_));
 sky130_fd_sc_hd__o2bb2ai_2 _27954_ (.A1_N(_18411_),
    .A2_N(_23080_),
    .B1(_23077_),
    .B2(_23075_),
    .Y(_24748_));
 sky130_fd_sc_hd__nand3_2 _27955_ (.A(_24744_),
    .B(_24747_),
    .C(_24748_),
    .Y(_24749_));
 sky130_fd_sc_hd__o211a_1 _27956_ (.A1(_24735_),
    .A2(_24738_),
    .B1(_18422_),
    .C1(_24742_),
    .X(_24750_));
 sky130_fd_sc_hd__a21oi_1 _27957_ (.A1(_24746_),
    .A2(_24742_),
    .B1(_18423_),
    .Y(_24751_));
 sky130_fd_sc_hd__o21bai_2 _27958_ (.A1(_24750_),
    .A2(_24751_),
    .B1_N(_24748_),
    .Y(_24752_));
 sky130_fd_sc_hd__nand3b_1 _27959_ (.A_N(_24733_),
    .B(_24749_),
    .C(_24752_),
    .Y(_24753_));
 sky130_fd_sc_hd__a21bo_1 _27960_ (.A1(_24749_),
    .A2(_24752_),
    .B1_N(_24733_),
    .X(_24755_));
 sky130_fd_sc_hd__nand3b_1 _27961_ (.A_N(_24730_),
    .B(_24753_),
    .C(_24755_),
    .Y(_24756_));
 sky130_fd_sc_hd__a21o_1 _27962_ (.A1(_24749_),
    .A2(_24752_),
    .B1(_24733_),
    .X(_24757_));
 sky130_fd_sc_hd__nand3_1 _27963_ (.A(_24733_),
    .B(_24749_),
    .C(_24752_),
    .Y(_24758_));
 sky130_fd_sc_hd__nand3_1 _27964_ (.A(_24757_),
    .B(_24758_),
    .C(_24730_),
    .Y(_24759_));
 sky130_fd_sc_hd__or3b_1 _27965_ (.A(_01798_),
    .B(_07118_),
    .C_N(_22402_),
    .X(_24760_));
 sky130_fd_sc_hd__nand4_1 _27966_ (.A(_24756_),
    .B(_24094_),
    .C(_24759_),
    .D(_24760_),
    .Y(_24761_));
 sky130_fd_sc_hd__and3_1 _27967_ (.A(_16722_),
    .B(_24094_),
    .C(_22413_),
    .X(_24762_));
 sky130_fd_sc_hd__clkbuf_2 _27968_ (.A(_07118_),
    .X(_24763_));
 sky130_fd_sc_hd__o2bb2ai_1 _27969_ (.A1_N(_24759_),
    .A2_N(_24756_),
    .B1(_24762_),
    .B2(_24763_),
    .Y(_24764_));
 sky130_fd_sc_hd__nand2_1 _27970_ (.A(_24761_),
    .B(_24764_),
    .Y(_24766_));
 sky130_fd_sc_hd__a21oi_1 _27971_ (.A1(_23100_),
    .A2(_23101_),
    .B1(_24766_),
    .Y(_24767_));
 sky130_fd_sc_hd__and3_1 _27972_ (.A(_23102_),
    .B(_21479_),
    .C(_23101_),
    .X(_24768_));
 sky130_fd_sc_hd__a21boi_1 _27973_ (.A1(_23097_),
    .A2(_22424_),
    .B1_N(_23100_),
    .Y(_24769_));
 sky130_fd_sc_hd__nand2_1 _27974_ (.A(_24766_),
    .B(_24769_),
    .Y(_24770_));
 sky130_fd_sc_hd__nand3b_1 _27975_ (.A_N(_24767_),
    .B(_24768_),
    .C(_24770_),
    .Y(_24771_));
 sky130_fd_sc_hd__nand2_1 _27976_ (.A(_23101_),
    .B(_23102_),
    .Y(_24772_));
 sky130_fd_sc_hd__a21boi_1 _27977_ (.A1(_24761_),
    .A2(_24764_),
    .B1_N(_24769_),
    .Y(_24773_));
 sky130_fd_sc_hd__o22ai_1 _27978_ (.A1(_21476_),
    .A2(_24772_),
    .B1(_24773_),
    .B2(_24767_),
    .Y(_24774_));
 sky130_fd_sc_hd__nand2_1 _27979_ (.A(_24771_),
    .B(_24774_),
    .Y(_24775_));
 sky130_fd_sc_hd__nand2_1 _27980_ (.A(_23103_),
    .B(_23104_),
    .Y(_24777_));
 sky130_fd_sc_hd__o32ai_1 _27981_ (.A1(_20595_),
    .A2(_21446_),
    .A3(_21482_),
    .B1(_20622_),
    .B2(_21485_),
    .Y(_24778_));
 sky130_fd_sc_hd__a2bb2oi_1 _27982_ (.A1_N(_21477_),
    .A2_N(_24772_),
    .B1(_24777_),
    .B2(_24778_),
    .Y(_24779_));
 sky130_fd_sc_hd__or2_1 _27983_ (.A(_24775_),
    .B(_24779_),
    .X(_24780_));
 sky130_fd_sc_hd__o41ai_4 _27984_ (.A1(_21489_),
    .A2(_21500_),
    .A3(_21501_),
    .A4(_23064_),
    .B1(_23068_),
    .Y(_24781_));
 sky130_fd_sc_hd__and2_1 _27985_ (.A(_18405_),
    .B(net391),
    .X(_24782_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _27986_ (.A(\delay_line[14][9] ),
    .X(_24783_));
 sky130_fd_sc_hd__o21ai_2 _27987_ (.A1(_18405_),
    .A2(net391),
    .B1(_24783_),
    .Y(_24784_));
 sky130_fd_sc_hd__a21oi_2 _27988_ (.A1(_21491_),
    .A2(_18406_),
    .B1(_23056_),
    .Y(_24785_));
 sky130_fd_sc_hd__nor2_1 _27989_ (.A(_23052_),
    .B(_19450_),
    .Y(_24786_));
 sky130_fd_sc_hd__o21bai_2 _27990_ (.A1(_24782_),
    .A2(_24786_),
    .B1_N(_24783_),
    .Y(_24788_));
 sky130_fd_sc_hd__o211ai_4 _27991_ (.A1(_24782_),
    .A2(_24784_),
    .B1(_24785_),
    .C1(_24788_),
    .Y(_24789_));
 sky130_fd_sc_hd__a21o_1 _27992_ (.A1(_23052_),
    .A2(_19450_),
    .B1(_24784_),
    .X(_24790_));
 sky130_fd_sc_hd__a21o_1 _27993_ (.A1(_24790_),
    .A2(_24788_),
    .B1(_24785_),
    .X(_24791_));
 sky130_fd_sc_hd__a21oi_1 _27994_ (.A1(_16832_),
    .A2(_18406_),
    .B1(_01765_),
    .Y(_24792_));
 sky130_fd_sc_hd__and3_1 _27995_ (.A(net393),
    .B(_21491_),
    .C(_23052_),
    .X(_24793_));
 sky130_fd_sc_hd__nor2_1 _27996_ (.A(_24792_),
    .B(_24793_),
    .Y(_24794_));
 sky130_fd_sc_hd__a21bo_1 _27997_ (.A1(_24789_),
    .A2(_24791_),
    .B1_N(_24794_),
    .X(_24795_));
 sky130_fd_sc_hd__o211ai_1 _27998_ (.A1(_24792_),
    .A2(_24793_),
    .B1(_24789_),
    .C1(_24791_),
    .Y(_24796_));
 sky130_fd_sc_hd__o21ba_1 _27999_ (.A1(_23061_),
    .A2(_23059_),
    .B1_N(_23058_),
    .X(_24797_));
 sky130_fd_sc_hd__a21o_1 _28000_ (.A1(_24795_),
    .A2(_24796_),
    .B1(_24797_),
    .X(_24799_));
 sky130_fd_sc_hd__nand3_1 _28001_ (.A(_24795_),
    .B(_24796_),
    .C(_24797_),
    .Y(_24800_));
 sky130_fd_sc_hd__nand4_1 _28002_ (.A(_24799_),
    .B(_24061_),
    .C(_24800_),
    .D(_21495_),
    .Y(_24801_));
 sky130_fd_sc_hd__a32o_1 _28003_ (.A1(_24061_),
    .A2(_16832_),
    .A3(_07184_),
    .B1(_24800_),
    .B2(_24799_),
    .X(_24802_));
 sky130_fd_sc_hd__and4bb_1 _28004_ (.A_N(_21499_),
    .B_N(_23064_),
    .C(_24801_),
    .D(_24802_),
    .X(_24803_));
 sky130_fd_sc_hd__a2bb2o_1 _28005_ (.A1_N(_21499_),
    .A2_N(_23064_),
    .B1(_24801_),
    .B2(_24802_),
    .X(_24804_));
 sky130_fd_sc_hd__or2b_1 _28006_ (.A(_24803_),
    .B_N(_24804_),
    .X(_24805_));
 sky130_fd_sc_hd__xnor2_2 _28007_ (.A(_24781_),
    .B(_24805_),
    .Y(_24806_));
 sky130_fd_sc_hd__nand2_1 _28008_ (.A(_24779_),
    .B(_24775_),
    .Y(_24807_));
 sky130_fd_sc_hd__nand3_2 _28009_ (.A(_24780_),
    .B(_24806_),
    .C(_24807_),
    .Y(_24808_));
 sky130_fd_sc_hd__a21o_1 _28010_ (.A1(_24807_),
    .A2(_24780_),
    .B1(_24806_),
    .X(_24810_));
 sky130_fd_sc_hd__and2_1 _28011_ (.A(_24808_),
    .B(_24810_),
    .X(_24811_));
 sky130_fd_sc_hd__o21ai_1 _28012_ (.A1(_16601_),
    .A2(_23020_),
    .B1(_23017_),
    .Y(_24812_));
 sky130_fd_sc_hd__and2_1 _28013_ (.A(\delay_line[16][5] ),
    .B(net385),
    .X(_24813_));
 sky130_fd_sc_hd__or2_1 _28014_ (.A(\delay_line[16][5] ),
    .B(\delay_line[16][6] ),
    .X(_24814_));
 sky130_fd_sc_hd__nand3b_1 _28015_ (.A_N(_24813_),
    .B(_18399_),
    .C(_24814_),
    .Y(_24815_));
 sky130_fd_sc_hd__buf_1 _28016_ (.A(net385),
    .X(_24816_));
 sky130_fd_sc_hd__nor2_1 _28017_ (.A(_23016_),
    .B(_24816_),
    .Y(_24817_));
 sky130_fd_sc_hd__o21bai_1 _28018_ (.A1(_24817_),
    .A2(_24813_),
    .B1_N(_21514_),
    .Y(_24818_));
 sky130_fd_sc_hd__clkbuf_2 _28019_ (.A(\delay_line[16][9] ),
    .X(_24819_));
 sky130_fd_sc_hd__clkbuf_2 _28020_ (.A(_24819_),
    .X(_24821_));
 sky130_fd_sc_hd__nand3_2 _28021_ (.A(_24815_),
    .B(_24818_),
    .C(_24821_),
    .Y(_24822_));
 sky130_fd_sc_hd__buf_1 _28022_ (.A(_24822_),
    .X(_24823_));
 sky130_fd_sc_hd__a21o_1 _28023_ (.A1(_24815_),
    .A2(_24818_),
    .B1(_24821_),
    .X(_24824_));
 sky130_fd_sc_hd__a21o_1 _28024_ (.A1(_24823_),
    .A2(_24824_),
    .B1(_23027_),
    .X(_24825_));
 sky130_fd_sc_hd__nand3_1 _28025_ (.A(_23027_),
    .B(_24823_),
    .C(_24824_),
    .Y(_24826_));
 sky130_fd_sc_hd__nand3_1 _28026_ (.A(_24812_),
    .B(_24825_),
    .C(_24826_),
    .Y(_24827_));
 sky130_fd_sc_hd__nand3_1 _28027_ (.A(_23030_),
    .B(_24823_),
    .C(_24824_),
    .Y(_24828_));
 sky130_fd_sc_hd__a32o_1 _28028_ (.A1(_23026_),
    .A2(_23019_),
    .A3(_23022_),
    .B1(_24822_),
    .B2(_24824_),
    .X(_24829_));
 sky130_fd_sc_hd__o2111ai_2 _28029_ (.A1(_16601_),
    .A2(_23020_),
    .B1(_23017_),
    .C1(_24828_),
    .D1(_24829_),
    .Y(_24830_));
 sky130_fd_sc_hd__nand2_1 _28030_ (.A(_24827_),
    .B(_24830_),
    .Y(_24832_));
 sky130_fd_sc_hd__a21boi_1 _28031_ (.A1(_23031_),
    .A2(_23032_),
    .B1_N(_23028_),
    .Y(_24833_));
 sky130_fd_sc_hd__nand2_1 _28032_ (.A(_24832_),
    .B(_24833_),
    .Y(_24834_));
 sky130_fd_sc_hd__buf_1 _28033_ (.A(_18400_),
    .X(_24835_));
 sky130_fd_sc_hd__o211a_1 _28034_ (.A1(_16612_),
    .A2(_24835_),
    .B1(_21536_),
    .C1(_24127_),
    .X(_24836_));
 sky130_fd_sc_hd__o21a_1 _28035_ (.A1(_07217_),
    .A2(_21519_),
    .B1(_16645_),
    .X(_24837_));
 sky130_fd_sc_hd__nor2_1 _28036_ (.A(_24836_),
    .B(_24837_),
    .Y(_24838_));
 sky130_fd_sc_hd__nand3b_1 _28037_ (.A_N(_24833_),
    .B(_24827_),
    .C(_24830_),
    .Y(_24839_));
 sky130_fd_sc_hd__nand3_2 _28038_ (.A(_24834_),
    .B(_24838_),
    .C(_24839_),
    .Y(_24840_));
 sky130_fd_sc_hd__a2bb2o_1 _28039_ (.A1_N(_24836_),
    .A2_N(_24837_),
    .B1(_24839_),
    .B2(_24834_),
    .X(_24841_));
 sky130_fd_sc_hd__a21bo_1 _28040_ (.A1(_23036_),
    .A2(_21511_),
    .B1_N(_23035_),
    .X(_24843_));
 sky130_fd_sc_hd__a21oi_1 _28041_ (.A1(_24840_),
    .A2(_24841_),
    .B1(_24843_),
    .Y(_24844_));
 sky130_fd_sc_hd__and3_1 _28042_ (.A(_24843_),
    .B(_24840_),
    .C(_24841_),
    .X(_24845_));
 sky130_fd_sc_hd__or2_1 _28043_ (.A(_24844_),
    .B(_24845_),
    .X(_24846_));
 sky130_fd_sc_hd__a22oi_4 _28044_ (.A1(_23044_),
    .A2(_23043_),
    .B1(_23042_),
    .B2(_23041_),
    .Y(_24847_));
 sky130_fd_sc_hd__xor2_2 _28045_ (.A(_24846_),
    .B(_24847_),
    .X(_24848_));
 sky130_fd_sc_hd__xnor2_2 _28046_ (.A(_24811_),
    .B(_24848_),
    .Y(_24849_));
 sky130_fd_sc_hd__a21o_2 _28047_ (.A1(_23108_),
    .A2(_23112_),
    .B1(_24849_),
    .X(_24850_));
 sky130_fd_sc_hd__or2_1 _28048_ (.A(_23105_),
    .B(_23107_),
    .X(_24851_));
 sky130_fd_sc_hd__o211ai_4 _28049_ (.A1(_23070_),
    .A2(_24851_),
    .B1(_23112_),
    .C1(_24849_),
    .Y(_24852_));
 sky130_fd_sc_hd__nand2_1 _28050_ (.A(_24850_),
    .B(_24852_),
    .Y(_24854_));
 sky130_fd_sc_hd__xnor2_2 _28051_ (.A(_24729_),
    .B(_24854_),
    .Y(_24855_));
 sky130_fd_sc_hd__and3_1 _28052_ (.A(_23115_),
    .B(_24623_),
    .C(_24855_),
    .X(_24856_));
 sky130_fd_sc_hd__a21oi_4 _28053_ (.A1(_23115_),
    .A2(_24623_),
    .B1(_24855_),
    .Y(_24857_));
 sky130_fd_sc_hd__nor2_2 _28054_ (.A(_24856_),
    .B(_24857_),
    .Y(_24858_));
 sky130_fd_sc_hd__xnor2_1 _28055_ (.A(_24621_),
    .B(_24858_),
    .Y(_24859_));
 sky130_fd_sc_hd__or2b_1 _28056_ (.A(_24495_),
    .B_N(_24859_),
    .X(_24860_));
 sky130_fd_sc_hd__or2b_1 _28057_ (.A(_24859_),
    .B_N(_24495_),
    .X(_24861_));
 sky130_fd_sc_hd__nand2_1 _28058_ (.A(_24860_),
    .B(_24861_),
    .Y(_24862_));
 sky130_fd_sc_hd__xnor2_1 _28059_ (.A(_24493_),
    .B(_24862_),
    .Y(_24863_));
 sky130_fd_sc_hd__a21o_1 _28060_ (.A1(_23121_),
    .A2(_23302_),
    .B1(_24863_),
    .X(_24865_));
 sky130_fd_sc_hd__o211ai_1 _28061_ (.A1(_23123_),
    .A2(_23301_),
    .B1(_24863_),
    .C1(_23121_),
    .Y(_24866_));
 sky130_fd_sc_hd__nand2_1 _28062_ (.A(_24865_),
    .B(_24866_),
    .Y(_24867_));
 sky130_fd_sc_hd__o21a_1 _28063_ (.A1(_23300_),
    .A2(_23299_),
    .B1(_23298_),
    .X(_24868_));
 sky130_fd_sc_hd__nand2_1 _28064_ (.A(_23422_),
    .B(_23424_),
    .Y(_24869_));
 sky130_fd_sc_hd__or3b_1 _28065_ (.A(_23417_),
    .B(_23342_),
    .C_N(_23416_),
    .X(_24870_));
 sky130_fd_sc_hd__or2_1 _28066_ (.A(_23239_),
    .B(_23240_),
    .X(_24871_));
 sky130_fd_sc_hd__a21boi_1 _28067_ (.A1(_23335_),
    .A2(_21098_),
    .B1_N(_23336_),
    .Y(_24872_));
 sky130_fd_sc_hd__buf_1 _28068_ (.A(_18633_),
    .X(_24873_));
 sky130_fd_sc_hd__buf_1 _28069_ (.A(\delay_line[34][6] ),
    .X(_24874_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28070_ (.A(_24874_),
    .X(_24876_));
 sky130_fd_sc_hd__a21boi_1 _28071_ (.A1(_24873_),
    .A2(_24876_),
    .B1_N(_05403_),
    .Y(_24877_));
 sky130_fd_sc_hd__and3b_1 _28072_ (.A_N(_05403_),
    .B(_18633_),
    .C(_24874_),
    .X(_24878_));
 sky130_fd_sc_hd__nor2_1 _28073_ (.A(_21085_),
    .B(\delay_line[34][10] ),
    .Y(_24879_));
 sky130_fd_sc_hd__buf_1 _28074_ (.A(\delay_line[34][10] ),
    .X(_24880_));
 sky130_fd_sc_hd__nand2_1 _28075_ (.A(_21085_),
    .B(_24880_),
    .Y(_24881_));
 sky130_fd_sc_hd__nand3b_1 _28076_ (.A_N(_24879_),
    .B(_23317_),
    .C(_24881_),
    .Y(_24882_));
 sky130_fd_sc_hd__and2_1 _28077_ (.A(_21085_),
    .B(\delay_line[34][10] ),
    .X(_24883_));
 sky130_fd_sc_hd__o21ai_2 _28078_ (.A1(_24883_),
    .A2(_24879_),
    .B1(_23313_),
    .Y(_24884_));
 sky130_fd_sc_hd__nor2_1 _28079_ (.A(_24874_),
    .B(_20741_),
    .Y(_24885_));
 sky130_fd_sc_hd__and2_1 _28080_ (.A(_19553_),
    .B(_20743_),
    .X(_24887_));
 sky130_fd_sc_hd__nor2_1 _28081_ (.A(_24885_),
    .B(_24887_),
    .Y(_24888_));
 sky130_fd_sc_hd__a21bo_1 _28082_ (.A1(_24882_),
    .A2(_24884_),
    .B1_N(_24888_),
    .X(_24889_));
 sky130_fd_sc_hd__o211ai_1 _28083_ (.A1(_24885_),
    .A2(_24887_),
    .B1(_24882_),
    .C1(_24884_),
    .Y(_24890_));
 sky130_fd_sc_hd__nand4_1 _28084_ (.A(_23316_),
    .B(_23327_),
    .C(_24889_),
    .D(_24890_),
    .Y(_24891_));
 sky130_fd_sc_hd__a22o_1 _28085_ (.A1(_23316_),
    .A2(_23327_),
    .B1(_24889_),
    .B2(_24890_),
    .X(_24892_));
 sky130_fd_sc_hd__a2bb2o_1 _28086_ (.A1_N(_24877_),
    .A2_N(_24878_),
    .B1(_24891_),
    .B2(_24892_),
    .X(_24893_));
 sky130_fd_sc_hd__nor2_1 _28087_ (.A(_24877_),
    .B(_24878_),
    .Y(_24894_));
 sky130_fd_sc_hd__nand3_2 _28088_ (.A(_24892_),
    .B(_24894_),
    .C(_24891_),
    .Y(_24895_));
 sky130_fd_sc_hd__nand2_1 _28089_ (.A(_23329_),
    .B(_23332_),
    .Y(_24896_));
 sky130_fd_sc_hd__a21oi_1 _28090_ (.A1(_24893_),
    .A2(_24895_),
    .B1(_24896_),
    .Y(_24898_));
 sky130_fd_sc_hd__nand3_1 _28091_ (.A(_24896_),
    .B(_24893_),
    .C(_24895_),
    .Y(_24899_));
 sky130_fd_sc_hd__or4bb_1 _28092_ (.A(_02249_),
    .B(_24898_),
    .C_N(_24899_),
    .D_N(_20737_),
    .X(_24900_));
 sky130_fd_sc_hd__and3_1 _28093_ (.A(_24896_),
    .B(_24893_),
    .C(_24895_),
    .X(_24901_));
 sky130_fd_sc_hd__o22ai_1 _28094_ (.A1(_02260_),
    .A2(_21097_),
    .B1(_24898_),
    .B2(_24901_),
    .Y(_24902_));
 sky130_fd_sc_hd__nand2_1 _28095_ (.A(_24900_),
    .B(_24902_),
    .Y(_24903_));
 sky130_fd_sc_hd__xor2_1 _28096_ (.A(_24872_),
    .B(_24903_),
    .X(_24904_));
 sky130_fd_sc_hd__nand2_1 _28097_ (.A(_23340_),
    .B(_23310_),
    .Y(_24905_));
 sky130_fd_sc_hd__nor2_1 _28098_ (.A(_23310_),
    .B(_23340_),
    .Y(_24906_));
 sky130_fd_sc_hd__a31o_1 _28099_ (.A1(_24905_),
    .A2(_21108_),
    .A3(_21109_),
    .B1(_24906_),
    .X(_24907_));
 sky130_fd_sc_hd__xor2_1 _28100_ (.A(_24904_),
    .B(_24907_),
    .X(_24909_));
 sky130_fd_sc_hd__a21boi_2 _28101_ (.A1(_21175_),
    .A2(_23380_),
    .B1_N(_23379_),
    .Y(_24910_));
 sky130_fd_sc_hd__nand3_2 _28102_ (.A(_23346_),
    .B(_23376_),
    .C(_23374_),
    .Y(_24911_));
 sky130_fd_sc_hd__nand2_1 _28103_ (.A(_23376_),
    .B(_24911_),
    .Y(_24912_));
 sky130_fd_sc_hd__buf_1 _28104_ (.A(net312),
    .X(_24913_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28105_ (.A(_23350_),
    .X(_24914_));
 sky130_fd_sc_hd__nor3_1 _28106_ (.A(_02161_),
    .B(_24913_),
    .C(_24914_),
    .Y(_24915_));
 sky130_fd_sc_hd__o21a_1 _28107_ (.A1(_23352_),
    .A2(_24914_),
    .B1(_19570_),
    .X(_24916_));
 sky130_fd_sc_hd__o22ai_2 _28108_ (.A1(_23367_),
    .A2(_00568_),
    .B1(_24915_),
    .B2(_24916_),
    .Y(_24917_));
 sky130_fd_sc_hd__nor2_1 _28109_ (.A(_19570_),
    .B(_24913_),
    .Y(_24918_));
 sky130_fd_sc_hd__a2111o_1 _28110_ (.A1(_17822_),
    .A2(_24918_),
    .B1(_23367_),
    .C1(_00557_),
    .D1(_24916_),
    .X(_24920_));
 sky130_fd_sc_hd__clkbuf_2 _28111_ (.A(_23349_),
    .X(_24921_));
 sky130_fd_sc_hd__clkbuf_2 _28112_ (.A(\delay_line[33][10] ),
    .X(_24922_));
 sky130_fd_sc_hd__and2b_1 _28113_ (.A_N(\delay_line[33][6] ),
    .B(net312),
    .X(_24923_));
 sky130_fd_sc_hd__and2b_1 _28114_ (.A_N(\delay_line[33][5] ),
    .B(\delay_line[33][6] ),
    .X(_24924_));
 sky130_fd_sc_hd__nor3_2 _28115_ (.A(_24922_),
    .B(_24923_),
    .C(_24924_),
    .Y(_24925_));
 sky130_fd_sc_hd__o21a_1 _28116_ (.A1(_24923_),
    .A2(_24924_),
    .B1(_24922_),
    .X(_24926_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28117_ (.A(_24926_),
    .X(_24927_));
 sky130_fd_sc_hd__a211o_1 _28118_ (.A1(_24921_),
    .A2(_23355_),
    .B1(_24925_),
    .C1(_24927_),
    .X(_24928_));
 sky130_fd_sc_hd__o211ai_2 _28119_ (.A1(_24925_),
    .A2(_24927_),
    .B1(_24921_),
    .C1(_23355_),
    .Y(_24929_));
 sky130_fd_sc_hd__nand4_2 _28120_ (.A(_24917_),
    .B(_24920_),
    .C(_24928_),
    .D(_24929_),
    .Y(_24931_));
 sky130_fd_sc_hd__a211oi_1 _28121_ (.A1(_24921_),
    .A2(_23355_),
    .B1(_24925_),
    .C1(_24927_),
    .Y(_24932_));
 sky130_fd_sc_hd__o211a_1 _28122_ (.A1(_24925_),
    .A2(_24927_),
    .B1(_24921_),
    .C1(_23355_),
    .X(_24933_));
 sky130_fd_sc_hd__nand2_1 _28123_ (.A(_24917_),
    .B(_24920_),
    .Y(_24934_));
 sky130_fd_sc_hd__o21ai_1 _28124_ (.A1(_24932_),
    .A2(_24933_),
    .B1(_24934_),
    .Y(_24935_));
 sky130_fd_sc_hd__a21bo_1 _28125_ (.A1(_23365_),
    .A2(_23369_),
    .B1_N(_23363_),
    .X(_24936_));
 sky130_fd_sc_hd__a21o_1 _28126_ (.A1(_24931_),
    .A2(_24935_),
    .B1(_24936_),
    .X(_24937_));
 sky130_fd_sc_hd__nand3_1 _28127_ (.A(_24936_),
    .B(_24931_),
    .C(_24935_),
    .Y(_24938_));
 sky130_fd_sc_hd__nand4_1 _28128_ (.A(_24937_),
    .B(_24938_),
    .C(_05348_),
    .D(_19572_),
    .Y(_24939_));
 sky130_fd_sc_hd__a32o_1 _28129_ (.A1(_00590_),
    .A2(_02183_),
    .A3(_05348_),
    .B1(_24937_),
    .B2(_24938_),
    .X(_24940_));
 sky130_fd_sc_hd__nand2_2 _28130_ (.A(_24939_),
    .B(_24940_),
    .Y(_24942_));
 sky130_fd_sc_hd__xor2_2 _28131_ (.A(_24912_),
    .B(_24942_),
    .X(_24943_));
 sky130_fd_sc_hd__and2_1 _28132_ (.A(_24910_),
    .B(_24943_),
    .X(_24944_));
 sky130_fd_sc_hd__nor2_1 _28133_ (.A(_24943_),
    .B(_24910_),
    .Y(_24945_));
 sky130_fd_sc_hd__and2_1 _28134_ (.A(_23408_),
    .B(_23384_),
    .X(_24946_));
 sky130_fd_sc_hd__buf_1 _28135_ (.A(_23405_),
    .X(_24947_));
 sky130_fd_sc_hd__a41o_1 _28136_ (.A1(_23407_),
    .A2(_21140_),
    .A3(_21139_),
    .A4(_21138_),
    .B1(_24947_),
    .X(_24948_));
 sky130_fd_sc_hd__nand2_2 _28137_ (.A(_05216_),
    .B(_18659_),
    .Y(_24949_));
 sky130_fd_sc_hd__nand2_1 _28138_ (.A(_18672_),
    .B(_02106_),
    .Y(_24950_));
 sky130_fd_sc_hd__and4_2 _28139_ (.A(_24523_),
    .B(_24949_),
    .C(_24950_),
    .D(_05304_),
    .X(_24951_));
 sky130_fd_sc_hd__o2bb2a_1 _28140_ (.A1_N(_24949_),
    .A2_N(_24950_),
    .B1(_24457_),
    .B2(_05260_),
    .X(_24953_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28141_ (.A(\delay_line[32][9] ),
    .X(_24954_));
 sky130_fd_sc_hd__nor2_1 _28142_ (.A(_24954_),
    .B(\delay_line[32][10] ),
    .Y(_24955_));
 sky130_fd_sc_hd__buf_1 _28143_ (.A(\delay_line[32][10] ),
    .X(_24956_));
 sky130_fd_sc_hd__nand2_1 _28144_ (.A(_24954_),
    .B(_24956_),
    .Y(_24957_));
 sky130_fd_sc_hd__nand3b_1 _28145_ (.A_N(_24955_),
    .B(_24957_),
    .C(_21115_),
    .Y(_24958_));
 sky130_fd_sc_hd__and2_1 _28146_ (.A(_24954_),
    .B(\delay_line[32][10] ),
    .X(_24959_));
 sky130_fd_sc_hd__o21ai_1 _28147_ (.A1(_24955_),
    .A2(_24959_),
    .B1(_21113_),
    .Y(_24960_));
 sky130_fd_sc_hd__nor2_1 _28148_ (.A(\delay_line[32][8] ),
    .B(_24954_),
    .Y(_24961_));
 sky130_fd_sc_hd__nand2_1 _28149_ (.A(_21115_),
    .B(_23389_),
    .Y(_24962_));
 sky130_fd_sc_hd__o21ai_1 _28150_ (.A1(_20689_),
    .A2(_24961_),
    .B1(_24962_),
    .Y(_24964_));
 sky130_fd_sc_hd__and3_1 _28151_ (.A(_24958_),
    .B(_24960_),
    .C(_24964_),
    .X(_24965_));
 sky130_fd_sc_hd__a21o_1 _28152_ (.A1(_24958_),
    .A2(_24960_),
    .B1(_24964_),
    .X(_24966_));
 sky130_fd_sc_hd__nand3b_2 _28153_ (.A_N(_24965_),
    .B(_24966_),
    .C(_21126_),
    .Y(_24967_));
 sky130_fd_sc_hd__a21oi_1 _28154_ (.A1(_24958_),
    .A2(_24960_),
    .B1(_24964_),
    .Y(_24968_));
 sky130_fd_sc_hd__buf_1 _28155_ (.A(_20690_),
    .X(_24969_));
 sky130_fd_sc_hd__o21ai_2 _28156_ (.A1(_24965_),
    .A2(_24968_),
    .B1(_24969_),
    .Y(_24970_));
 sky130_fd_sc_hd__clkbuf_2 _28157_ (.A(_23393_),
    .X(_24971_));
 sky130_fd_sc_hd__a31o_1 _28158_ (.A1(_21114_),
    .A2(_23391_),
    .A3(_24971_),
    .B1(_23394_),
    .X(_24972_));
 sky130_fd_sc_hd__a21oi_1 _28159_ (.A1(_24967_),
    .A2(_24970_),
    .B1(_24972_),
    .Y(_24973_));
 sky130_fd_sc_hd__and3_1 _28160_ (.A(_24972_),
    .B(_24967_),
    .C(_24970_),
    .X(_24975_));
 sky130_fd_sc_hd__o22ai_2 _28161_ (.A1(_24951_),
    .A2(_24953_),
    .B1(_24973_),
    .B2(_24975_),
    .Y(_24976_));
 sky130_fd_sc_hd__a21o_1 _28162_ (.A1(_24967_),
    .A2(_24970_),
    .B1(_24972_),
    .X(_24977_));
 sky130_fd_sc_hd__nand3_1 _28163_ (.A(_24972_),
    .B(_24967_),
    .C(_24970_),
    .Y(_24978_));
 sky130_fd_sc_hd__nor2_1 _28164_ (.A(_24951_),
    .B(_24953_),
    .Y(_24979_));
 sky130_fd_sc_hd__nand3_1 _28165_ (.A(_24977_),
    .B(_24978_),
    .C(_24979_),
    .Y(_24980_));
 sky130_fd_sc_hd__o211ai_2 _28166_ (.A1(_23398_),
    .A2(_23401_),
    .B1(_24976_),
    .C1(_24980_),
    .Y(_24981_));
 sky130_fd_sc_hd__a211o_1 _28167_ (.A1(_24976_),
    .A2(_24980_),
    .B1(_23398_),
    .C1(_23401_),
    .X(_24982_));
 sky130_fd_sc_hd__a32o_1 _28168_ (.A1(_19587_),
    .A2(_23385_),
    .A3(_23386_),
    .B1(_24981_),
    .B2(_24982_),
    .X(_24983_));
 sky130_fd_sc_hd__nand3_1 _28169_ (.A(_24982_),
    .B(_23387_),
    .C(_24981_),
    .Y(_24984_));
 sky130_fd_sc_hd__nand2_2 _28170_ (.A(_24983_),
    .B(_24984_),
    .Y(_24986_));
 sky130_fd_sc_hd__xnor2_2 _28171_ (.A(_24948_),
    .B(_24986_),
    .Y(_24987_));
 sky130_fd_sc_hd__o21a_1 _28172_ (.A1(_24946_),
    .A2(_23410_),
    .B1(_24987_),
    .X(_24988_));
 sky130_fd_sc_hd__xnor2_1 _28173_ (.A(_23384_),
    .B(_23408_),
    .Y(_24989_));
 sky130_fd_sc_hd__a21o_1 _28174_ (.A1(_21145_),
    .A2(_21148_),
    .B1(_21151_),
    .X(_24990_));
 sky130_fd_sc_hd__o22ai_1 _28175_ (.A1(_20727_),
    .A2(_20726_),
    .B1(_20729_),
    .B2(_20725_),
    .Y(_24991_));
 sky130_fd_sc_hd__a21oi_1 _28176_ (.A1(_24990_),
    .A2(_24991_),
    .B1(_21157_),
    .Y(_24992_));
 sky130_fd_sc_hd__o21bai_1 _28177_ (.A1(_24989_),
    .A2(_24992_),
    .B1_N(_24946_),
    .Y(_24993_));
 sky130_fd_sc_hd__nor2_1 _28178_ (.A(_24987_),
    .B(_24993_),
    .Y(_24994_));
 sky130_fd_sc_hd__o22a_1 _28179_ (.A1(_24944_),
    .A2(_24945_),
    .B1(_24988_),
    .B2(_24994_),
    .X(_24995_));
 sky130_fd_sc_hd__nor4_1 _28180_ (.A(_24944_),
    .B(_24945_),
    .C(_24988_),
    .D(_24994_),
    .Y(_24997_));
 sky130_fd_sc_hd__nor2_1 _28181_ (.A(_24995_),
    .B(_24997_),
    .Y(_24998_));
 sky130_fd_sc_hd__and2_1 _28182_ (.A(_24909_),
    .B(_24998_),
    .X(_24999_));
 sky130_fd_sc_hd__nor2_1 _28183_ (.A(_24909_),
    .B(_24998_),
    .Y(_25000_));
 sky130_fd_sc_hd__or2_2 _28184_ (.A(_24999_),
    .B(_25000_),
    .X(_25001_));
 sky130_fd_sc_hd__o211ai_1 _28185_ (.A1(_24871_),
    .A2(_23286_),
    .B1(_23290_),
    .C1(_25001_),
    .Y(_25002_));
 sky130_fd_sc_hd__a21o_2 _28186_ (.A1(_23288_),
    .A2(_23290_),
    .B1(_25001_),
    .X(_25003_));
 sky130_fd_sc_hd__nand2_2 _28187_ (.A(_25002_),
    .B(_25003_),
    .Y(_25004_));
 sky130_fd_sc_hd__a21o_1 _28188_ (.A1(_23416_),
    .A2(_24870_),
    .B1(_25004_),
    .X(_25005_));
 sky130_fd_sc_hd__o211ai_1 _28189_ (.A1(_23417_),
    .A2(_23342_),
    .B1(_23416_),
    .C1(_25004_),
    .Y(_25006_));
 sky130_fd_sc_hd__nand2_1 _28190_ (.A(_25005_),
    .B(_25006_),
    .Y(_25008_));
 sky130_fd_sc_hd__and2b_1 _28191_ (.A_N(_24869_),
    .B(_25008_),
    .X(_25009_));
 sky130_fd_sc_hd__and2b_1 _28192_ (.A_N(_25008_),
    .B(_24869_),
    .X(_25010_));
 sky130_fd_sc_hd__nor2_1 _28193_ (.A(_25009_),
    .B(_25010_),
    .Y(_25011_));
 sky130_fd_sc_hd__nand2_1 _28194_ (.A(net281),
    .B(_23443_),
    .Y(_25012_));
 sky130_fd_sc_hd__nor2_1 _28195_ (.A(_23443_),
    .B(\delay_line[39][10] ),
    .Y(_25013_));
 sky130_fd_sc_hd__and2_1 _28196_ (.A(_23443_),
    .B(\delay_line[39][10] ),
    .X(_25014_));
 sky130_fd_sc_hd__or3_1 _28197_ (.A(_23445_),
    .B(_25013_),
    .C(_25014_),
    .X(_25015_));
 sky130_fd_sc_hd__o21ai_1 _28198_ (.A1(_25013_),
    .A2(_25014_),
    .B1(_23445_),
    .Y(_25016_));
 sky130_fd_sc_hd__nand2_1 _28199_ (.A(_25015_),
    .B(_25016_),
    .Y(_25017_));
 sky130_fd_sc_hd__a21oi_2 _28200_ (.A1(_25012_),
    .A2(_23449_),
    .B1(_25017_),
    .Y(_25019_));
 sky130_fd_sc_hd__a311oi_2 _28201_ (.A1(_23444_),
    .A2(_25012_),
    .A3(_25017_),
    .B1(_20986_),
    .C1(_25019_),
    .Y(_25020_));
 sky130_fd_sc_hd__and3_1 _28202_ (.A(_25012_),
    .B(_23449_),
    .C(_25017_),
    .X(_25021_));
 sky130_fd_sc_hd__o21a_1 _28203_ (.A1(_25019_),
    .A2(_25021_),
    .B1(_20986_),
    .X(_25022_));
 sky130_fd_sc_hd__or2_1 _28204_ (.A(_25020_),
    .B(_25022_),
    .X(_25023_));
 sky130_fd_sc_hd__or2b_1 _28205_ (.A(_23452_),
    .B_N(_25023_),
    .X(_25024_));
 sky130_fd_sc_hd__o21bai_1 _28206_ (.A1(_23452_),
    .A2(_23453_),
    .B1_N(_25023_),
    .Y(_25025_));
 sky130_fd_sc_hd__o221a_2 _28207_ (.A1(_25024_),
    .A2(_23453_),
    .B1(_23459_),
    .B2(_23462_),
    .C1(_25025_),
    .X(_25026_));
 sky130_fd_sc_hd__o21a_1 _28208_ (.A1(_23453_),
    .A2(_25024_),
    .B1(_25025_),
    .X(_25027_));
 sky130_fd_sc_hd__or3_1 _28209_ (.A(_23459_),
    .B(_23462_),
    .C(_25027_),
    .X(_25028_));
 sky130_fd_sc_hd__inv_2 _28210_ (.A(_25028_),
    .Y(_25030_));
 sky130_fd_sc_hd__nor2_1 _28211_ (.A(_23434_),
    .B(\delay_line[38][10] ),
    .Y(_25031_));
 sky130_fd_sc_hd__and2_2 _28212_ (.A(_23434_),
    .B(\delay_line[38][10] ),
    .X(_25032_));
 sky130_fd_sc_hd__nor2_1 _28213_ (.A(_25031_),
    .B(_25032_),
    .Y(_25033_));
 sky130_fd_sc_hd__clkbuf_2 _28214_ (.A(_25033_),
    .X(_25034_));
 sky130_fd_sc_hd__o21ai_1 _28215_ (.A1(_23429_),
    .A2(net286),
    .B1(_21005_),
    .Y(_25035_));
 sky130_fd_sc_hd__and3_1 _28216_ (.A(_25034_),
    .B(_25035_),
    .C(_23432_),
    .X(_25036_));
 sky130_fd_sc_hd__a21oi_1 _28217_ (.A1(_23432_),
    .A2(_25035_),
    .B1(_25034_),
    .Y(_25037_));
 sky130_fd_sc_hd__a41o_1 _28218_ (.A1(_19649_),
    .A2(_23434_),
    .A3(_21006_),
    .A4(_23433_),
    .B1(_23439_),
    .X(_25038_));
 sky130_fd_sc_hd__or3_1 _28219_ (.A(_25036_),
    .B(_25037_),
    .C(_25038_),
    .X(_25039_));
 sky130_fd_sc_hd__o21ai_2 _28220_ (.A1(_25036_),
    .A2(_25037_),
    .B1(_25038_),
    .Y(_25041_));
 sky130_fd_sc_hd__nand2_1 _28221_ (.A(_25039_),
    .B(_25041_),
    .Y(_25042_));
 sky130_fd_sc_hd__o21a_1 _28222_ (.A1(_25026_),
    .A2(_25030_),
    .B1(_25042_),
    .X(_25043_));
 sky130_fd_sc_hd__inv_2 _28223_ (.A(_25043_),
    .Y(_25044_));
 sky130_fd_sc_hd__inv_2 _28224_ (.A(\delay_line[40][9] ),
    .Y(_25045_));
 sky130_fd_sc_hd__a31o_1 _28225_ (.A1(\delay_line[40][7] ),
    .A2(_23464_),
    .A3(_25045_),
    .B1(_23468_),
    .X(_25046_));
 sky130_fd_sc_hd__or3b_2 _28226_ (.A(\delay_line[40][10] ),
    .B(_25045_),
    .C_N(_21019_),
    .X(_25047_));
 sky130_fd_sc_hd__or3b_1 _28227_ (.A(_21019_),
    .B(_25045_),
    .C_N(\delay_line[40][10] ),
    .X(_25048_));
 sky130_fd_sc_hd__o211a_1 _28228_ (.A1(_23465_),
    .A2(\delay_line[40][10] ),
    .B1(_25047_),
    .C1(_25048_),
    .X(_25049_));
 sky130_fd_sc_hd__nand2_1 _28229_ (.A(_20771_),
    .B(_25049_),
    .Y(_25050_));
 sky130_fd_sc_hd__or2_1 _28230_ (.A(_20771_),
    .B(_25049_),
    .X(_25052_));
 sky130_fd_sc_hd__and3_1 _28231_ (.A(_25046_),
    .B(_25050_),
    .C(_25052_),
    .X(_25053_));
 sky130_fd_sc_hd__a21oi_1 _28232_ (.A1(_25050_),
    .A2(_25052_),
    .B1(_25046_),
    .Y(_25054_));
 sky130_fd_sc_hd__o211ai_1 _28233_ (.A1(net272),
    .A2(_23470_),
    .B1(_21020_),
    .C1(_21023_),
    .Y(_25055_));
 sky130_fd_sc_hd__a21oi_1 _28234_ (.A1(_25055_),
    .A2(_23473_),
    .B1(_23472_),
    .Y(_25056_));
 sky130_fd_sc_hd__or3_1 _28235_ (.A(_25053_),
    .B(_25054_),
    .C(_25056_),
    .X(_25057_));
 sky130_fd_sc_hd__o21ai_1 _28236_ (.A1(_25053_),
    .A2(_25054_),
    .B1(_25056_),
    .Y(_25058_));
 sky130_fd_sc_hd__and2_2 _28237_ (.A(_25057_),
    .B(_25058_),
    .X(_25059_));
 sky130_fd_sc_hd__or3_4 _28238_ (.A(_25042_),
    .B(_25026_),
    .C(_25030_),
    .X(_25060_));
 sky130_fd_sc_hd__and3_1 _28239_ (.A(_25044_),
    .B(_25059_),
    .C(_25060_),
    .X(_25061_));
 sky130_fd_sc_hd__a21oi_1 _28240_ (.A1(_25060_),
    .A2(_25044_),
    .B1(_25059_),
    .Y(_25063_));
 sky130_fd_sc_hd__or2_2 _28241_ (.A(_25061_),
    .B(_25063_),
    .X(_25064_));
 sky130_fd_sc_hd__a21oi_4 _28242_ (.A1(_23529_),
    .A2(_23518_),
    .B1(net116),
    .Y(_25065_));
 sky130_fd_sc_hd__or2b_1 _28243_ (.A(_21036_),
    .B_N(\delay_line[37][10] ),
    .X(_25066_));
 sky130_fd_sc_hd__or2b_1 _28244_ (.A(\delay_line[37][10] ),
    .B_N(_21036_),
    .X(_25067_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28245_ (.A(_23520_),
    .X(_25068_));
 sky130_fd_sc_hd__nor3_1 _28246_ (.A(_25068_),
    .B(_23522_),
    .C(_21035_),
    .Y(_25069_));
 sky130_fd_sc_hd__o2bb2a_1 _28247_ (.A1_N(_25066_),
    .A2_N(_25067_),
    .B1(_25069_),
    .B2(_25068_),
    .X(_25070_));
 sky130_fd_sc_hd__nor2_1 _28248_ (.A(_25068_),
    .B(_25069_),
    .Y(_25071_));
 sky130_fd_sc_hd__and3_1 _28249_ (.A(_25071_),
    .B(_25067_),
    .C(_25066_),
    .X(_25072_));
 sky130_fd_sc_hd__or2_2 _28250_ (.A(_25070_),
    .B(_25072_),
    .X(_25074_));
 sky130_fd_sc_hd__a41o_2 _28251_ (.A1(_23521_),
    .A2(_20817_),
    .A3(_21035_),
    .A4(_21037_),
    .B1(_23527_),
    .X(_25075_));
 sky130_fd_sc_hd__xnor2_4 _28252_ (.A(_25074_),
    .B(_25075_),
    .Y(_25076_));
 sky130_fd_sc_hd__buf_1 _28253_ (.A(\delay_line[36][6] ),
    .X(_25077_));
 sky130_fd_sc_hd__and3_1 _28254_ (.A(_25077_),
    .B(_20825_),
    .C(_21051_),
    .X(_25078_));
 sky130_fd_sc_hd__and2b_1 _28255_ (.A_N(_21049_),
    .B(net297),
    .X(_25079_));
 sky130_fd_sc_hd__and2b_1 _28256_ (.A_N(net297),
    .B(_21049_),
    .X(_25080_));
 sky130_fd_sc_hd__nor2_1 _28257_ (.A(_25079_),
    .B(_25080_),
    .Y(_25081_));
 sky130_fd_sc_hd__and3b_1 _28258_ (.A_N(_19715_),
    .B(_21049_),
    .C(_23486_),
    .X(_25082_));
 sky130_fd_sc_hd__or3_1 _28259_ (.A(_23484_),
    .B(_25081_),
    .C(_25082_),
    .X(_25083_));
 sky130_fd_sc_hd__o21ai_1 _28260_ (.A1(_23484_),
    .A2(_25082_),
    .B1(_25081_),
    .Y(_25085_));
 sky130_fd_sc_hd__o211a_1 _28261_ (.A1(_23490_),
    .A2(_25078_),
    .B1(_25083_),
    .C1(_25085_),
    .X(_25086_));
 sky130_fd_sc_hd__inv_2 _28262_ (.A(_25086_),
    .Y(_25087_));
 sky130_fd_sc_hd__a221o_1 _28263_ (.A1(_25077_),
    .A2(_23488_),
    .B1(_25085_),
    .B2(_25083_),
    .C1(_23490_),
    .X(_25088_));
 sky130_fd_sc_hd__nor2_1 _28264_ (.A(_05909_),
    .B(_23507_),
    .Y(_25089_));
 sky130_fd_sc_hd__nor3b_1 _28265_ (.A(_23497_),
    .B(_23498_),
    .C_N(_20838_),
    .Y(_25090_));
 sky130_fd_sc_hd__buf_1 _28266_ (.A(\delay_line[35][10] ),
    .X(_25091_));
 sky130_fd_sc_hd__nor2_1 _28267_ (.A(_23496_),
    .B(_25091_),
    .Y(_25092_));
 sky130_fd_sc_hd__and2_1 _28268_ (.A(\delay_line[35][9] ),
    .B(\delay_line[35][10] ),
    .X(_25093_));
 sky130_fd_sc_hd__or3b_1 _28269_ (.A(_25092_),
    .B(_25093_),
    .C_N(_23495_),
    .X(_25094_));
 sky130_fd_sc_hd__o21bai_1 _28270_ (.A1(_25092_),
    .A2(_25093_),
    .B1_N(_23495_),
    .Y(_25096_));
 sky130_fd_sc_hd__o211a_1 _28271_ (.A1(_23498_),
    .A2(_25090_),
    .B1(_25094_),
    .C1(_25096_),
    .X(_25097_));
 sky130_fd_sc_hd__clkbuf_2 _28272_ (.A(_23496_),
    .X(_25098_));
 sky130_fd_sc_hd__a221oi_2 _28273_ (.A1(_23503_),
    .A2(_25098_),
    .B1(_25094_),
    .B2(_25096_),
    .C1(_25090_),
    .Y(_25099_));
 sky130_fd_sc_hd__nor3b_2 _28274_ (.A(_25097_),
    .B(_25099_),
    .C_N(_23501_),
    .Y(_25100_));
 sky130_fd_sc_hd__o21bai_1 _28275_ (.A1(_25097_),
    .A2(_25099_),
    .B1_N(_23501_),
    .Y(_25101_));
 sky130_fd_sc_hd__inv_2 _28276_ (.A(_25101_),
    .Y(_25102_));
 sky130_fd_sc_hd__or3_1 _28277_ (.A(_19697_),
    .B(_25100_),
    .C(_25102_),
    .X(_25103_));
 sky130_fd_sc_hd__o21ai_1 _28278_ (.A1(_25100_),
    .A2(_25102_),
    .B1(_19697_),
    .Y(_25104_));
 sky130_fd_sc_hd__o211ai_2 _28279_ (.A1(_23505_),
    .A2(_25089_),
    .B1(_25103_),
    .C1(_25104_),
    .Y(_25105_));
 sky130_fd_sc_hd__a211o_1 _28280_ (.A1(_25103_),
    .A2(_25104_),
    .B1(_23505_),
    .C1(_25089_),
    .X(_25107_));
 sky130_fd_sc_hd__a221o_1 _28281_ (.A1(_25105_),
    .A2(_25107_),
    .B1(_23512_),
    .B2(_23511_),
    .C1(_23509_),
    .X(_25108_));
 sky130_fd_sc_hd__nand2_1 _28282_ (.A(_25105_),
    .B(_25107_),
    .Y(_25109_));
 sky130_fd_sc_hd__a21oi_1 _28283_ (.A1(_23512_),
    .A2(_23511_),
    .B1(_23509_),
    .Y(_25110_));
 sky130_fd_sc_hd__or2_1 _28284_ (.A(_25109_),
    .B(_25110_),
    .X(_25111_));
 sky130_fd_sc_hd__nand4_1 _28285_ (.A(_25087_),
    .B(_25088_),
    .C(_25108_),
    .D(_25111_),
    .Y(_25112_));
 sky130_fd_sc_hd__a22o_1 _28286_ (.A1(_25087_),
    .A2(_25088_),
    .B1(_25108_),
    .B2(_25111_),
    .X(_25113_));
 sky130_fd_sc_hd__and2_1 _28287_ (.A(_25112_),
    .B(_25113_),
    .X(_25114_));
 sky130_fd_sc_hd__xnor2_4 _28288_ (.A(_25076_),
    .B(_25114_),
    .Y(_25115_));
 sky130_fd_sc_hd__xor2_4 _28289_ (.A(_25065_),
    .B(_25115_),
    .X(_25116_));
 sky130_fd_sc_hd__xor2_4 _28290_ (.A(_25064_),
    .B(_25116_),
    .X(_25118_));
 sky130_fd_sc_hd__xnor2_1 _28291_ (.A(_25011_),
    .B(_25118_),
    .Y(_25119_));
 sky130_fd_sc_hd__nor2_1 _28292_ (.A(_24868_),
    .B(_25119_),
    .Y(_25120_));
 sky130_fd_sc_hd__a21boi_1 _28293_ (.A1(_23308_),
    .A2(_23427_),
    .B1_N(_23538_),
    .Y(_25121_));
 sky130_fd_sc_hd__a21o_1 _28294_ (.A1(_25119_),
    .A2(_24868_),
    .B1(_25121_),
    .X(_25122_));
 sky130_fd_sc_hd__o211a_1 _28295_ (.A1(_23300_),
    .A2(_23299_),
    .B1(_23298_),
    .C1(_25119_),
    .X(_25123_));
 sky130_fd_sc_hd__o21ai_1 _28296_ (.A1(_25120_),
    .A2(_25123_),
    .B1(_25121_),
    .Y(_25124_));
 sky130_fd_sc_hd__o21ai_1 _28297_ (.A1(_25120_),
    .A2(_25122_),
    .B1(_25124_),
    .Y(_25125_));
 sky130_fd_sc_hd__or2_1 _28298_ (.A(_24867_),
    .B(_25125_),
    .X(_25126_));
 sky130_fd_sc_hd__nand2_1 _28299_ (.A(_24867_),
    .B(_25125_),
    .Y(_25127_));
 sky130_fd_sc_hd__nand2_2 _28300_ (.A(_25126_),
    .B(_25127_),
    .Y(_25129_));
 sky130_fd_sc_hd__xor2_2 _28301_ (.A(_24309_),
    .B(_25129_),
    .X(_25130_));
 sky130_fd_sc_hd__a21oi_4 _28302_ (.A1(_24307_),
    .A2(_24308_),
    .B1(_25130_),
    .Y(_25131_));
 sky130_fd_sc_hd__nor2_1 _28303_ (.A(_22805_),
    .B(_23631_),
    .Y(_25132_));
 sky130_fd_sc_hd__a21oi_2 _28304_ (.A1(_24301_),
    .A2(_24305_),
    .B1(_24306_),
    .Y(_25133_));
 sky130_fd_sc_hd__nand2_1 _28305_ (.A(_24308_),
    .B(_25130_),
    .Y(_25134_));
 sky130_fd_sc_hd__o22ai_4 _28306_ (.A1(_23547_),
    .A2(_25132_),
    .B1(_25133_),
    .B2(_25134_),
    .Y(_25135_));
 sky130_fd_sc_hd__inv_2 _28307_ (.A(_22788_),
    .Y(_25136_));
 sky130_fd_sc_hd__o211a_1 _28308_ (.A1(_22793_),
    .A2(_25136_),
    .B1(_24301_),
    .C1(_24305_),
    .X(_25137_));
 sky130_fd_sc_hd__inv_2 _28309_ (.A(_25130_),
    .Y(_25138_));
 sky130_fd_sc_hd__o21ai_1 _28310_ (.A1(_25133_),
    .A2(_25137_),
    .B1(_25138_),
    .Y(_25140_));
 sky130_fd_sc_hd__a31oi_1 _28311_ (.A1(_24301_),
    .A2(_24305_),
    .A3(_24306_),
    .B1(_25138_),
    .Y(_25141_));
 sky130_fd_sc_hd__nand2_1 _28312_ (.A(_25141_),
    .B(_24307_),
    .Y(_25142_));
 sky130_fd_sc_hd__or2_1 _28313_ (.A(_23547_),
    .B(_25132_),
    .X(_25143_));
 sky130_fd_sc_hd__a21o_1 _28314_ (.A1(_25140_),
    .A2(_25142_),
    .B1(_25143_),
    .X(_25144_));
 sky130_fd_sc_hd__o221ai_2 _28315_ (.A1(_23743_),
    .A2(_23744_),
    .B1(_25131_),
    .B2(_25135_),
    .C1(_25144_),
    .Y(_25145_));
 sky130_fd_sc_hd__nand2_1 _28316_ (.A(_24307_),
    .B(_24308_),
    .Y(_25146_));
 sky130_fd_sc_hd__a21oi_1 _28317_ (.A1(_25146_),
    .A2(_25138_),
    .B1(_25135_),
    .Y(_25147_));
 sky130_fd_sc_hd__a21oi_2 _28318_ (.A1(_25140_),
    .A2(_25142_),
    .B1(_25143_),
    .Y(_25148_));
 sky130_fd_sc_hd__nor2_1 _28319_ (.A(_23743_),
    .B(_23744_),
    .Y(_25149_));
 sky130_fd_sc_hd__o21ai_1 _28320_ (.A1(_25147_),
    .A2(_25148_),
    .B1(_25149_),
    .Y(_25151_));
 sky130_fd_sc_hd__nand3b_2 _28321_ (.A_N(_23675_),
    .B(_25145_),
    .C(_25151_),
    .Y(_25152_));
 sky130_fd_sc_hd__nand2_1 _28322_ (.A(_23741_),
    .B(_23677_),
    .Y(_25153_));
 sky130_fd_sc_hd__or2b_2 _28323_ (.A(_23743_),
    .B_N(_25153_),
    .X(_25154_));
 sky130_fd_sc_hd__o21ai_1 _28324_ (.A1(_25147_),
    .A2(_25148_),
    .B1(_25154_),
    .Y(_25155_));
 sky130_fd_sc_hd__o211ai_1 _28325_ (.A1(_25131_),
    .A2(_25135_),
    .B1(_25149_),
    .C1(_25144_),
    .Y(_25156_));
 sky130_fd_sc_hd__nand3_2 _28326_ (.A(_23675_),
    .B(_25155_),
    .C(_25156_),
    .Y(_25157_));
 sky130_fd_sc_hd__nand3_1 _28327_ (.A(_23614_),
    .B(_23615_),
    .C(_23618_),
    .Y(_25158_));
 sky130_fd_sc_hd__clkbuf_2 _28328_ (.A(_23602_),
    .X(_25159_));
 sky130_fd_sc_hd__and2b_1 _28329_ (.A_N(_25159_),
    .B(_20964_),
    .X(_25160_));
 sky130_fd_sc_hd__o21a_1 _28330_ (.A1(_22194_),
    .A2(_20967_),
    .B1(_25160_),
    .X(_25162_));
 sky130_fd_sc_hd__nor2_1 _28331_ (.A(_19825_),
    .B(_00854_),
    .Y(_25163_));
 sky130_fd_sc_hd__and2_1 _28332_ (.A(_00843_),
    .B(_18811_),
    .X(_25164_));
 sky130_fd_sc_hd__or4_2 _28333_ (.A(_22139_),
    .B(_25163_),
    .C(_18722_),
    .D(_25164_),
    .X(_25165_));
 sky130_fd_sc_hd__a2bb2o_1 _28334_ (.A1_N(_25164_),
    .A2_N(_25163_),
    .B1(_04931_),
    .B2(_22177_),
    .X(_25166_));
 sky130_fd_sc_hd__nand2_1 _28335_ (.A(_25165_),
    .B(_25166_),
    .Y(_25167_));
 sky130_fd_sc_hd__xor2_2 _28336_ (.A(_25162_),
    .B(_25167_),
    .X(_25168_));
 sky130_fd_sc_hd__a21oi_2 _28337_ (.A1(_23601_),
    .A2(_23609_),
    .B1(_25168_),
    .Y(_25169_));
 sky130_fd_sc_hd__inv_2 _28338_ (.A(_25169_),
    .Y(_25170_));
 sky130_fd_sc_hd__nand3_1 _28339_ (.A(_23601_),
    .B(_23609_),
    .C(_25168_),
    .Y(_25171_));
 sky130_fd_sc_hd__and3_1 _28340_ (.A(_25170_),
    .B(net259),
    .C(_25171_),
    .X(_25173_));
 sky130_fd_sc_hd__a21oi_1 _28341_ (.A1(_25171_),
    .A2(_25170_),
    .B1(net259),
    .Y(_25174_));
 sky130_fd_sc_hd__o211a_1 _28342_ (.A1(_25173_),
    .A2(_25174_),
    .B1(_23643_),
    .C1(_23645_),
    .X(_25175_));
 sky130_fd_sc_hd__a211oi_1 _28343_ (.A1(_23643_),
    .A2(_23645_),
    .B1(_25173_),
    .C1(_25174_),
    .Y(_25176_));
 sky130_fd_sc_hd__or2_1 _28344_ (.A(_25175_),
    .B(_25176_),
    .X(_25177_));
 sky130_fd_sc_hd__a21oi_1 _28345_ (.A1(_23614_),
    .A2(_25158_),
    .B1(_25177_),
    .Y(_25178_));
 sky130_fd_sc_hd__nand3_1 _28346_ (.A(_23614_),
    .B(_25158_),
    .C(_25177_),
    .Y(_25179_));
 sky130_fd_sc_hd__and2b_1 _28347_ (.A_N(_25178_),
    .B(_25179_),
    .X(_25180_));
 sky130_fd_sc_hd__xor2_1 _28348_ (.A(_23647_),
    .B(_25180_),
    .X(_25181_));
 sky130_fd_sc_hd__a21o_1 _28349_ (.A1(_25152_),
    .A2(_25157_),
    .B1(_25181_),
    .X(_25182_));
 sky130_fd_sc_hd__nand3_1 _28350_ (.A(_25152_),
    .B(_25181_),
    .C(_25157_),
    .Y(_25184_));
 sky130_fd_sc_hd__nand3_1 _28351_ (.A(_23674_),
    .B(_25182_),
    .C(_25184_),
    .Y(_25185_));
 sky130_fd_sc_hd__xnor2_1 _28352_ (.A(_23647_),
    .B(_25180_),
    .Y(_25186_));
 sky130_fd_sc_hd__a21o_1 _28353_ (.A1(_25152_),
    .A2(_25157_),
    .B1(_25186_),
    .X(_25187_));
 sky130_fd_sc_hd__and2_1 _28354_ (.A(_23628_),
    .B(_23673_),
    .X(_25188_));
 sky130_fd_sc_hd__nand3_1 _28355_ (.A(_25152_),
    .B(_25157_),
    .C(_25186_),
    .Y(_25189_));
 sky130_fd_sc_hd__nand3_2 _28356_ (.A(_25187_),
    .B(_25188_),
    .C(_25189_),
    .Y(_25190_));
 sky130_fd_sc_hd__or3_1 _28357_ (.A(_23636_),
    .B(_23647_),
    .C(_23648_),
    .X(_25191_));
 sky130_fd_sc_hd__o21ai_2 _28358_ (.A1(_22187_),
    .A2(_23650_),
    .B1(_25191_),
    .Y(_25192_));
 sky130_fd_sc_hd__a21oi_1 _28359_ (.A1(_25185_),
    .A2(_25190_),
    .B1(_25192_),
    .Y(_25193_));
 sky130_fd_sc_hd__inv_2 _28360_ (.A(_25192_),
    .Y(_25195_));
 sky130_fd_sc_hd__nand2_1 _28361_ (.A(_25185_),
    .B(_25190_),
    .Y(_25196_));
 sky130_fd_sc_hd__a32o_1 _28362_ (.A1(_23656_),
    .A2(_23658_),
    .A3(_23659_),
    .B1(_23657_),
    .B2(_23663_),
    .X(_25197_));
 sky130_fd_sc_hd__o21ai_1 _28363_ (.A1(_25195_),
    .A2(_25196_),
    .B1(_25197_),
    .Y(_25198_));
 sky130_fd_sc_hd__a21o_1 _28364_ (.A1(_25185_),
    .A2(_25190_),
    .B1(_25195_),
    .X(_25199_));
 sky130_fd_sc_hd__inv_2 _28365_ (.A(_25197_),
    .Y(_25200_));
 sky130_fd_sc_hd__o2111ai_1 _28366_ (.A1(_22187_),
    .A2(_23650_),
    .B1(_25185_),
    .C1(_25190_),
    .D1(_25191_),
    .Y(_25201_));
 sky130_fd_sc_hd__nand3_1 _28367_ (.A(_25199_),
    .B(_25200_),
    .C(_25201_),
    .Y(_25202_));
 sky130_fd_sc_hd__o21ai_2 _28368_ (.A1(_25193_),
    .A2(_25198_),
    .B1(_25202_),
    .Y(_25203_));
 sky130_fd_sc_hd__xnor2_2 _28369_ (.A(_23672_),
    .B(_25203_),
    .Y(_00004_));
 sky130_fd_sc_hd__a2bb2oi_2 _28370_ (.A1_N(_25193_),
    .A2_N(_25198_),
    .B1(_25202_),
    .B2(_23672_),
    .Y(_25205_));
 sky130_fd_sc_hd__o22a_1 _28371_ (.A1(_25131_),
    .A2(_25135_),
    .B1(_25154_),
    .B2(_25148_),
    .X(_25206_));
 sky130_fd_sc_hd__buf_1 _28372_ (.A(_24274_),
    .X(_25207_));
 sky130_fd_sc_hd__nand2_1 _28373_ (.A(_24299_),
    .B(_24293_),
    .Y(_25208_));
 sky130_fd_sc_hd__o221a_1 _28374_ (.A1(_23539_),
    .A2(_24295_),
    .B1(_25207_),
    .B2(_25208_),
    .C1(_24304_),
    .X(_25209_));
 sky130_fd_sc_hd__inv_2 _28375_ (.A(_24306_),
    .Y(_25210_));
 sky130_fd_sc_hd__a31oi_1 _28376_ (.A1(_24294_),
    .A2(_24296_),
    .A3(_24300_),
    .B1(_25210_),
    .Y(_25211_));
 sky130_fd_sc_hd__a21bo_1 _28377_ (.A1(_23571_),
    .A2(_23697_),
    .B1_N(_23696_),
    .X(_25212_));
 sky130_fd_sc_hd__or3_1 _28378_ (.A(_24280_),
    .B(_24289_),
    .C(_24290_),
    .X(_25213_));
 sky130_fd_sc_hd__or3b_1 _28379_ (.A(_23683_),
    .B(_23684_),
    .C_N(_23560_),
    .X(_25214_));
 sky130_fd_sc_hd__buf_1 _28380_ (.A(_23682_),
    .X(_25216_));
 sky130_fd_sc_hd__clkbuf_2 _28381_ (.A(\delay_line[20][11] ),
    .X(_25217_));
 sky130_fd_sc_hd__nor2_1 _28382_ (.A(_23682_),
    .B(_25217_),
    .Y(_25218_));
 sky130_fd_sc_hd__and2_1 _28383_ (.A(\delay_line[20][10] ),
    .B(_25217_),
    .X(_25219_));
 sky130_fd_sc_hd__nor2_2 _28384_ (.A(_25218_),
    .B(_25219_),
    .Y(_25220_));
 sky130_fd_sc_hd__and3_1 _28385_ (.A(_23681_),
    .B(_25216_),
    .C(_25220_),
    .X(_25221_));
 sky130_fd_sc_hd__o2bb2a_1 _28386_ (.A1_N(_23681_),
    .A2_N(_25216_),
    .B1(_25218_),
    .B2(_25219_),
    .X(_25222_));
 sky130_fd_sc_hd__xnor2_1 _28387_ (.A(_19795_),
    .B(_23561_),
    .Y(_25223_));
 sky130_fd_sc_hd__clkbuf_2 _28388_ (.A(_25223_),
    .X(_25224_));
 sky130_fd_sc_hd__nor3_2 _28389_ (.A(_25221_),
    .B(_25222_),
    .C(_25224_),
    .Y(_25225_));
 sky130_fd_sc_hd__o21a_1 _28390_ (.A1(_25221_),
    .A2(_25222_),
    .B1(_25224_),
    .X(_25227_));
 sky130_fd_sc_hd__a211oi_2 _28391_ (.A1(_25214_),
    .A2(_23690_),
    .B1(_25225_),
    .C1(_25227_),
    .Y(_25228_));
 sky130_fd_sc_hd__o221a_1 _28392_ (.A1(_23688_),
    .A2(_23691_),
    .B1(_25227_),
    .B2(_25225_),
    .C1(_25214_),
    .X(_25229_));
 sky130_fd_sc_hd__a211o_1 _28393_ (.A1(_24285_),
    .A2(_25213_),
    .B1(_25228_),
    .C1(_25229_),
    .X(_25230_));
 sky130_fd_sc_hd__o211ai_2 _28394_ (.A1(_25228_),
    .A2(_25229_),
    .B1(_24285_),
    .C1(_25213_),
    .Y(_25231_));
 sky130_fd_sc_hd__and3_1 _28395_ (.A(_25230_),
    .B(_25231_),
    .C(_23694_),
    .X(_25232_));
 sky130_fd_sc_hd__a21oi_1 _28396_ (.A1(_25230_),
    .A2(_25231_),
    .B1(_23694_),
    .Y(_25233_));
 sky130_fd_sc_hd__nor2_1 _28397_ (.A(_25232_),
    .B(_25233_),
    .Y(_25234_));
 sky130_fd_sc_hd__xnor2_1 _28398_ (.A(_25212_),
    .B(_25234_),
    .Y(_25235_));
 sky130_fd_sc_hd__buf_1 _28399_ (.A(_23719_),
    .X(_25236_));
 sky130_fd_sc_hd__buf_2 _28400_ (.A(_23592_),
    .X(_25238_));
 sky130_fd_sc_hd__o211a_1 _28401_ (.A1(_25236_),
    .A2(_25238_),
    .B1(_19819_),
    .C1(_10767_),
    .X(_25239_));
 sky130_fd_sc_hd__clkbuf_2 _28402_ (.A(_23719_),
    .X(_25240_));
 sky130_fd_sc_hd__a211oi_2 _28403_ (.A1(_10767_),
    .A2(_19819_),
    .B1(_25238_),
    .C1(_25240_),
    .Y(_25241_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28404_ (.A(net376),
    .X(_25242_));
 sky130_fd_sc_hd__nand2_1 _28405_ (.A(_25159_),
    .B(_25242_),
    .Y(_25243_));
 sky130_fd_sc_hd__o31a_1 _28406_ (.A1(_23726_),
    .A2(_25239_),
    .A3(_25241_),
    .B1(_25243_),
    .X(_25244_));
 sky130_fd_sc_hd__nor4_2 _28407_ (.A(_25243_),
    .B(_25239_),
    .C(_25241_),
    .D(_23726_),
    .Y(_25245_));
 sky130_fd_sc_hd__or2_2 _28408_ (.A(_25244_),
    .B(_25245_),
    .X(_25246_));
 sky130_fd_sc_hd__or2_2 _28409_ (.A(\delay_line[17][10] ),
    .B(\delay_line[17][11] ),
    .X(_25247_));
 sky130_fd_sc_hd__buf_1 _28410_ (.A(\delay_line[17][11] ),
    .X(_25249_));
 sky130_fd_sc_hd__nand2_1 _28411_ (.A(_23719_),
    .B(_25249_),
    .Y(_25250_));
 sky130_fd_sc_hd__buf_2 _28412_ (.A(_25250_),
    .X(_25251_));
 sky130_fd_sc_hd__nor2_1 _28413_ (.A(_18744_),
    .B(_10954_),
    .Y(_25252_));
 sky130_fd_sc_hd__and3b_1 _28414_ (.A_N(_04821_),
    .B(_04843_),
    .C(_18744_),
    .X(_25253_));
 sky130_fd_sc_hd__o2bb2a_1 _28415_ (.A1_N(_25247_),
    .A2_N(_25251_),
    .B1(_25252_),
    .B2(_25253_),
    .X(_25254_));
 sky130_fd_sc_hd__nand2_1 _28416_ (.A(_10954_),
    .B(_18744_),
    .Y(_25255_));
 sky130_fd_sc_hd__and2_1 _28417_ (.A(_25247_),
    .B(_25250_),
    .X(_25256_));
 sky130_fd_sc_hd__and3b_1 _28418_ (.A_N(_25252_),
    .B(_25255_),
    .C(_25256_),
    .X(_25257_));
 sky130_fd_sc_hd__nor2_1 _28419_ (.A(_25254_),
    .B(_25257_),
    .Y(_25258_));
 sky130_fd_sc_hd__a21oi_2 _28420_ (.A1(_19790_),
    .A2(_23555_),
    .B1(_20929_),
    .Y(_25260_));
 sky130_fd_sc_hd__and2_1 _28421_ (.A(_20928_),
    .B(_25260_),
    .X(_25261_));
 sky130_fd_sc_hd__nor2_1 _28422_ (.A(_25260_),
    .B(_20928_),
    .Y(_25262_));
 sky130_fd_sc_hd__or3_1 _28423_ (.A(_20947_),
    .B(_25261_),
    .C(_25262_),
    .X(_25263_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28424_ (.A(_20947_),
    .X(_25264_));
 sky130_fd_sc_hd__o21ai_1 _28425_ (.A1(_25261_),
    .A2(_25262_),
    .B1(_25264_),
    .Y(_25265_));
 sky130_fd_sc_hd__a211oi_1 _28426_ (.A1(_25263_),
    .A2(_25265_),
    .B1(_23708_),
    .C1(_23711_),
    .Y(_25266_));
 sky130_fd_sc_hd__o211a_1 _28427_ (.A1(_23708_),
    .A2(_23711_),
    .B1(_25263_),
    .C1(_25265_),
    .X(_25267_));
 sky130_fd_sc_hd__nor2_1 _28428_ (.A(_25266_),
    .B(_25267_),
    .Y(_25268_));
 sky130_fd_sc_hd__or2_2 _28429_ (.A(_25258_),
    .B(_25268_),
    .X(_25269_));
 sky130_fd_sc_hd__or3b_2 _28430_ (.A(_25266_),
    .B(_25267_),
    .C_N(_25258_),
    .X(_25271_));
 sky130_fd_sc_hd__a221oi_4 _28431_ (.A1(_23713_),
    .A2(_23714_),
    .B1(_25269_),
    .B2(_25271_),
    .C1(_23729_),
    .Y(_25272_));
 sky130_fd_sc_hd__o211ai_4 _28432_ (.A1(_23716_),
    .A2(_23729_),
    .B1(_25271_),
    .C1(_25269_),
    .Y(_25273_));
 sky130_fd_sc_hd__or2b_1 _28433_ (.A(_25272_),
    .B_N(_25273_),
    .X(_25274_));
 sky130_fd_sc_hd__xor2_2 _28434_ (.A(_25246_),
    .B(_25274_),
    .X(_25275_));
 sky130_fd_sc_hd__xor2_1 _28435_ (.A(_25235_),
    .B(_25275_),
    .X(_25276_));
 sky130_fd_sc_hd__o21bai_2 _28436_ (.A1(_25209_),
    .A2(_25211_),
    .B1_N(_25276_),
    .Y(_25277_));
 sky130_fd_sc_hd__o21ai_1 _28437_ (.A1(_25207_),
    .A2(_25208_),
    .B1(_24304_),
    .Y(_25278_));
 sky130_fd_sc_hd__a31o_1 _28438_ (.A1(_24294_),
    .A2(_24296_),
    .A3(_24300_),
    .B1(_25210_),
    .X(_25279_));
 sky130_fd_sc_hd__o211ai_2 _28439_ (.A1(_24296_),
    .A2(_25278_),
    .B1(_25276_),
    .C1(_25279_),
    .Y(_25280_));
 sky130_fd_sc_hd__o21bai_2 _28440_ (.A1(_23702_),
    .A2(_23736_),
    .B1_N(_23701_),
    .Y(_25282_));
 sky130_fd_sc_hd__a21o_1 _28441_ (.A1(_25277_),
    .A2(_25280_),
    .B1(_25282_),
    .X(_25283_));
 sky130_fd_sc_hd__nand3_1 _28442_ (.A(_25282_),
    .B(_25277_),
    .C(_25280_),
    .Y(_25284_));
 sky130_fd_sc_hd__nand2_1 _28443_ (.A(_25283_),
    .B(_25284_),
    .Y(_25285_));
 sky130_fd_sc_hd__o22ai_1 _28444_ (.A1(_25129_),
    .A2(_24309_),
    .B1(_25133_),
    .B2(_25134_),
    .Y(_25286_));
 sky130_fd_sc_hd__o21ba_1 _28445_ (.A1(_25121_),
    .A2(_25123_),
    .B1_N(_25120_),
    .X(_25287_));
 sky130_fd_sc_hd__nand2_1 _28446_ (.A(_24263_),
    .B(_24272_),
    .Y(_25288_));
 sky130_fd_sc_hd__or2b_1 _28447_ (.A(_25065_),
    .B_N(_25115_),
    .X(_25289_));
 sky130_fd_sc_hd__o21ai_2 _28448_ (.A1(_25064_),
    .A2(_25116_),
    .B1(_25289_),
    .Y(_25290_));
 sky130_fd_sc_hd__inv_2 _28449_ (.A(_25290_),
    .Y(_25291_));
 sky130_fd_sc_hd__inv_2 _28450_ (.A(_25060_),
    .Y(_25293_));
 sky130_fd_sc_hd__or2_1 _28451_ (.A(_23966_),
    .B(_23993_),
    .X(_25294_));
 sky130_fd_sc_hd__nand2_1 _28452_ (.A(_23952_),
    .B(_23954_),
    .Y(_25295_));
 sky130_fd_sc_hd__clkbuf_2 _28453_ (.A(\delay_line[7][11] ),
    .X(_25296_));
 sky130_fd_sc_hd__clkbuf_2 _28454_ (.A(_25296_),
    .X(_25297_));
 sky130_fd_sc_hd__nand2_1 _28455_ (.A(_18844_),
    .B(_25297_),
    .Y(_25298_));
 sky130_fd_sc_hd__or2_1 _28456_ (.A(_25296_),
    .B(_18844_),
    .X(_25299_));
 sky130_fd_sc_hd__or4bb_1 _28457_ (.A(_09009_),
    .B(_11866_),
    .C_N(_25298_),
    .D_N(_25299_),
    .X(_25300_));
 sky130_fd_sc_hd__a2bb2o_1 _28458_ (.A1_N(_11899_),
    .A2_N(_11866_),
    .B1(_25298_),
    .B2(_25299_),
    .X(_25301_));
 sky130_fd_sc_hd__nand2_1 _28459_ (.A(_25300_),
    .B(_25301_),
    .Y(_25302_));
 sky130_fd_sc_hd__a21oi_1 _28460_ (.A1(_23950_),
    .A2(_25295_),
    .B1(_25302_),
    .Y(_25304_));
 sky130_fd_sc_hd__and3_1 _28461_ (.A(_23950_),
    .B(_25302_),
    .C(_25295_),
    .X(_25305_));
 sky130_fd_sc_hd__nor2_1 _28462_ (.A(_25304_),
    .B(_25305_),
    .Y(_25306_));
 sky130_fd_sc_hd__xnor2_1 _28463_ (.A(_23933_),
    .B(_25306_),
    .Y(_25307_));
 sky130_fd_sc_hd__buf_1 _28464_ (.A(\delay_line[8][11] ),
    .X(_25308_));
 sky130_fd_sc_hd__nor2b_1 _28465_ (.A(_08657_),
    .B_N(_25308_),
    .Y(_25309_));
 sky130_fd_sc_hd__buf_1 _28466_ (.A(_25309_),
    .X(_25310_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28467_ (.A(_25308_),
    .X(_25311_));
 sky130_fd_sc_hd__and2b_1 _28468_ (.A_N(_25311_),
    .B(_18053_),
    .X(_25312_));
 sky130_fd_sc_hd__clkbuf_2 _28469_ (.A(\delay_line[8][9] ),
    .X(_25313_));
 sky130_fd_sc_hd__and3b_1 _28470_ (.A_N(_02876_),
    .B(_18055_),
    .C(_25313_),
    .X(_25315_));
 sky130_fd_sc_hd__o22ai_1 _28471_ (.A1(_25310_),
    .A2(_25312_),
    .B1(_25315_),
    .B2(_18054_),
    .Y(_25316_));
 sky130_fd_sc_hd__or4_1 _28472_ (.A(_18054_),
    .B(_25310_),
    .C(_25312_),
    .D(_25315_),
    .X(_25317_));
 sky130_fd_sc_hd__or3_1 _28473_ (.A(_21869_),
    .B(_22503_),
    .C(_23943_),
    .X(_25318_));
 sky130_fd_sc_hd__and3_1 _28474_ (.A(_25318_),
    .B(_18044_),
    .C(_23948_),
    .X(_25319_));
 sky130_fd_sc_hd__a21oi_1 _28475_ (.A1(_23948_),
    .A2(_25318_),
    .B1(_18044_),
    .Y(_25320_));
 sky130_fd_sc_hd__or2_1 _28476_ (.A(_25319_),
    .B(_25320_),
    .X(_25321_));
 sky130_fd_sc_hd__and3_1 _28477_ (.A(_25316_),
    .B(_25317_),
    .C(_25321_),
    .X(_25322_));
 sky130_fd_sc_hd__a21oi_1 _28478_ (.A1(_25316_),
    .A2(_25317_),
    .B1(_25321_),
    .Y(_25323_));
 sky130_fd_sc_hd__nor2_1 _28479_ (.A(_25322_),
    .B(_25323_),
    .Y(_25324_));
 sky130_fd_sc_hd__a32o_1 _28480_ (.A1(_23956_),
    .A2(_23959_),
    .A3(_23955_),
    .B1(_23957_),
    .B2(_18058_),
    .X(_25326_));
 sky130_fd_sc_hd__and2_1 _28481_ (.A(_25324_),
    .B(_25326_),
    .X(_25327_));
 sky130_fd_sc_hd__nor2_1 _28482_ (.A(_25326_),
    .B(_25324_),
    .Y(_25328_));
 sky130_fd_sc_hd__or2_1 _28483_ (.A(_25327_),
    .B(_25328_),
    .X(_25329_));
 sky130_fd_sc_hd__nor2_1 _28484_ (.A(_25307_),
    .B(_25329_),
    .Y(_25330_));
 sky130_fd_sc_hd__nand2_1 _28485_ (.A(_25307_),
    .B(_25329_),
    .Y(_25331_));
 sky130_fd_sc_hd__or2b_1 _28486_ (.A(_25330_),
    .B_N(_25331_),
    .X(_25332_));
 sky130_fd_sc_hd__a21bo_1 _28487_ (.A1(_23968_),
    .A2(_23987_),
    .B1_N(_23989_),
    .X(_25333_));
 sky130_fd_sc_hd__a31o_1 _28488_ (.A1(_23980_),
    .A2(_23977_),
    .A3(_23979_),
    .B1(_23986_),
    .X(_25334_));
 sky130_fd_sc_hd__o21ai_1 _28489_ (.A1(_23757_),
    .A2(_23767_),
    .B1(_23765_),
    .Y(_25335_));
 sky130_fd_sc_hd__buf_2 _28490_ (.A(_22440_),
    .X(_25337_));
 sky130_fd_sc_hd__and3_1 _28491_ (.A(_23976_),
    .B(_25337_),
    .C(_23969_),
    .X(_25338_));
 sky130_fd_sc_hd__nand2_2 _28492_ (.A(_23974_),
    .B(_23971_),
    .Y(_25339_));
 sky130_fd_sc_hd__a211oi_1 _28493_ (.A1(_25339_),
    .A2(_22439_),
    .B1(_17915_),
    .C1(_23978_),
    .Y(_25340_));
 sky130_fd_sc_hd__buf_2 _28494_ (.A(\delay_line[9][10] ),
    .X(_25341_));
 sky130_fd_sc_hd__a21oi_1 _28495_ (.A1(_23974_),
    .A2(_25341_),
    .B1(_23970_),
    .Y(_25342_));
 sky130_fd_sc_hd__o21a_1 _28496_ (.A1(_23972_),
    .A2(_25342_),
    .B1(_17915_),
    .X(_25343_));
 sky130_fd_sc_hd__or2_1 _28497_ (.A(_25340_),
    .B(_25343_),
    .X(_25344_));
 sky130_fd_sc_hd__nand2_1 _28498_ (.A(_23752_),
    .B(_23754_),
    .Y(_25345_));
 sky130_fd_sc_hd__xnor2_1 _28499_ (.A(_25344_),
    .B(_25345_),
    .Y(_25346_));
 sky130_fd_sc_hd__xnor2_1 _28500_ (.A(_25338_),
    .B(_25346_),
    .Y(_25348_));
 sky130_fd_sc_hd__or2_1 _28501_ (.A(_25335_),
    .B(_25348_),
    .X(_25349_));
 sky130_fd_sc_hd__nand2_1 _28502_ (.A(_25348_),
    .B(_25335_),
    .Y(_25350_));
 sky130_fd_sc_hd__nand2_1 _28503_ (.A(_25349_),
    .B(_25350_),
    .Y(_25351_));
 sky130_fd_sc_hd__xnor2_1 _28504_ (.A(_25334_),
    .B(_25351_),
    .Y(_25352_));
 sky130_fd_sc_hd__or2_1 _28505_ (.A(_25333_),
    .B(_25352_),
    .X(_25353_));
 sky130_fd_sc_hd__nand2_1 _28506_ (.A(_25352_),
    .B(_25333_),
    .Y(_25354_));
 sky130_fd_sc_hd__nand2_1 _28507_ (.A(_25353_),
    .B(_25354_),
    .Y(_25355_));
 sky130_fd_sc_hd__or2_2 _28508_ (.A(_25332_),
    .B(_25355_),
    .X(_25356_));
 sky130_fd_sc_hd__nand2_1 _28509_ (.A(_25332_),
    .B(_25355_),
    .Y(_25357_));
 sky130_fd_sc_hd__a21boi_1 _28510_ (.A1(_23782_),
    .A2(_23783_),
    .B1_N(_23785_),
    .Y(_25359_));
 sky130_fd_sc_hd__a21boi_2 _28511_ (.A1(_25356_),
    .A2(_25357_),
    .B1_N(_25359_),
    .Y(_25360_));
 sky130_fd_sc_hd__nand3b_2 _28512_ (.A_N(_25359_),
    .B(_25356_),
    .C(_25357_),
    .Y(_25361_));
 sky130_fd_sc_hd__or2b_2 _28513_ (.A(_25360_),
    .B_N(_25361_),
    .X(_25362_));
 sky130_fd_sc_hd__o211a_2 _28514_ (.A1(_23991_),
    .A2(_23992_),
    .B1(_25294_),
    .C1(_25362_),
    .X(_25363_));
 sky130_fd_sc_hd__o21a_2 _28515_ (.A1(_23991_),
    .A2(_23992_),
    .B1(_25294_),
    .X(_25364_));
 sky130_fd_sc_hd__nor2_2 _28516_ (.A(_25364_),
    .B(_25362_),
    .Y(_25365_));
 sky130_fd_sc_hd__a211oi_2 _28517_ (.A1(_22464_),
    .A2(_22471_),
    .B1(_23777_),
    .C1(_23778_),
    .Y(_25366_));
 sky130_fd_sc_hd__nor2_1 _28518_ (.A(_23768_),
    .B(_23781_),
    .Y(_25367_));
 sky130_fd_sc_hd__a31o_1 _28519_ (.A1(_23802_),
    .A2(_23803_),
    .A3(_23805_),
    .B1(_23807_),
    .X(_25368_));
 sky130_fd_sc_hd__clkbuf_2 _28520_ (.A(\delay_line[10][11] ),
    .X(_25370_));
 sky130_fd_sc_hd__and3_1 _28521_ (.A(_12174_),
    .B(_18987_),
    .C(_25370_),
    .X(_25371_));
 sky130_fd_sc_hd__clkbuf_2 _28522_ (.A(_22392_),
    .X(_25372_));
 sky130_fd_sc_hd__clkbuf_2 _28523_ (.A(_23798_),
    .X(_25373_));
 sky130_fd_sc_hd__nand2_1 _28524_ (.A(_25372_),
    .B(_25373_),
    .Y(_25374_));
 sky130_fd_sc_hd__clkbuf_2 _28525_ (.A(\delay_line[10][11] ),
    .X(_25375_));
 sky130_fd_sc_hd__clkbuf_2 _28526_ (.A(_25375_),
    .X(_25376_));
 sky130_fd_sc_hd__a21oi_1 _28527_ (.A1(_12174_),
    .A2(_18988_),
    .B1(_25376_),
    .Y(_25377_));
 sky130_fd_sc_hd__nor4_1 _28528_ (.A(_23795_),
    .B(_25371_),
    .C(_25374_),
    .D(_25377_),
    .Y(_25378_));
 sky130_fd_sc_hd__o22a_1 _28529_ (.A1(_25374_),
    .A2(_23795_),
    .B1(_25371_),
    .B2(_25377_),
    .X(_25379_));
 sky130_fd_sc_hd__nor2_1 _28530_ (.A(_25378_),
    .B(_25379_),
    .Y(_25381_));
 sky130_fd_sc_hd__xnor2_1 _28531_ (.A(_23770_),
    .B(_25381_),
    .Y(_25382_));
 sky130_fd_sc_hd__or2_1 _28532_ (.A(_23776_),
    .B(_23777_),
    .X(_25383_));
 sky130_fd_sc_hd__xor2_1 _28533_ (.A(_25382_),
    .B(_25383_),
    .X(_25384_));
 sky130_fd_sc_hd__nor2_1 _28534_ (.A(_17921_),
    .B(_22448_),
    .Y(_25385_));
 sky130_fd_sc_hd__and2_1 _28535_ (.A(_17919_),
    .B(_22447_),
    .X(_25386_));
 sky130_fd_sc_hd__or3b_2 _28536_ (.A(_25385_),
    .B(_25386_),
    .C_N(_21801_),
    .X(_25387_));
 sky130_fd_sc_hd__o21bai_1 _28537_ (.A1(_25385_),
    .A2(_25386_),
    .B1_N(_22458_),
    .Y(_25388_));
 sky130_fd_sc_hd__nand3b_2 _28538_ (.A_N(_23761_),
    .B(_25387_),
    .C(_25388_),
    .Y(_25389_));
 sky130_fd_sc_hd__a21bo_1 _28539_ (.A1(_25387_),
    .A2(_25388_),
    .B1_N(_23761_),
    .X(_25390_));
 sky130_fd_sc_hd__clkbuf_2 _28540_ (.A(net412),
    .X(_25392_));
 sky130_fd_sc_hd__or2b_2 _28541_ (.A(_21817_),
    .B_N(net418),
    .X(_25393_));
 sky130_fd_sc_hd__or2b_1 _28542_ (.A(net418),
    .B_N(_21817_),
    .X(_25394_));
 sky130_fd_sc_hd__a22o_1 _28543_ (.A1(_17919_),
    .A2(_25392_),
    .B1(_25393_),
    .B2(_25394_),
    .X(_25395_));
 sky130_fd_sc_hd__clkbuf_2 _28544_ (.A(net413),
    .X(_25396_));
 sky130_fd_sc_hd__nand4_4 _28545_ (.A(_25393_),
    .B(_25394_),
    .C(_17921_),
    .D(_21821_),
    .Y(_25397_));
 sky130_fd_sc_hd__nand4_4 _28546_ (.A(_17910_),
    .B(_25395_),
    .C(_25396_),
    .D(_25397_),
    .Y(_25398_));
 sky130_fd_sc_hd__a22o_1 _28547_ (.A1(_25396_),
    .A2(_17910_),
    .B1(_25395_),
    .B2(_25397_),
    .X(_25399_));
 sky130_fd_sc_hd__a22o_1 _28548_ (.A1(_25389_),
    .A2(_25390_),
    .B1(_25398_),
    .B2(_25399_),
    .X(_25400_));
 sky130_fd_sc_hd__nand4_4 _28549_ (.A(_25389_),
    .B(_25390_),
    .C(_25398_),
    .D(_25399_),
    .Y(_25401_));
 sky130_fd_sc_hd__nand3_1 _28550_ (.A(_25384_),
    .B(_25400_),
    .C(_25401_),
    .Y(_25403_));
 sky130_fd_sc_hd__a21o_1 _28551_ (.A1(_25401_),
    .A2(_25400_),
    .B1(_25384_),
    .X(_25404_));
 sky130_fd_sc_hd__and2_1 _28552_ (.A(_25403_),
    .B(_25404_),
    .X(_25405_));
 sky130_fd_sc_hd__xnor2_1 _28553_ (.A(_25368_),
    .B(_25405_),
    .Y(_25406_));
 sky130_fd_sc_hd__nor3_1 _28554_ (.A(_25366_),
    .B(_25367_),
    .C(_25406_),
    .Y(_25407_));
 sky130_fd_sc_hd__o21a_1 _28555_ (.A1(_25366_),
    .A2(_25367_),
    .B1(_25406_),
    .X(_25408_));
 sky130_fd_sc_hd__nand3_2 _28556_ (.A(_22330_),
    .B(_22288_),
    .C(_22290_),
    .Y(_25409_));
 sky130_fd_sc_hd__o22a_2 _28557_ (.A1(_22294_),
    .A2(_22295_),
    .B1(_23832_),
    .B2(_23834_),
    .X(_25410_));
 sky130_fd_sc_hd__nand2_2 _28558_ (.A(_25409_),
    .B(_25410_),
    .Y(_25411_));
 sky130_fd_sc_hd__nor2_2 _28559_ (.A(_19993_),
    .B(_23833_),
    .Y(_25412_));
 sky130_fd_sc_hd__or3b_2 _28560_ (.A(_25412_),
    .B(_23831_),
    .C_N(_23827_),
    .X(_25414_));
 sky130_fd_sc_hd__o21a_2 _28561_ (.A1(_23826_),
    .A2(_23835_),
    .B1(_25414_),
    .X(_25415_));
 sky130_fd_sc_hd__clkbuf_2 _28562_ (.A(\delay_line[4][8] ),
    .X(_25416_));
 sky130_fd_sc_hd__nand2_1 _28563_ (.A(_23833_),
    .B(_25416_),
    .Y(_25417_));
 sky130_fd_sc_hd__or2b_2 _28564_ (.A(\delay_line[4][8] ),
    .B_N(\delay_line[4][6] ),
    .X(_25418_));
 sky130_fd_sc_hd__nor2b_4 _28565_ (.A(_22280_),
    .B_N(_23827_),
    .Y(_25419_));
 sky130_fd_sc_hd__a21oi_2 _28566_ (.A1(_25412_),
    .A2(_23829_),
    .B1(_25419_),
    .Y(_25420_));
 sky130_fd_sc_hd__a21oi_4 _28567_ (.A1(_25417_),
    .A2(_25418_),
    .B1(_25420_),
    .Y(_25421_));
 sky130_fd_sc_hd__and3_2 _28568_ (.A(_25420_),
    .B(_25418_),
    .C(_25417_),
    .X(_25422_));
 sky130_fd_sc_hd__nor2_2 _28569_ (.A(_25421_),
    .B(_25422_),
    .Y(_25423_));
 sky130_fd_sc_hd__nand3_4 _28570_ (.A(_25411_),
    .B(_25415_),
    .C(_25423_),
    .Y(_25425_));
 sky130_fd_sc_hd__o21ai_4 _28571_ (.A1(_23826_),
    .A2(_23835_),
    .B1(_25414_),
    .Y(_25426_));
 sky130_fd_sc_hd__o22ai_2 _28572_ (.A1(_22294_),
    .A2(_22295_),
    .B1(_23832_),
    .B2(_23834_),
    .Y(_25427_));
 sky130_fd_sc_hd__a21oi_4 _28573_ (.A1(_22328_),
    .A2(_22330_),
    .B1(_25427_),
    .Y(_25428_));
 sky130_fd_sc_hd__o22ai_4 _28574_ (.A1(_25421_),
    .A2(_25422_),
    .B1(_25426_),
    .B2(_25428_),
    .Y(_25429_));
 sky130_fd_sc_hd__nor2b_2 _28575_ (.A(_23839_),
    .B_N(_20002_),
    .Y(_25430_));
 sky130_fd_sc_hd__clkbuf_2 _28576_ (.A(_23842_),
    .X(_25431_));
 sky130_fd_sc_hd__o21ai_1 _28577_ (.A1(_25430_),
    .A2(_22309_),
    .B1(_25431_),
    .Y(_25432_));
 sky130_fd_sc_hd__buf_2 _28578_ (.A(\delay_line[11][9] ),
    .X(_25433_));
 sky130_fd_sc_hd__nand2b_1 _28579_ (.A_N(_20003_),
    .B(_25433_),
    .Y(_25434_));
 sky130_fd_sc_hd__nand2b_1 _28580_ (.A_N(\delay_line[11][9] ),
    .B(_20003_),
    .Y(_25436_));
 sky130_fd_sc_hd__nand2_2 _28581_ (.A(_25434_),
    .B(_25436_),
    .Y(_25437_));
 sky130_fd_sc_hd__nand2_1 _28582_ (.A(_25432_),
    .B(_25437_),
    .Y(_25438_));
 sky130_fd_sc_hd__xnor2_2 _28583_ (.A(_20003_),
    .B(_25433_),
    .Y(_25439_));
 sky130_fd_sc_hd__o211ai_2 _28584_ (.A1(_22313_),
    .A2(_25430_),
    .B1(_25431_),
    .C1(_25439_),
    .Y(_25440_));
 sky130_fd_sc_hd__nand2_1 _28585_ (.A(_25438_),
    .B(_25440_),
    .Y(_25441_));
 sky130_fd_sc_hd__o2bb2ai_1 _28586_ (.A1_N(_23846_),
    .A2_N(_23849_),
    .B1(_22311_),
    .B2(_23843_),
    .Y(_25442_));
 sky130_fd_sc_hd__nand2_2 _28587_ (.A(_25441_),
    .B(_25442_),
    .Y(_25443_));
 sky130_fd_sc_hd__and4b_1 _28588_ (.A_N(_23838_),
    .B(_23840_),
    .C(_25431_),
    .D(_22313_),
    .X(_25444_));
 sky130_fd_sc_hd__a211o_1 _28589_ (.A1(_23849_),
    .A2(_23846_),
    .B1(_25444_),
    .C1(_25441_),
    .X(_25445_));
 sky130_fd_sc_hd__a22oi_4 _28590_ (.A1(_25425_),
    .A2(_25429_),
    .B1(_25443_),
    .B2(_25445_),
    .Y(_00041_));
 sky130_fd_sc_hd__buf_2 _28591_ (.A(_25429_),
    .X(_00042_));
 sky130_fd_sc_hd__a41o_1 _28592_ (.A1(_25425_),
    .A2(_00042_),
    .A3(_25443_),
    .A4(_25445_),
    .B1(\delay_line[0][11] ),
    .X(_00043_));
 sky130_fd_sc_hd__a21o_1 _28593_ (.A1(_23849_),
    .A2(_23846_),
    .B1(_25441_),
    .X(_00044_));
 sky130_fd_sc_hd__o2111a_2 _28594_ (.A1(_25444_),
    .A2(_00044_),
    .B1(_25443_),
    .C1(_25425_),
    .D1(_25429_),
    .X(_00045_));
 sky130_fd_sc_hd__buf_1 _28595_ (.A(\delay_line[0][11] ),
    .X(_00046_));
 sky130_fd_sc_hd__o21ai_1 _28596_ (.A1(_00045_),
    .A2(_00041_),
    .B1(_00046_),
    .Y(_00047_));
 sky130_fd_sc_hd__o211ai_2 _28597_ (.A1(_00041_),
    .A2(_00043_),
    .B1(_23862_),
    .C1(_00047_),
    .Y(_00048_));
 sky130_fd_sc_hd__nor2b_1 _28598_ (.A(_18934_),
    .B_N(_23839_),
    .Y(_00049_));
 sky130_fd_sc_hd__or4_1 _28599_ (.A(_22304_),
    .B(_25430_),
    .C(_00049_),
    .D(_23838_),
    .X(_00050_));
 sky130_fd_sc_hd__and2_1 _28600_ (.A(_25438_),
    .B(_25440_),
    .X(_00052_));
 sky130_fd_sc_hd__a21oi_1 _28601_ (.A1(_23858_),
    .A2(_00050_),
    .B1(_00052_),
    .Y(_00053_));
 sky130_fd_sc_hd__o311a_1 _28602_ (.A1(_22311_),
    .A2(_25430_),
    .A3(_00049_),
    .B1(_00052_),
    .C1(_23858_),
    .X(_00054_));
 sky130_fd_sc_hd__o2bb2ai_2 _28603_ (.A1_N(_25425_),
    .A2_N(_00042_),
    .B1(_00053_),
    .B2(_00054_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand2_1 _28604_ (.A(_00055_),
    .B(_00046_),
    .Y(_00056_));
 sky130_fd_sc_hd__o21bai_2 _28605_ (.A1(_00045_),
    .A2(_00041_),
    .B1_N(\delay_line[0][11] ),
    .Y(_00057_));
 sky130_fd_sc_hd__o211ai_4 _28606_ (.A1(_00056_),
    .A2(_00045_),
    .B1(_23865_),
    .C1(_00057_),
    .Y(_00058_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28607_ (.A(\delay_line[0][10] ),
    .X(_00059_));
 sky130_fd_sc_hd__clkbuf_2 _28608_ (.A(_00059_),
    .X(_00060_));
 sky130_fd_sc_hd__a21oi_2 _28609_ (.A1(_00048_),
    .A2(_00058_),
    .B1(_00060_),
    .Y(_00061_));
 sky130_fd_sc_hd__o2111ai_1 _28610_ (.A1(_25444_),
    .A2(_00044_),
    .B1(_25443_),
    .C1(_25425_),
    .D1(_00042_),
    .Y(_00063_));
 sky130_fd_sc_hd__a21boi_1 _28611_ (.A1(_00063_),
    .A2(_00055_),
    .B1_N(_00046_),
    .Y(_00064_));
 sky130_fd_sc_hd__nor2_1 _28612_ (.A(_00041_),
    .B(_00043_),
    .Y(_00065_));
 sky130_fd_sc_hd__o311a_1 _28613_ (.A1(_23865_),
    .A2(_00064_),
    .A3(_00065_),
    .B1(_00060_),
    .C1(_00058_),
    .X(_00066_));
 sky130_fd_sc_hd__a21boi_2 _28614_ (.A1(_23868_),
    .A2(_23871_),
    .B1_N(_23864_),
    .Y(_00067_));
 sky130_fd_sc_hd__inv_2 _28615_ (.A(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__o21bai_4 _28616_ (.A1(_00061_),
    .A2(_00066_),
    .B1_N(_00068_),
    .Y(_00069_));
 sky130_fd_sc_hd__a21o_1 _28617_ (.A1(_00048_),
    .A2(_00058_),
    .B1(_00060_),
    .X(_00070_));
 sky130_fd_sc_hd__o31a_1 _28618_ (.A1(_23865_),
    .A2(_00064_),
    .A3(_00065_),
    .B1(_00059_),
    .X(_00071_));
 sky130_fd_sc_hd__nand2_1 _28619_ (.A(_00071_),
    .B(_00058_),
    .Y(_00072_));
 sky130_fd_sc_hd__nand3_4 _28620_ (.A(_00068_),
    .B(_00070_),
    .C(_00072_),
    .Y(_00074_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28621_ (.A(_22323_),
    .X(_00075_));
 sky130_fd_sc_hd__clkbuf_2 _28622_ (.A(_00075_),
    .X(_00076_));
 sky130_fd_sc_hd__clkbuf_2 _28623_ (.A(_00059_),
    .X(_00077_));
 sky130_fd_sc_hd__xor2_1 _28624_ (.A(_19986_),
    .B(\delay_line[13][11] ),
    .X(_00078_));
 sky130_fd_sc_hd__a21boi_2 _28625_ (.A1(_00076_),
    .A2(_00077_),
    .B1_N(_00078_),
    .Y(_00079_));
 sky130_fd_sc_hd__and3b_1 _28626_ (.A_N(_00078_),
    .B(_00060_),
    .C(_00076_),
    .X(_00080_));
 sky130_fd_sc_hd__o2bb2ai_1 _28627_ (.A1_N(_00069_),
    .A2_N(_00074_),
    .B1(_00079_),
    .B2(_00080_),
    .Y(_00081_));
 sky130_fd_sc_hd__and3_1 _28628_ (.A(_00075_),
    .B(_00059_),
    .C(_00078_),
    .X(_00082_));
 sky130_fd_sc_hd__a21oi_1 _28629_ (.A1(_00076_),
    .A2(_00077_),
    .B1(_00078_),
    .Y(_00083_));
 sky130_fd_sc_hd__o211ai_1 _28630_ (.A1(_00082_),
    .A2(_00083_),
    .B1(_00069_),
    .C1(_00074_),
    .Y(_00085_));
 sky130_fd_sc_hd__a32o_2 _28631_ (.A1(_23875_),
    .A2(_23876_),
    .A3(_23877_),
    .B1(_23873_),
    .B2(_23882_),
    .X(_00086_));
 sky130_fd_sc_hd__inv_2 _28632_ (.A(_00086_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand3_1 _28633_ (.A(_00081_),
    .B(_00085_),
    .C(_00087_),
    .Y(_00088_));
 sky130_fd_sc_hd__o2bb2ai_2 _28634_ (.A1_N(_00069_),
    .A2_N(_00074_),
    .B1(_00082_),
    .B2(_00083_),
    .Y(_00089_));
 sky130_fd_sc_hd__o211ai_4 _28635_ (.A1(_00079_),
    .A2(_00080_),
    .B1(_00069_),
    .C1(_00074_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand3_2 _28636_ (.A(_00086_),
    .B(_00089_),
    .C(_00090_),
    .Y(_00091_));
 sky130_fd_sc_hd__buf_2 _28637_ (.A(_23884_),
    .X(_00092_));
 sky130_fd_sc_hd__buf_1 _28638_ (.A(\delay_line[13][10] ),
    .X(_00093_));
 sky130_fd_sc_hd__a21o_1 _28639_ (.A1(_22362_),
    .A2(_00093_),
    .B1(_23879_),
    .X(_00094_));
 sky130_fd_sc_hd__buf_2 _28640_ (.A(_00093_),
    .X(_00096_));
 sky130_fd_sc_hd__nand3_1 _28641_ (.A(_22363_),
    .B(_23879_),
    .C(_00096_),
    .Y(_00097_));
 sky130_fd_sc_hd__and3_1 _28642_ (.A(_00094_),
    .B(_18962_),
    .C(_00097_),
    .X(_00098_));
 sky130_fd_sc_hd__clkbuf_2 _28643_ (.A(_18962_),
    .X(_00099_));
 sky130_fd_sc_hd__a21oi_2 _28644_ (.A1(_00097_),
    .A2(_00094_),
    .B1(_00099_),
    .Y(_00100_));
 sky130_fd_sc_hd__a311oi_2 _28645_ (.A1(_19982_),
    .A2(_19983_),
    .A3(_00092_),
    .B1(_00098_),
    .C1(_00100_),
    .Y(_00101_));
 sky130_fd_sc_hd__o211a_1 _28646_ (.A1(_00098_),
    .A2(_00100_),
    .B1(_00092_),
    .C1(_23880_),
    .X(_00102_));
 sky130_fd_sc_hd__o2bb2ai_1 _28647_ (.A1_N(_00088_),
    .A2_N(_00091_),
    .B1(_00101_),
    .B2(_00102_),
    .Y(_00103_));
 sky130_fd_sc_hd__o211a_1 _28648_ (.A1(_23818_),
    .A2(_22370_),
    .B1(_23883_),
    .C1(_23888_),
    .X(_00104_));
 sky130_fd_sc_hd__o21a_1 _28649_ (.A1(_23816_),
    .A2(_23817_),
    .B1(_23894_),
    .X(_00105_));
 sky130_fd_sc_hd__nor2_1 _28650_ (.A(_00104_),
    .B(_00105_),
    .Y(_00107_));
 sky130_fd_sc_hd__buf_2 _28651_ (.A(_00092_),
    .X(_00108_));
 sky130_fd_sc_hd__nor2_1 _28652_ (.A(_00098_),
    .B(_00100_),
    .Y(_00109_));
 sky130_fd_sc_hd__and3_1 _28653_ (.A(_00108_),
    .B(_23880_),
    .C(_00109_),
    .X(_00110_));
 sky130_fd_sc_hd__o2bb2a_1 _28654_ (.A1_N(_00108_),
    .A2_N(_23880_),
    .B1(_00098_),
    .B2(_00100_),
    .X(_00111_));
 sky130_fd_sc_hd__o211ai_1 _28655_ (.A1(_00110_),
    .A2(_00111_),
    .B1(_00088_),
    .C1(_00091_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand3_1 _28656_ (.A(_00103_),
    .B(_00107_),
    .C(_00112_),
    .Y(_00113_));
 sky130_fd_sc_hd__clkbuf_2 _28657_ (.A(_00113_),
    .X(_00114_));
 sky130_fd_sc_hd__buf_6 _28658_ (.A(_00088_),
    .X(_00115_));
 sky130_fd_sc_hd__o211ai_2 _28659_ (.A1(_00101_),
    .A2(_00102_),
    .B1(_00115_),
    .C1(_00091_),
    .Y(_00116_));
 sky130_fd_sc_hd__o2bb2ai_1 _28660_ (.A1_N(_00115_),
    .A2_N(_00091_),
    .B1(_00110_),
    .B2(_00111_),
    .Y(_00118_));
 sky130_fd_sc_hd__o211ai_4 _28661_ (.A1(_00104_),
    .A2(_00105_),
    .B1(_00116_),
    .C1(_00118_),
    .Y(_00119_));
 sky130_fd_sc_hd__buf_1 _28662_ (.A(\delay_line[12][11] ),
    .X(_00120_));
 sky130_fd_sc_hd__buf_2 _28663_ (.A(_00120_),
    .X(_00121_));
 sky130_fd_sc_hd__nand3b_2 _28664_ (.A_N(_23798_),
    .B(\delay_line[12][10] ),
    .C(\delay_line[12][11] ),
    .Y(_00122_));
 sky130_fd_sc_hd__inv_2 _28665_ (.A(\delay_line[12][10] ),
    .Y(_00123_));
 sky130_fd_sc_hd__or3b_2 _28666_ (.A(_00120_),
    .B(_00123_),
    .C_N(_23798_),
    .X(_00124_));
 sky130_fd_sc_hd__o2111ai_4 _28667_ (.A1(_23795_),
    .A2(_00121_),
    .B1(_00122_),
    .C1(_18985_),
    .D1(_00124_),
    .Y(_00125_));
 sky130_fd_sc_hd__o21a_1 _28668_ (.A1(_23800_),
    .A2(_00120_),
    .B1(_00122_),
    .X(_00126_));
 sky130_fd_sc_hd__a21o_1 _28669_ (.A1(_00124_),
    .A2(_00126_),
    .B1(_18985_),
    .X(_00127_));
 sky130_fd_sc_hd__nand2_1 _28670_ (.A(_17978_),
    .B(_23794_),
    .Y(_00129_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28671_ (.A(_18915_),
    .X(_00130_));
 sky130_fd_sc_hd__a21o_1 _28672_ (.A1(_12746_),
    .A2(_00130_),
    .B1(_17978_),
    .X(_00131_));
 sky130_fd_sc_hd__nand4_2 _28673_ (.A(_00125_),
    .B(_00127_),
    .C(_00129_),
    .D(_00131_),
    .Y(_00132_));
 sky130_fd_sc_hd__a22o_1 _28674_ (.A1(_00125_),
    .A2(_00127_),
    .B1(_00129_),
    .B2(_00131_),
    .X(_00133_));
 sky130_fd_sc_hd__a211oi_1 _28675_ (.A1(_00132_),
    .A2(_00133_),
    .B1(_23814_),
    .C1(_23897_),
    .Y(_00134_));
 sky130_fd_sc_hd__o211ai_2 _28676_ (.A1(_23814_),
    .A2(_23897_),
    .B1(_00132_),
    .C1(_00133_),
    .Y(_00135_));
 sky130_fd_sc_hd__inv_2 _28677_ (.A(_00135_),
    .Y(_00136_));
 sky130_fd_sc_hd__or3_1 _28678_ (.A(_00134_),
    .B(_23803_),
    .C(_00136_),
    .X(_00137_));
 sky130_fd_sc_hd__inv_2 _28679_ (.A(_00137_),
    .Y(_00138_));
 sky130_fd_sc_hd__o21a_1 _28680_ (.A1(_00136_),
    .A2(_00134_),
    .B1(_23803_),
    .X(_00140_));
 sky130_fd_sc_hd__nor2_1 _28681_ (.A(_00138_),
    .B(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__clkbuf_2 _28682_ (.A(_00141_),
    .X(_00142_));
 sky130_fd_sc_hd__a21oi_2 _28683_ (.A1(_00114_),
    .A2(_00119_),
    .B1(_00142_),
    .Y(_00143_));
 sky130_fd_sc_hd__o211a_1 _28684_ (.A1(_22411_),
    .A2(_23810_),
    .B1(_23895_),
    .C1(_23900_),
    .X(_00144_));
 sky130_fd_sc_hd__o21a_1 _28685_ (.A1(_23909_),
    .A2(_23910_),
    .B1(_23908_),
    .X(_00145_));
 sky130_fd_sc_hd__nand3_1 _28686_ (.A(_00119_),
    .B(_00142_),
    .C(_00114_),
    .Y(_00146_));
 sky130_fd_sc_hd__o21ai_1 _28687_ (.A1(_00144_),
    .A2(_00145_),
    .B1(_00146_),
    .Y(_00147_));
 sky130_fd_sc_hd__nor2_1 _28688_ (.A(_00143_),
    .B(_00147_),
    .Y(_00148_));
 sky130_fd_sc_hd__or2_1 _28689_ (.A(_00101_),
    .B(_00102_),
    .X(_00149_));
 sky130_fd_sc_hd__a21oi_1 _28690_ (.A1(_00115_),
    .A2(_00091_),
    .B1(_00149_),
    .Y(_00151_));
 sky130_fd_sc_hd__o21ai_1 _28691_ (.A1(_00104_),
    .A2(_00105_),
    .B1(_00116_),
    .Y(_00152_));
 sky130_fd_sc_hd__o21ai_1 _28692_ (.A1(_00151_),
    .A2(_00152_),
    .B1(_00114_),
    .Y(_00153_));
 sky130_fd_sc_hd__o21ai_2 _28693_ (.A1(_00138_),
    .A2(_00140_),
    .B1(_00153_),
    .Y(_00154_));
 sky130_fd_sc_hd__a21o_1 _28694_ (.A1(_23908_),
    .A2(_23915_),
    .B1(_00144_),
    .X(_00155_));
 sky130_fd_sc_hd__a21oi_1 _28695_ (.A1(_00146_),
    .A2(_00154_),
    .B1(_00155_),
    .Y(_00156_));
 sky130_fd_sc_hd__o22ai_1 _28696_ (.A1(_25407_),
    .A2(_25408_),
    .B1(_00148_),
    .B2(_00156_),
    .Y(_00157_));
 sky130_fd_sc_hd__inv_2 _28697_ (.A(_23917_),
    .Y(_00158_));
 sky130_fd_sc_hd__a21oi_1 _28698_ (.A1(_23790_),
    .A2(_23912_),
    .B1(_00158_),
    .Y(_00159_));
 sky130_fd_sc_hd__o21ba_1 _28699_ (.A1(_25366_),
    .A2(_25367_),
    .B1_N(_25406_),
    .X(_00160_));
 sky130_fd_sc_hd__clkbuf_2 _28700_ (.A(_00160_),
    .X(_00162_));
 sky130_fd_sc_hd__o211a_1 _28701_ (.A1(_23768_),
    .A2(_23781_),
    .B1(_25406_),
    .C1(_23780_),
    .X(_00163_));
 sky130_fd_sc_hd__o211a_1 _28702_ (.A1(_00151_),
    .A2(_00152_),
    .B1(_00141_),
    .C1(_00113_),
    .X(_00164_));
 sky130_fd_sc_hd__a21oi_1 _28703_ (.A1(_23908_),
    .A2(_23915_),
    .B1(_00144_),
    .Y(_00165_));
 sky130_fd_sc_hd__o21ai_2 _28704_ (.A1(_00164_),
    .A2(_00143_),
    .B1(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__o221ai_2 _28705_ (.A1(_00162_),
    .A2(_00163_),
    .B1(_00143_),
    .B2(_00147_),
    .C1(_00166_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand3_2 _28706_ (.A(_00157_),
    .B(_00159_),
    .C(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__clkbuf_2 _28707_ (.A(_00168_),
    .X(_00169_));
 sky130_fd_sc_hd__a31oi_2 _28708_ (.A1(_00114_),
    .A2(_00119_),
    .A3(_00142_),
    .B1(_00165_),
    .Y(_00170_));
 sky130_fd_sc_hd__a2bb2oi_1 _28709_ (.A1_N(_25407_),
    .A2_N(_25408_),
    .B1(_00154_),
    .B2(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__buf_6 _28710_ (.A(_00166_),
    .X(_00173_));
 sky130_fd_sc_hd__a21oi_1 _28711_ (.A1(_00171_),
    .A2(_00173_),
    .B1(_00159_),
    .Y(_00174_));
 sky130_fd_sc_hd__o22ai_1 _28712_ (.A1(_00162_),
    .A2(_00163_),
    .B1(_00148_),
    .B2(_00156_),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _28713_ (.A(_00174_),
    .B(_00175_),
    .Y(_00176_));
 sky130_fd_sc_hd__a2bb2oi_4 _28714_ (.A1_N(_25363_),
    .A2_N(_25365_),
    .B1(_00169_),
    .B2(_00176_),
    .Y(_00177_));
 sky130_fd_sc_hd__inv_2 _28715_ (.A(_24126_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _28716_ (.A(_00170_),
    .B(_00154_),
    .Y(_00179_));
 sky130_fd_sc_hd__a2bb2oi_2 _28717_ (.A1_N(_00162_),
    .A2_N(_00163_),
    .B1(_00179_),
    .B2(_00173_),
    .Y(_00180_));
 sky130_fd_sc_hd__a311oi_2 _28718_ (.A1(_23911_),
    .A2(_23791_),
    .A3(_23906_),
    .B1(_23788_),
    .C1(_23787_),
    .Y(_00181_));
 sky130_fd_sc_hd__o2bb2ai_2 _28719_ (.A1_N(_00173_),
    .A2_N(_00171_),
    .B1(_00158_),
    .B2(_00181_),
    .Y(_00182_));
 sky130_fd_sc_hd__xor2_2 _28720_ (.A(_25364_),
    .B(_25362_),
    .X(_00184_));
 sky130_fd_sc_hd__o211ai_4 _28721_ (.A1(_00180_),
    .A2(_00182_),
    .B1(_00184_),
    .C1(_00168_),
    .Y(_00185_));
 sky130_fd_sc_hd__o21ai_4 _28722_ (.A1(_24125_),
    .A2(_00178_),
    .B1(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__nor2_2 _28723_ (.A(_00177_),
    .B(_00186_),
    .Y(_00187_));
 sky130_fd_sc_hd__o21ai_1 _28724_ (.A1(_00180_),
    .A2(_00182_),
    .B1(_00169_),
    .Y(_00188_));
 sky130_fd_sc_hd__o21ai_4 _28725_ (.A1(_25363_),
    .A2(_25365_),
    .B1(_00188_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _28726_ (.A(_24007_),
    .B(_24126_),
    .Y(_00190_));
 sky130_fd_sc_hd__a21oi_4 _28727_ (.A1(_00189_),
    .A2(_00185_),
    .B1(_00190_),
    .Y(_00191_));
 sky130_fd_sc_hd__a311o_2 _28728_ (.A1(_21928_),
    .A2(_21929_),
    .A3(_22618_),
    .B1(_22617_),
    .C1(_24109_),
    .X(_00192_));
 sky130_fd_sc_hd__o21ai_4 _28729_ (.A1(_24078_),
    .A2(_24110_),
    .B1(_00192_),
    .Y(_00193_));
 sky130_fd_sc_hd__o21ai_2 _28730_ (.A1(_22481_),
    .A2(_22491_),
    .B1(_23994_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_2 _28731_ (.A(_13460_),
    .B(\delay_line[5][11] ),
    .Y(_00196_));
 sky130_fd_sc_hd__or2_1 _28732_ (.A(\delay_line[5][11] ),
    .B(_13460_),
    .X(_00197_));
 sky130_fd_sc_hd__nand3_1 _28733_ (.A(_00196_),
    .B(_00197_),
    .C(net430),
    .Y(_00198_));
 sky130_fd_sc_hd__a21o_1 _28734_ (.A1(_00196_),
    .A2(_00197_),
    .B1(net430),
    .X(_00199_));
 sky130_fd_sc_hd__a22o_2 _28735_ (.A1(_24058_),
    .A2(_21979_),
    .B1(_00198_),
    .B2(_00199_),
    .X(_00200_));
 sky130_fd_sc_hd__clkbuf_2 _28736_ (.A(_00198_),
    .X(_00201_));
 sky130_fd_sc_hd__nand4_2 _28737_ (.A(_00199_),
    .B(_24059_),
    .C(_24058_),
    .D(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand4_1 _28738_ (.A(_24045_),
    .B(_24048_),
    .C(_00200_),
    .D(_00202_),
    .Y(_00203_));
 sky130_fd_sc_hd__a22o_1 _28739_ (.A1(_24045_),
    .A2(_24048_),
    .B1(_00200_),
    .B2(_00202_),
    .X(_00204_));
 sky130_fd_sc_hd__nand2_1 _28740_ (.A(_00203_),
    .B(_00204_),
    .Y(_00206_));
 sky130_fd_sc_hd__clkbuf_2 _28741_ (.A(\delay_line[3][11] ),
    .X(_00207_));
 sky130_fd_sc_hd__xnor2_1 _28742_ (.A(_18104_),
    .B(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__xnor2_1 _28743_ (.A(_24041_),
    .B(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__xnor2_1 _28744_ (.A(_00206_),
    .B(_00209_),
    .Y(_00210_));
 sky130_fd_sc_hd__clkbuf_2 _28745_ (.A(_22606_),
    .X(_00211_));
 sky130_fd_sc_hd__nand3b_2 _28746_ (.A_N(_22596_),
    .B(\delay_line[6][10] ),
    .C(_22604_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand3b_2 _28747_ (.A_N(\delay_line[6][10] ),
    .B(_22596_),
    .C(_22604_),
    .Y(_00213_));
 sky130_fd_sc_hd__o211a_1 _28748_ (.A1(_00211_),
    .A2(_24084_),
    .B1(_00212_),
    .C1(_00213_),
    .X(_00214_));
 sky130_fd_sc_hd__o211a_1 _28749_ (.A1(_22604_),
    .A2(_24084_),
    .B1(_21979_),
    .C1(_00213_),
    .X(_00215_));
 sky130_fd_sc_hd__a2bb2o_1 _28750_ (.A1_N(_24059_),
    .A2_N(_00214_),
    .B1(_00215_),
    .B2(_00212_),
    .X(_00217_));
 sky130_fd_sc_hd__a21o_1 _28751_ (.A1(_24088_),
    .A2(_24096_),
    .B1(_00217_),
    .X(_00218_));
 sky130_fd_sc_hd__nand3_1 _28752_ (.A(_24088_),
    .B(_24096_),
    .C(_00217_),
    .Y(_00219_));
 sky130_fd_sc_hd__and3_1 _28753_ (.A(_00218_),
    .B(_24066_),
    .C(_00219_),
    .X(_00220_));
 sky130_fd_sc_hd__a21oi_1 _28754_ (.A1(_00219_),
    .A2(_00218_),
    .B1(_24066_),
    .Y(_00221_));
 sky130_fd_sc_hd__a211oi_1 _28755_ (.A1(_24068_),
    .A2(_24070_),
    .B1(_00220_),
    .C1(_00221_),
    .Y(_00222_));
 sky130_fd_sc_hd__o211a_1 _28756_ (.A1(_00220_),
    .A2(_00221_),
    .B1(_24068_),
    .C1(_24070_),
    .X(_00223_));
 sky130_fd_sc_hd__or3_1 _28757_ (.A(_00210_),
    .B(_00222_),
    .C(_00223_),
    .X(_00224_));
 sky130_fd_sc_hd__o21ai_1 _28758_ (.A1(_00222_),
    .A2(_00223_),
    .B1(_00210_),
    .Y(_00225_));
 sky130_fd_sc_hd__a32o_1 _28759_ (.A1(_24057_),
    .A2(_24069_),
    .A3(_24070_),
    .B1(_24073_),
    .B2(_24056_),
    .X(_00226_));
 sky130_fd_sc_hd__a21oi_1 _28760_ (.A1(_00224_),
    .A2(_00225_),
    .B1(_00226_),
    .Y(_00228_));
 sky130_fd_sc_hd__and3_1 _28761_ (.A(_00226_),
    .B(_00224_),
    .C(_00225_),
    .X(_00229_));
 sky130_fd_sc_hd__a21oi_1 _28762_ (.A1(_24030_),
    .A2(_24014_),
    .B1(_24026_),
    .Y(_00230_));
 sky130_fd_sc_hd__or2_1 _28763_ (.A(\delay_line[2][11] ),
    .B(_22638_),
    .X(_00231_));
 sky130_fd_sc_hd__nand2_1 _28764_ (.A(_22640_),
    .B(\delay_line[2][11] ),
    .Y(_00232_));
 sky130_fd_sc_hd__a22o_1 _28765_ (.A1(_24016_),
    .A2(_22674_),
    .B1(_00231_),
    .B2(_00232_),
    .X(_00233_));
 sky130_fd_sc_hd__nand4_2 _28766_ (.A(_22674_),
    .B(_00231_),
    .C(_24016_),
    .D(_00232_),
    .Y(_00234_));
 sky130_fd_sc_hd__and3_1 _28767_ (.A(_00233_),
    .B(_24043_),
    .C(_00234_),
    .X(_00235_));
 sky130_fd_sc_hd__a21oi_1 _28768_ (.A1(_00234_),
    .A2(_00233_),
    .B1(_24043_),
    .Y(_00236_));
 sky130_fd_sc_hd__o211ai_1 _28769_ (.A1(_00235_),
    .A2(_00236_),
    .B1(_24019_),
    .C1(_24024_),
    .Y(_00237_));
 sky130_fd_sc_hd__a211o_1 _28770_ (.A1(_24019_),
    .A2(_24024_),
    .B1(_00235_),
    .C1(_00236_),
    .X(_00239_));
 sky130_fd_sc_hd__nand2_1 _28771_ (.A(_00237_),
    .B(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__o21ba_1 _28772_ (.A1(_24054_),
    .A2(_24052_),
    .B1_N(_24051_),
    .X(_00241_));
 sky130_fd_sc_hd__xnor2_1 _28773_ (.A(_00240_),
    .B(_00241_),
    .Y(_00242_));
 sky130_fd_sc_hd__or2_1 _28774_ (.A(_00230_),
    .B(_00242_),
    .X(_00243_));
 sky130_fd_sc_hd__nand2_1 _28775_ (.A(_00242_),
    .B(_00230_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _28776_ (.A(_00243_),
    .B(_00244_),
    .Y(_00245_));
 sky130_fd_sc_hd__o21ai_1 _28777_ (.A1(_00228_),
    .A2(_00229_),
    .B1(_00245_),
    .Y(_00246_));
 sky130_fd_sc_hd__or3_1 _28778_ (.A(_00228_),
    .B(_00245_),
    .C(_00229_),
    .X(_00247_));
 sky130_fd_sc_hd__nand2_2 _28779_ (.A(_00246_),
    .B(_00247_),
    .Y(_00248_));
 sky130_fd_sc_hd__o21a_1 _28780_ (.A1(_24082_),
    .A2(_24103_),
    .B1(_24107_),
    .X(_00250_));
 sky130_fd_sc_hd__a21o_1 _28781_ (.A1(_23941_),
    .A2(_23965_),
    .B1(_23963_),
    .X(_00251_));
 sky130_fd_sc_hd__buf_1 _28782_ (.A(_18025_),
    .X(_00252_));
 sky130_fd_sc_hd__clkbuf_2 _28783_ (.A(\delay_line[7][6] ),
    .X(_00253_));
 sky130_fd_sc_hd__nand2_1 _28784_ (.A(_22591_),
    .B(net427),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2b_1 _28785_ (.A_N(net427),
    .B(_08965_),
    .Y(_00255_));
 sky130_fd_sc_hd__a22o_1 _28786_ (.A1(_00252_),
    .A2(_00253_),
    .B1(_00254_),
    .B2(_00255_),
    .X(_00256_));
 sky130_fd_sc_hd__nand4_2 _28787_ (.A(_00254_),
    .B(_00255_),
    .C(_18026_),
    .D(_00253_),
    .Y(_00257_));
 sky130_fd_sc_hd__and3_1 _28788_ (.A(_00256_),
    .B(_24086_),
    .C(_00257_),
    .X(_00258_));
 sky130_fd_sc_hd__o2bb2a_1 _28789_ (.A1_N(_00257_),
    .A2_N(_00256_),
    .B1(_21906_),
    .B2(_21910_),
    .X(_00259_));
 sky130_fd_sc_hd__clkbuf_2 _28790_ (.A(\delay_line[7][7] ),
    .X(_00261_));
 sky130_fd_sc_hd__nor2_1 _28791_ (.A(_24092_),
    .B(_00261_),
    .Y(_00262_));
 sky130_fd_sc_hd__and2_1 _28792_ (.A(_24092_),
    .B(_00261_),
    .X(_00263_));
 sky130_fd_sc_hd__o21bai_1 _28793_ (.A1(_00262_),
    .A2(_00263_),
    .B1_N(_00252_),
    .Y(_00264_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28794_ (.A(_00261_),
    .X(_00265_));
 sky130_fd_sc_hd__nand2_1 _28795_ (.A(_24092_),
    .B(_00265_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand3b_1 _28796_ (.A_N(_00262_),
    .B(_00266_),
    .C(_18026_),
    .Y(_00267_));
 sky130_fd_sc_hd__clkbuf_2 _28797_ (.A(_24091_),
    .X(_00268_));
 sky130_fd_sc_hd__and4_1 _28798_ (.A(_00264_),
    .B(_00267_),
    .C(_00268_),
    .D(_24093_),
    .X(_00269_));
 sky130_fd_sc_hd__a22oi_1 _28799_ (.A1(_00268_),
    .A2(_24093_),
    .B1(_00264_),
    .B2(_00267_),
    .Y(_00270_));
 sky130_fd_sc_hd__or4_2 _28800_ (.A(_00258_),
    .B(_00259_),
    .C(_00269_),
    .D(_00270_),
    .X(_00272_));
 sky130_fd_sc_hd__o22ai_1 _28801_ (.A1(_00258_),
    .A2(_00259_),
    .B1(_00269_),
    .B2(_00270_),
    .Y(_00273_));
 sky130_fd_sc_hd__o21bai_1 _28802_ (.A1(_22528_),
    .A2(_23935_),
    .B1_N(_23937_),
    .Y(_00274_));
 sky130_fd_sc_hd__and3_1 _28803_ (.A(_00272_),
    .B(_00273_),
    .C(_00274_),
    .X(_00275_));
 sky130_fd_sc_hd__a21oi_1 _28804_ (.A1(_00272_),
    .A2(_00273_),
    .B1(_00274_),
    .Y(_00276_));
 sky130_fd_sc_hd__o21bai_1 _28805_ (.A1(_00275_),
    .A2(_00276_),
    .B1_N(_24097_),
    .Y(_00277_));
 sky130_fd_sc_hd__or3b_1 _28806_ (.A(_00275_),
    .B(_00276_),
    .C_N(_24097_),
    .X(_00278_));
 sky130_fd_sc_hd__and3_1 _28807_ (.A(_00251_),
    .B(_00277_),
    .C(_00278_),
    .X(_00279_));
 sky130_fd_sc_hd__a21oi_1 _28808_ (.A1(_00277_),
    .A2(_00278_),
    .B1(_00251_),
    .Y(_00280_));
 sky130_fd_sc_hd__a21boi_1 _28809_ (.A1(_22608_),
    .A2(_24100_),
    .B1_N(_24099_),
    .Y(_00281_));
 sky130_fd_sc_hd__o21a_1 _28810_ (.A1(_00279_),
    .A2(_00280_),
    .B1(_00281_),
    .X(_00283_));
 sky130_fd_sc_hd__nor3_1 _28811_ (.A(_00281_),
    .B(_00279_),
    .C(_00280_),
    .Y(_00284_));
 sky130_fd_sc_hd__nor3_1 _28812_ (.A(_00250_),
    .B(_00283_),
    .C(_00284_),
    .Y(_00285_));
 sky130_fd_sc_hd__o21ai_1 _28813_ (.A1(_00283_),
    .A2(_00284_),
    .B1(_00250_),
    .Y(_00286_));
 sky130_fd_sc_hd__and2b_1 _28814_ (.A_N(_00285_),
    .B(_00286_),
    .X(_00287_));
 sky130_fd_sc_hd__xor2_4 _28815_ (.A(_00248_),
    .B(_00287_),
    .X(_00288_));
 sky130_fd_sc_hd__a21o_2 _28816_ (.A1(_00195_),
    .A2(_24003_),
    .B1(_00288_),
    .X(_00289_));
 sky130_fd_sc_hd__o211ai_2 _28817_ (.A1(_23927_),
    .A2(_23996_),
    .B1(_00195_),
    .C1(_00288_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_2 _28818_ (.A(_00289_),
    .B(_00290_),
    .Y(_00291_));
 sky130_fd_sc_hd__xor2_4 _28819_ (.A(_00193_),
    .B(_00291_),
    .X(_00292_));
 sky130_fd_sc_hd__inv_2 _28820_ (.A(_00292_),
    .Y(_00294_));
 sky130_fd_sc_hd__o21ai_2 _28821_ (.A1(_00187_),
    .A2(_00191_),
    .B1(_00294_),
    .Y(_00295_));
 sky130_fd_sc_hd__a21oi_2 _28822_ (.A1(_24119_),
    .A2(_24010_),
    .B1(_24129_),
    .Y(_00296_));
 sky130_fd_sc_hd__and3_2 _28823_ (.A(_00192_),
    .B(_24112_),
    .C(_00291_),
    .X(_00297_));
 sky130_fd_sc_hd__and3_2 _28824_ (.A(_00193_),
    .B(_00289_),
    .C(_00290_),
    .X(_00298_));
 sky130_fd_sc_hd__o211a_1 _28825_ (.A1(_00180_),
    .A2(_00182_),
    .B1(_00184_),
    .C1(_00169_),
    .X(_00299_));
 sky130_fd_sc_hd__o21bai_4 _28826_ (.A1(_00177_),
    .A2(_00299_),
    .B1_N(_00190_),
    .Y(_00300_));
 sky130_fd_sc_hd__o221ai_4 _28827_ (.A1(_00297_),
    .A2(_00298_),
    .B1(_00177_),
    .B2(_00186_),
    .C1(_00300_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand3_1 _28828_ (.A(_00295_),
    .B(_00296_),
    .C(_00301_),
    .Y(_00302_));
 sky130_fd_sc_hd__clkbuf_2 _28829_ (.A(_00302_),
    .X(_00303_));
 sky130_fd_sc_hd__o21bai_4 _28830_ (.A1(_00177_),
    .A2(_00186_),
    .B1_N(_00292_),
    .Y(_00305_));
 sky130_fd_sc_hd__buf_2 _28831_ (.A(_00191_),
    .X(_00306_));
 sky130_fd_sc_hd__a21o_2 _28832_ (.A1(_24119_),
    .A2(_24010_),
    .B1(_24129_),
    .X(_00307_));
 sky130_fd_sc_hd__o22ai_2 _28833_ (.A1(_00297_),
    .A2(_00298_),
    .B1(_00187_),
    .B2(_00306_),
    .Y(_00308_));
 sky130_fd_sc_hd__o211ai_4 _28834_ (.A1(_00305_),
    .A2(_00306_),
    .B1(_00307_),
    .C1(_00308_),
    .Y(_00309_));
 sky130_fd_sc_hd__nor2_2 _28835_ (.A(_24117_),
    .B(_24115_),
    .Y(_00310_));
 sky130_fd_sc_hd__inv_2 _28836_ (.A(_24168_),
    .Y(_00311_));
 sky130_fd_sc_hd__a21oi_1 _28837_ (.A1(_24166_),
    .A2(_22231_),
    .B1(_00311_),
    .Y(_00312_));
 sky130_fd_sc_hd__a21oi_1 _28838_ (.A1(_22657_),
    .A2(_22661_),
    .B1(_24031_),
    .Y(_00313_));
 sky130_fd_sc_hd__a21o_1 _28839_ (.A1(_20186_),
    .A2(_22234_),
    .B1(_22239_),
    .X(_00314_));
 sky130_fd_sc_hd__and2_1 _28840_ (.A(_00314_),
    .B(_22024_),
    .X(_00316_));
 sky130_fd_sc_hd__nor2b_1 _28841_ (.A(net448),
    .B_N(net449),
    .Y(_00317_));
 sky130_fd_sc_hd__nor2b_1 _28842_ (.A(net449),
    .B_N(net448),
    .Y(_00318_));
 sky130_fd_sc_hd__clkbuf_2 _28843_ (.A(_00318_),
    .X(_00319_));
 sky130_fd_sc_hd__nor3_1 _28844_ (.A(net442),
    .B(_00317_),
    .C(_00319_),
    .Y(_00320_));
 sky130_fd_sc_hd__o21a_1 _28845_ (.A1(_00317_),
    .A2(_00318_),
    .B1(net442),
    .X(_00321_));
 sky130_fd_sc_hd__nor3_1 _28846_ (.A(_00320_),
    .B(_24152_),
    .C(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__o2bb2a_1 _28847_ (.A1_N(net440),
    .A2_N(_24151_),
    .B1(_00321_),
    .B2(_00320_),
    .X(_00323_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28848_ (.A(\delay_line[1][10] ),
    .X(_00324_));
 sky130_fd_sc_hd__o2bb2a_1 _28849_ (.A1_N(_20193_),
    .A2_N(_00324_),
    .B1(_22234_),
    .B2(_22239_),
    .X(_00325_));
 sky130_fd_sc_hd__and4b_1 _28850_ (.A_N(_22234_),
    .B(_22236_),
    .C(_20193_),
    .D(_00324_),
    .X(_00327_));
 sky130_fd_sc_hd__o21ai_1 _28851_ (.A1(_22023_),
    .A2(_22235_),
    .B1(_22024_),
    .Y(_00328_));
 sky130_fd_sc_hd__o211a_1 _28852_ (.A1(_00325_),
    .A2(_00327_),
    .B1(_22236_),
    .C1(_00328_),
    .X(_00329_));
 sky130_fd_sc_hd__a211oi_1 _28853_ (.A1(_22236_),
    .A2(_00328_),
    .B1(_00325_),
    .C1(_00327_),
    .Y(_00330_));
 sky130_fd_sc_hd__or4_1 _28854_ (.A(_00322_),
    .B(_00323_),
    .C(_00329_),
    .D(_00330_),
    .X(_00331_));
 sky130_fd_sc_hd__o22ai_1 _28855_ (.A1(_00322_),
    .A2(_00323_),
    .B1(_00329_),
    .B2(_00330_),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _28856_ (.A(_24154_),
    .B(_24164_),
    .Y(_00333_));
 sky130_fd_sc_hd__a21oi_1 _28857_ (.A1(_00331_),
    .A2(_00332_),
    .B1(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__and3_1 _28858_ (.A(_00333_),
    .B(_00331_),
    .C(_00332_),
    .X(_00335_));
 sky130_fd_sc_hd__nor2_1 _28859_ (.A(_00334_),
    .B(_00335_),
    .Y(_00336_));
 sky130_fd_sc_hd__xnor2_1 _28860_ (.A(_00316_),
    .B(_00336_),
    .Y(_00338_));
 sky130_fd_sc_hd__nor3b_1 _28861_ (.A(_00313_),
    .B(_24034_),
    .C_N(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__o21ba_1 _28862_ (.A1(_00313_),
    .A2(_24034_),
    .B1_N(_00338_),
    .X(_00340_));
 sky130_fd_sc_hd__or3_1 _28863_ (.A(_00312_),
    .B(_00339_),
    .C(_00340_),
    .X(_00341_));
 sky130_fd_sc_hd__o21ai_1 _28864_ (.A1(_00339_),
    .A2(_00340_),
    .B1(_00312_),
    .Y(_00342_));
 sky130_fd_sc_hd__a221o_1 _28865_ (.A1(_24036_),
    .A2(_24076_),
    .B1(_00341_),
    .B2(_00342_),
    .C1(_24075_),
    .X(_00343_));
 sky130_fd_sc_hd__a21o_1 _28866_ (.A1(_24036_),
    .A2(_24076_),
    .B1(_24075_),
    .X(_00344_));
 sky130_fd_sc_hd__nand3_2 _28867_ (.A(_00344_),
    .B(_00341_),
    .C(_00342_),
    .Y(_00345_));
 sky130_fd_sc_hd__nand2_1 _28868_ (.A(_22247_),
    .B(_22249_),
    .Y(_00346_));
 sky130_fd_sc_hd__a21boi_1 _28869_ (.A1(_00346_),
    .A2(_24172_),
    .B1_N(_24173_),
    .Y(_00347_));
 sky130_fd_sc_hd__inv_2 _28870_ (.A(_00347_),
    .Y(_00349_));
 sky130_fd_sc_hd__a21o_1 _28871_ (.A1(_00343_),
    .A2(_00345_),
    .B1(_00349_),
    .X(_00350_));
 sky130_fd_sc_hd__nand3_2 _28872_ (.A(_00343_),
    .B(_00345_),
    .C(_00349_),
    .Y(_00351_));
 sky130_fd_sc_hd__a21bo_1 _28873_ (.A1(_24179_),
    .A2(_24145_),
    .B1_N(_24178_),
    .X(_00352_));
 sky130_fd_sc_hd__a21oi_1 _28874_ (.A1(_00350_),
    .A2(_00351_),
    .B1(_00352_),
    .Y(_00353_));
 sky130_fd_sc_hd__nand3_1 _28875_ (.A(_00352_),
    .B(_00350_),
    .C(_00351_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2b_1 _28876_ (.A_N(_00353_),
    .B(_00354_),
    .Y(_00355_));
 sky130_fd_sc_hd__xnor2_2 _28877_ (.A(_00310_),
    .B(_00355_),
    .Y(_00356_));
 sky130_fd_sc_hd__o21a_1 _28878_ (.A1(_24144_),
    .A2(_24180_),
    .B1(_00356_),
    .X(_00357_));
 sky130_fd_sc_hd__or2_1 _28879_ (.A(_24144_),
    .B(_24180_),
    .X(_00358_));
 sky130_fd_sc_hd__nor2_2 _28880_ (.A(_00358_),
    .B(_00356_),
    .Y(_00360_));
 sky130_fd_sc_hd__nor2_2 _28881_ (.A(_00357_),
    .B(_00360_),
    .Y(_00361_));
 sky130_fd_sc_hd__a21oi_4 _28882_ (.A1(_00303_),
    .A2(_00309_),
    .B1(_00361_),
    .Y(_00362_));
 sky130_fd_sc_hd__o211ai_4 _28883_ (.A1(_24125_),
    .A2(_00178_),
    .B1(_00189_),
    .C1(_00185_),
    .Y(_00363_));
 sky130_fd_sc_hd__a21oi_2 _28884_ (.A1(_00363_),
    .A2(_00300_),
    .B1(_00294_),
    .Y(_00364_));
 sky130_fd_sc_hd__o21ai_2 _28885_ (.A1(_00306_),
    .A2(_00305_),
    .B1(_00307_),
    .Y(_00365_));
 sky130_fd_sc_hd__o211ai_2 _28886_ (.A1(_00364_),
    .A2(_00365_),
    .B1(_00361_),
    .C1(_00303_),
    .Y(_00366_));
 sky130_fd_sc_hd__o21ai_1 _28887_ (.A1(_24188_),
    .A2(_24196_),
    .B1(_24135_),
    .Y(_00367_));
 sky130_fd_sc_hd__nand2_1 _28888_ (.A(_00366_),
    .B(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__nor2_1 _28889_ (.A(_00362_),
    .B(_00368_),
    .Y(_00369_));
 sky130_fd_sc_hd__o21ai_1 _28890_ (.A1(_00364_),
    .A2(_00365_),
    .B1(_00302_),
    .Y(_00371_));
 sky130_fd_sc_hd__o21ai_2 _28891_ (.A1(_00357_),
    .A2(_00360_),
    .B1(_00371_),
    .Y(_00372_));
 sky130_fd_sc_hd__a21oi_2 _28892_ (.A1(_00372_),
    .A2(_00366_),
    .B1(_00367_),
    .Y(_00373_));
 sky130_fd_sc_hd__o22a_1 _28893_ (.A1(_24183_),
    .A2(_24185_),
    .B1(_00369_),
    .B2(_00373_),
    .X(_00374_));
 sky130_fd_sc_hd__nand2_1 _28894_ (.A(_24141_),
    .B(_24195_),
    .Y(_00375_));
 sky130_fd_sc_hd__a31oi_1 _28895_ (.A1(_00303_),
    .A2(_00309_),
    .A3(_00361_),
    .B1(_00375_),
    .Y(_00376_));
 sky130_fd_sc_hd__a31o_1 _28896_ (.A1(_22701_),
    .A2(_24143_),
    .A3(_24181_),
    .B1(_24185_),
    .X(_00377_));
 sky130_fd_sc_hd__a21oi_2 _28897_ (.A1(_00376_),
    .A2(_00372_),
    .B1(_00377_),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_2 _28898_ (.A(_24195_),
    .Y(_00379_));
 sky130_fd_sc_hd__o211a_1 _28899_ (.A1(_00364_),
    .A2(_00365_),
    .B1(_00361_),
    .C1(_00303_),
    .X(_00380_));
 sky130_fd_sc_hd__o22ai_4 _28900_ (.A1(_24196_),
    .A2(_00379_),
    .B1(_00362_),
    .B2(_00380_),
    .Y(_00382_));
 sky130_fd_sc_hd__a22o_1 _28901_ (.A1(_24194_),
    .A2(_24210_),
    .B1(_00378_),
    .B2(_00382_),
    .X(_00383_));
 sky130_fd_sc_hd__o21ai_1 _28902_ (.A1(_00369_),
    .A2(_00373_),
    .B1(_24186_),
    .Y(_00384_));
 sky130_fd_sc_hd__o31a_1 _28903_ (.A1(_22266_),
    .A2(_24202_),
    .A3(_24211_),
    .B1(_24194_),
    .X(_00385_));
 sky130_fd_sc_hd__o211ai_2 _28904_ (.A1(_00362_),
    .A2(_00368_),
    .B1(_00377_),
    .C1(_00382_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand3_2 _28905_ (.A(_00384_),
    .B(_00385_),
    .C(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__o21a_1 _28906_ (.A1(_00374_),
    .A2(_00383_),
    .B1(_00387_),
    .X(_00388_));
 sky130_fd_sc_hd__o22ai_2 _28907_ (.A1(_24207_),
    .A2(_24217_),
    .B1(_24231_),
    .B2(_24232_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_2 _28908_ (.A(_00388_),
    .B(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__o21ai_2 _28909_ (.A1(_00374_),
    .A2(_00383_),
    .B1(_00387_),
    .Y(_00391_));
 sky130_fd_sc_hd__o211ai_4 _28910_ (.A1(_24232_),
    .A2(_24231_),
    .B1(_24213_),
    .C1(_00391_),
    .Y(_00393_));
 sky130_fd_sc_hd__nor2_1 _28911_ (.A(net348),
    .B(\delay_line[23][11] ),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_2 _28912_ (.A(\delay_line[23][11] ),
    .Y(_00395_));
 sky130_fd_sc_hd__nor2_1 _28913_ (.A(_24238_),
    .B(_00395_),
    .Y(_00396_));
 sky130_fd_sc_hd__nor2_1 _28914_ (.A(_00394_),
    .B(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand3_2 _28915_ (.A(_00390_),
    .B(_00393_),
    .C(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__clkbuf_2 _28916_ (.A(_00396_),
    .X(_00399_));
 sky130_fd_sc_hd__nand2_1 _28917_ (.A(_00391_),
    .B(_00389_),
    .Y(_00400_));
 sky130_fd_sc_hd__o21a_1 _28918_ (.A1(_22720_),
    .A2(_23747_),
    .B1(_24200_),
    .X(_00401_));
 sky130_fd_sc_hd__a31o_2 _28919_ (.A1(_24190_),
    .A2(_24191_),
    .A3(_24189_),
    .B1(_00401_),
    .X(_00402_));
 sky130_fd_sc_hd__nand2_2 _28920_ (.A(_00386_),
    .B(_00384_),
    .Y(_00404_));
 sky130_fd_sc_hd__a21oi_1 _28921_ (.A1(_24194_),
    .A2(_00401_),
    .B1(_24205_),
    .Y(_00405_));
 sky130_fd_sc_hd__a22oi_4 _28922_ (.A1(_24194_),
    .A2(_24210_),
    .B1(_00378_),
    .B2(_00382_),
    .Y(_00406_));
 sky130_fd_sc_hd__o22ai_4 _28923_ (.A1(_24183_),
    .A2(_24185_),
    .B1(_00369_),
    .B2(_00373_),
    .Y(_00407_));
 sky130_fd_sc_hd__a22oi_4 _28924_ (.A1(_24209_),
    .A2(_00405_),
    .B1(_00406_),
    .B2(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__o211ai_4 _28925_ (.A1(_00402_),
    .A2(_00404_),
    .B1(_00408_),
    .C1(_24224_),
    .Y(_00409_));
 sky130_fd_sc_hd__o211ai_2 _28926_ (.A1(_00394_),
    .A2(_00399_),
    .B1(_00400_),
    .C1(_00409_),
    .Y(_00410_));
 sky130_fd_sc_hd__o211ai_4 _28927_ (.A1(_25293_),
    .A2(_25061_),
    .B1(_00398_),
    .C1(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__o211ai_1 _28928_ (.A1(_00394_),
    .A2(_00399_),
    .B1(_00390_),
    .C1(_00393_),
    .Y(_00412_));
 sky130_fd_sc_hd__a21oi_1 _28929_ (.A1(_25059_),
    .A2(_25044_),
    .B1(_25293_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand3_1 _28930_ (.A(_00400_),
    .B(_00409_),
    .C(_00397_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand3_2 _28931_ (.A(_00412_),
    .B(_00413_),
    .C(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__a21oi_1 _28932_ (.A1(_24240_),
    .A2(_24252_),
    .B1(_24245_),
    .Y(_00417_));
 sky130_fd_sc_hd__a21boi_2 _28933_ (.A1(_00411_),
    .A2(_00416_),
    .B1_N(_00417_),
    .Y(_00418_));
 sky130_fd_sc_hd__o211a_2 _28934_ (.A1(_24245_),
    .A2(_24236_),
    .B1(_00411_),
    .C1(_00416_),
    .X(_00419_));
 sky130_fd_sc_hd__nor3_2 _28935_ (.A(_25291_),
    .B(_00418_),
    .C(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__a21bo_1 _28936_ (.A1(_00411_),
    .A2(_00416_),
    .B1_N(_00417_),
    .X(_00421_));
 sky130_fd_sc_hd__o211ai_2 _28937_ (.A1(_24245_),
    .A2(_24236_),
    .B1(_00411_),
    .C1(_00416_),
    .Y(_00422_));
 sky130_fd_sc_hd__a21oi_1 _28938_ (.A1(_00421_),
    .A2(_00422_),
    .B1(_25290_),
    .Y(_00423_));
 sky130_fd_sc_hd__o21ai_2 _28939_ (.A1(_24254_),
    .A2(_24249_),
    .B1(_24257_),
    .Y(_00424_));
 sky130_fd_sc_hd__o21ai_1 _28940_ (.A1(_00420_),
    .A2(_00423_),
    .B1(_00424_),
    .Y(_00426_));
 sky130_fd_sc_hd__nand3_1 _28941_ (.A(_25290_),
    .B(_00421_),
    .C(_00422_),
    .Y(_00427_));
 sky130_fd_sc_hd__o21ai_2 _28942_ (.A1(_00418_),
    .A2(_00419_),
    .B1(_25291_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand4_2 _28943_ (.A(_24257_),
    .B(_24258_),
    .C(_00427_),
    .D(_00428_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand4_4 _28944_ (.A(_24267_),
    .B(_25288_),
    .C(_00426_),
    .D(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__a22oi_1 _28945_ (.A1(_24257_),
    .A2(_24258_),
    .B1(_00427_),
    .B2(_00428_),
    .Y(_00431_));
 sky130_fd_sc_hd__nor3_1 _28946_ (.A(_00424_),
    .B(_00420_),
    .C(_00423_),
    .Y(_00432_));
 sky130_fd_sc_hd__o2bb2ai_2 _28947_ (.A1_N(_24267_),
    .A2_N(_25288_),
    .B1(_00431_),
    .B2(_00432_),
    .Y(_00433_));
 sky130_fd_sc_hd__mux2_1 _28948_ (.A0(_04623_),
    .A1(_15427_),
    .S(_24289_),
    .X(_00434_));
 sky130_fd_sc_hd__clkbuf_2 _28949_ (.A(_22129_),
    .X(_00435_));
 sky130_fd_sc_hd__buf_2 _28950_ (.A(_24250_),
    .X(_00437_));
 sky130_fd_sc_hd__nand2_2 _28951_ (.A(_22782_),
    .B(_24241_),
    .Y(_00438_));
 sky130_fd_sc_hd__or2_1 _28952_ (.A(_22782_),
    .B(_24241_),
    .X(_00439_));
 sky130_fd_sc_hd__a22o_1 _28953_ (.A1(_00435_),
    .A2(_00437_),
    .B1(_00438_),
    .B2(_00439_),
    .X(_00440_));
 sky130_fd_sc_hd__nand4_4 _28954_ (.A(_00439_),
    .B(_00437_),
    .C(_00435_),
    .D(_00438_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand3_1 _28955_ (.A(_00434_),
    .B(_00440_),
    .C(_00441_),
    .Y(_00442_));
 sky130_fd_sc_hd__inv_2 _28956_ (.A(_00442_),
    .Y(_00443_));
 sky130_fd_sc_hd__a21oi_1 _28957_ (.A1(_00441_),
    .A2(_00440_),
    .B1(_00434_),
    .Y(_00444_));
 sky130_fd_sc_hd__o2bb2ai_1 _28958_ (.A1_N(_00430_),
    .A2_N(_00433_),
    .B1(_00443_),
    .B2(_00444_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _28959_ (.A(_00441_),
    .B(_00440_),
    .Y(_00446_));
 sky130_fd_sc_hd__nor2_1 _28960_ (.A(_00446_),
    .B(_00434_),
    .Y(_00448_));
 sky130_fd_sc_hd__and2_1 _28961_ (.A(_00434_),
    .B(_00446_),
    .X(_00449_));
 sky130_fd_sc_hd__clkbuf_2 _28962_ (.A(_00433_),
    .X(_00450_));
 sky130_fd_sc_hd__o211ai_1 _28963_ (.A1(_00448_),
    .A2(_00449_),
    .B1(_00430_),
    .C1(_00450_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand3b_1 _28964_ (.A_N(_25287_),
    .B(_00445_),
    .C(_00451_),
    .Y(_00452_));
 sky130_fd_sc_hd__clkbuf_2 _28965_ (.A(_00452_),
    .X(_00453_));
 sky130_fd_sc_hd__o2bb2ai_1 _28966_ (.A1_N(_00430_),
    .A2_N(_00433_),
    .B1(_00448_),
    .B2(_00449_),
    .Y(_00454_));
 sky130_fd_sc_hd__o211ai_1 _28967_ (.A1(_00443_),
    .A2(_00444_),
    .B1(_00430_),
    .C1(_00450_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand3_2 _28968_ (.A(_00454_),
    .B(_00455_),
    .C(_25287_),
    .Y(_00456_));
 sky130_fd_sc_hd__or2_1 _28969_ (.A(_24288_),
    .B(_24291_),
    .X(_00457_));
 sky130_fd_sc_hd__o32a_1 _28970_ (.A1(_24268_),
    .A2(_24273_),
    .A3(_24298_),
    .B1(_00457_),
    .B2(_24279_),
    .X(_00459_));
 sky130_fd_sc_hd__a21bo_1 _28971_ (.A1(_00453_),
    .A2(_00456_),
    .B1_N(_00459_),
    .X(_00460_));
 sky130_fd_sc_hd__nor2_1 _28972_ (.A(_00457_),
    .B(_24279_),
    .Y(_00461_));
 sky130_fd_sc_hd__o211ai_1 _28973_ (.A1(_25207_),
    .A2(_00461_),
    .B1(_00453_),
    .C1(_00456_),
    .Y(_00462_));
 sky130_fd_sc_hd__o21a_1 _28974_ (.A1(_24493_),
    .A2(_24862_),
    .B1(_24861_),
    .X(_00463_));
 sky130_fd_sc_hd__o21ai_4 _28975_ (.A1(_24539_),
    .A2(_24498_),
    .B1(_24538_),
    .Y(_00464_));
 sky130_fd_sc_hd__clkbuf_2 _28976_ (.A(_06799_),
    .X(_00465_));
 sky130_fd_sc_hd__o2bb2a_1 _28977_ (.A1_N(_17150_),
    .A2_N(_06777_),
    .B1(_22836_),
    .B2(_17182_),
    .X(_00466_));
 sky130_fd_sc_hd__a32oi_2 _28978_ (.A1(_24510_),
    .A2(_24514_),
    .A3(_24515_),
    .B1(_24519_),
    .B2(_00466_),
    .Y(_00467_));
 sky130_fd_sc_hd__and2b_1 _28979_ (.A_N(_17171_),
    .B(_17248_),
    .X(_00468_));
 sky130_fd_sc_hd__nand3b_2 _28980_ (.A_N(_17248_),
    .B(_17171_),
    .C(_17139_),
    .Y(_00470_));
 sky130_fd_sc_hd__and3_1 _28981_ (.A(_17259_),
    .B(_00470_),
    .C(_17182_),
    .X(_00471_));
 sky130_fd_sc_hd__and2_1 _28982_ (.A(_22814_),
    .B(\delay_line[25][11] ),
    .X(_00472_));
 sky130_fd_sc_hd__buf_1 _28983_ (.A(_00472_),
    .X(_00473_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _28984_ (.A(\delay_line[25][11] ),
    .X(_00474_));
 sky130_fd_sc_hd__o211ai_2 _28985_ (.A1(_22819_),
    .A2(_00474_),
    .B1(_24505_),
    .C1(_21563_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _28986_ (.A(_22814_),
    .B(\delay_line[25][11] ),
    .Y(_00476_));
 sky130_fd_sc_hd__o21bai_2 _28987_ (.A1(_00472_),
    .A2(_00476_),
    .B1_N(_24503_),
    .Y(_00477_));
 sky130_fd_sc_hd__o211a_1 _28988_ (.A1(_00473_),
    .A2(_00475_),
    .B1(_21569_),
    .C1(_00477_),
    .X(_00478_));
 sky130_fd_sc_hd__a21o_1 _28989_ (.A1(_22819_),
    .A2(_00474_),
    .B1(_00475_),
    .X(_00479_));
 sky130_fd_sc_hd__a21o_1 _28990_ (.A1(_00479_),
    .A2(_00477_),
    .B1(_21569_),
    .X(_00481_));
 sky130_fd_sc_hd__o2bb2ai_1 _28991_ (.A1_N(_24507_),
    .A2_N(_24509_),
    .B1(_24506_),
    .B2(_24504_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand3b_2 _28992_ (.A_N(_00478_),
    .B(_00481_),
    .C(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__buf_1 _28993_ (.A(_21569_),
    .X(_00484_));
 sky130_fd_sc_hd__a21oi_1 _28994_ (.A1(_00479_),
    .A2(_00477_),
    .B1(_00484_),
    .Y(_00485_));
 sky130_fd_sc_hd__o21bai_2 _28995_ (.A1(_00478_),
    .A2(_00485_),
    .B1_N(_00482_),
    .Y(_00486_));
 sky130_fd_sc_hd__o211ai_1 _28996_ (.A1(_00468_),
    .A2(_00471_),
    .B1(_00483_),
    .C1(_00486_),
    .Y(_00487_));
 sky130_fd_sc_hd__a31o_1 _28997_ (.A1(_17259_),
    .A2(_00470_),
    .A3(_17182_),
    .B1(_00468_),
    .X(_00488_));
 sky130_fd_sc_hd__a21o_1 _28998_ (.A1(_00483_),
    .A2(_00486_),
    .B1(_00488_),
    .X(_00489_));
 sky130_fd_sc_hd__nand3b_2 _28999_ (.A_N(_00467_),
    .B(_00487_),
    .C(_00489_),
    .Y(_00490_));
 sky130_fd_sc_hd__o211a_1 _29000_ (.A1(_00468_),
    .A2(_00471_),
    .B1(_00483_),
    .C1(_00486_),
    .X(_00492_));
 sky130_fd_sc_hd__a21oi_1 _29001_ (.A1(_00483_),
    .A2(_00486_),
    .B1(_00488_),
    .Y(_00493_));
 sky130_fd_sc_hd__o21ai_2 _29002_ (.A1(_00492_),
    .A2(_00493_),
    .B1(_00467_),
    .Y(_00494_));
 sky130_fd_sc_hd__o2111ai_4 _29003_ (.A1(_06821_),
    .A2(_00465_),
    .B1(_24499_),
    .C1(_00490_),
    .D1(_00494_),
    .Y(_00495_));
 sky130_fd_sc_hd__o21a_1 _29004_ (.A1(_06799_),
    .A2(_06821_),
    .B1(_24499_),
    .X(_00496_));
 sky130_fd_sc_hd__a21o_1 _29005_ (.A1(_00494_),
    .A2(_00490_),
    .B1(_00496_),
    .X(_00497_));
 sky130_fd_sc_hd__nand2_1 _29006_ (.A(_24528_),
    .B(_24529_),
    .Y(_00498_));
 sky130_fd_sc_hd__a21o_1 _29007_ (.A1(_00495_),
    .A2(_00497_),
    .B1(_00498_),
    .X(_00499_));
 sky130_fd_sc_hd__nand3_2 _29008_ (.A(_00498_),
    .B(_00495_),
    .C(_00497_),
    .Y(_00500_));
 sky130_fd_sc_hd__a21o_1 _29009_ (.A1(_00499_),
    .A2(_00500_),
    .B1(_24530_),
    .X(_00501_));
 sky130_fd_sc_hd__nand3_2 _29010_ (.A(_00499_),
    .B(_00500_),
    .C(_24530_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _29011_ (.A(_24529_),
    .B(_24531_),
    .Y(_00504_));
 sky130_fd_sc_hd__o31a_1 _29012_ (.A1(_22811_),
    .A2(_22830_),
    .A3(_22832_),
    .B1(_22835_),
    .X(_00505_));
 sky130_fd_sc_hd__o2bb2a_1 _29013_ (.A1_N(_00501_),
    .A2_N(_00503_),
    .B1(_00504_),
    .B2(_00505_),
    .X(_00506_));
 sky130_fd_sc_hd__and4b_1 _29014_ (.A_N(_00504_),
    .B(_24532_),
    .C(_00501_),
    .D(_00503_),
    .X(_00507_));
 sky130_fd_sc_hd__or2_2 _29015_ (.A(_00506_),
    .B(_00507_),
    .X(_00508_));
 sky130_fd_sc_hd__xor2_4 _29016_ (.A(_00464_),
    .B(_00508_),
    .X(_00509_));
 sky130_fd_sc_hd__and3_1 _29017_ (.A(_24565_),
    .B(_24562_),
    .C(_24561_),
    .X(_00510_));
 sky130_fd_sc_hd__a21o_1 _29018_ (.A1(_24569_),
    .A2(_24542_),
    .B1(_00510_),
    .X(_00511_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29019_ (.A(_19501_),
    .X(_00512_));
 sky130_fd_sc_hd__clkbuf_2 _29020_ (.A(_24543_),
    .X(_00514_));
 sky130_fd_sc_hd__a21oi_1 _29021_ (.A1(_00512_),
    .A2(_00514_),
    .B1(_24544_),
    .Y(_00515_));
 sky130_fd_sc_hd__inv_2 _29022_ (.A(net353),
    .Y(_00516_));
 sky130_fd_sc_hd__clkbuf_2 _29023_ (.A(_00516_),
    .X(_00517_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29024_ (.A(\delay_line[22][10] ),
    .X(_00518_));
 sky130_fd_sc_hd__nor2_1 _29025_ (.A(_20449_),
    .B(_00518_),
    .Y(_00519_));
 sky130_fd_sc_hd__inv_2 _29026_ (.A(_24543_),
    .Y(_00520_));
 sky130_fd_sc_hd__and2_1 _29027_ (.A(_20449_),
    .B(\delay_line[22][10] ),
    .X(_00521_));
 sky130_fd_sc_hd__nor4_1 _29028_ (.A(_00517_),
    .B(_00519_),
    .C(_00520_),
    .D(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__o22a_1 _29029_ (.A1(_00516_),
    .A2(_00520_),
    .B1(_00521_),
    .B2(_00519_),
    .X(_00523_));
 sky130_fd_sc_hd__nand2_1 _29030_ (.A(_24549_),
    .B(_17073_),
    .Y(_00525_));
 sky130_fd_sc_hd__o21a_1 _29031_ (.A1(net356),
    .A2(_17073_),
    .B1(_21600_),
    .X(_00526_));
 sky130_fd_sc_hd__a2bb2oi_1 _29032_ (.A1_N(_17084_),
    .A2_N(_21600_),
    .B1(_00525_),
    .B2(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__o21ai_1 _29033_ (.A1(_00522_),
    .A2(_00523_),
    .B1(_00527_),
    .Y(_00528_));
 sky130_fd_sc_hd__or4bb_1 _29034_ (.A(_00521_),
    .B(_00519_),
    .C_N(_19501_),
    .D_N(_24555_),
    .X(_00529_));
 sky130_fd_sc_hd__a2bb2o_1 _29035_ (.A1_N(_00521_),
    .A2_N(_00519_),
    .B1(_00512_),
    .B2(_00514_),
    .X(_00530_));
 sky130_fd_sc_hd__nand3b_1 _29036_ (.A_N(_00527_),
    .B(_00529_),
    .C(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__o211ai_1 _29037_ (.A1(_00515_),
    .A2(_24553_),
    .B1(_00528_),
    .C1(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__a31o_1 _29038_ (.A1(_24550_),
    .A2(_24554_),
    .A3(_24552_),
    .B1(_00515_),
    .X(_00533_));
 sky130_fd_sc_hd__a21o_1 _29039_ (.A1(_00528_),
    .A2(_00531_),
    .B1(_00533_),
    .X(_00534_));
 sky130_fd_sc_hd__o2111ai_1 _29040_ (.A1(_06876_),
    .A2(_22852_),
    .B1(_01424_),
    .C1(_00532_),
    .D1(_00534_),
    .Y(_00536_));
 sky130_fd_sc_hd__a22o_1 _29041_ (.A1(_24554_),
    .A2(_01413_),
    .B1(_00534_),
    .B2(_00532_),
    .X(_00537_));
 sky130_fd_sc_hd__nand2_1 _29042_ (.A(_24559_),
    .B(_24561_),
    .Y(_00538_));
 sky130_fd_sc_hd__a21oi_1 _29043_ (.A1(_00536_),
    .A2(_00537_),
    .B1(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__and3_1 _29044_ (.A(_00538_),
    .B(_00536_),
    .C(_00537_),
    .X(_00540_));
 sky130_fd_sc_hd__or4_1 _29045_ (.A(_24541_),
    .B(_24566_),
    .C(_00539_),
    .D(_00540_),
    .X(_00541_));
 sky130_fd_sc_hd__o22ai_2 _29046_ (.A1(_24541_),
    .A2(_24566_),
    .B1(_00539_),
    .B2(_00540_),
    .Y(_00542_));
 sky130_fd_sc_hd__and3_1 _29047_ (.A(_00511_),
    .B(_00541_),
    .C(_00542_),
    .X(_00543_));
 sky130_fd_sc_hd__a21oi_1 _29048_ (.A1(_00541_),
    .A2(_00542_),
    .B1(_00511_),
    .Y(_00544_));
 sky130_fd_sc_hd__o21ai_1 _29049_ (.A1(_19519_),
    .A2(_20464_),
    .B1(_18309_),
    .Y(_00545_));
 sky130_fd_sc_hd__o21ai_1 _29050_ (.A1(_18309_),
    .A2(_24575_),
    .B1(_00545_),
    .Y(_00547_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29051_ (.A(\delay_line[24][7] ),
    .X(_00548_));
 sky130_fd_sc_hd__and2_2 _29052_ (.A(\delay_line[24][6] ),
    .B(_00548_),
    .X(_00549_));
 sky130_fd_sc_hd__o21ai_2 _29053_ (.A1(_20463_),
    .A2(_00548_),
    .B1(_19512_),
    .Y(_00550_));
 sky130_fd_sc_hd__clkbuf_2 _29054_ (.A(\delay_line[24][10] ),
    .X(_00551_));
 sky130_fd_sc_hd__nor2_1 _29055_ (.A(_20463_),
    .B(_21619_),
    .Y(_00552_));
 sky130_fd_sc_hd__o21ai_2 _29056_ (.A1(_00549_),
    .A2(_00552_),
    .B1(_22877_),
    .Y(_00553_));
 sky130_fd_sc_hd__o211a_1 _29057_ (.A1(_00549_),
    .A2(_00550_),
    .B1(_00551_),
    .C1(_00553_),
    .X(_00554_));
 sky130_fd_sc_hd__a21o_1 _29058_ (.A1(_20464_),
    .A2(_21619_),
    .B1(_00550_),
    .X(_00555_));
 sky130_fd_sc_hd__a21oi_1 _29059_ (.A1(_00555_),
    .A2(_00553_),
    .B1(_00551_),
    .Y(_00556_));
 sky130_fd_sc_hd__o21bai_1 _29060_ (.A1(_00554_),
    .A2(_00556_),
    .B1_N(_24581_),
    .Y(_00558_));
 sky130_fd_sc_hd__clkbuf_2 _29061_ (.A(\delay_line[24][10] ),
    .X(_00559_));
 sky130_fd_sc_hd__clkbuf_2 _29062_ (.A(_00559_),
    .X(_00560_));
 sky130_fd_sc_hd__o211ai_2 _29063_ (.A1(_00549_),
    .A2(_00550_),
    .B1(_00560_),
    .C1(_00553_),
    .Y(_00561_));
 sky130_fd_sc_hd__a21o_1 _29064_ (.A1(_00555_),
    .A2(_00553_),
    .B1(_00560_),
    .X(_00562_));
 sky130_fd_sc_hd__nand3_1 _29065_ (.A(_24586_),
    .B(_00561_),
    .C(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand3_1 _29066_ (.A(_00547_),
    .B(_00558_),
    .C(_00563_),
    .Y(_00564_));
 sky130_fd_sc_hd__o21ai_1 _29067_ (.A1(_00554_),
    .A2(_00556_),
    .B1(_24586_),
    .Y(_00565_));
 sky130_fd_sc_hd__o21a_1 _29068_ (.A1(_18309_),
    .A2(_24575_),
    .B1(_00545_),
    .X(_00566_));
 sky130_fd_sc_hd__nand3b_1 _29069_ (.A_N(_24581_),
    .B(_00561_),
    .C(_00562_),
    .Y(_00567_));
 sky130_fd_sc_hd__nand3_1 _29070_ (.A(_00565_),
    .B(_00566_),
    .C(_00567_),
    .Y(_00569_));
 sky130_fd_sc_hd__a21oi_1 _29071_ (.A1(_24586_),
    .A2(_24584_),
    .B1(_22890_),
    .Y(_00570_));
 sky130_fd_sc_hd__o21ai_1 _29072_ (.A1(_24573_),
    .A2(_00570_),
    .B1(_24590_),
    .Y(_00571_));
 sky130_fd_sc_hd__a21o_1 _29073_ (.A1(_00564_),
    .A2(_00569_),
    .B1(_00571_),
    .X(_00572_));
 sky130_fd_sc_hd__xor2_1 _29074_ (.A(_19508_),
    .B(_24572_),
    .X(_00573_));
 sky130_fd_sc_hd__nand3_1 _29075_ (.A(_00571_),
    .B(_00564_),
    .C(_00569_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand3_1 _29076_ (.A(_00572_),
    .B(_00573_),
    .C(_00574_),
    .Y(_00575_));
 sky130_fd_sc_hd__a21o_1 _29077_ (.A1(_00574_),
    .A2(_00572_),
    .B1(_00573_),
    .X(_00576_));
 sky130_fd_sc_hd__o21bai_1 _29078_ (.A1(_24597_),
    .A2(_24594_),
    .B1_N(_24593_),
    .Y(_00577_));
 sky130_fd_sc_hd__a21o_1 _29079_ (.A1(_00575_),
    .A2(_00576_),
    .B1(_00577_),
    .X(_00578_));
 sky130_fd_sc_hd__nand3_1 _29080_ (.A(_00577_),
    .B(_00575_),
    .C(_00576_),
    .Y(_00580_));
 sky130_fd_sc_hd__and3_1 _29081_ (.A(_00578_),
    .B(_00580_),
    .C(_24596_),
    .X(_00581_));
 sky130_fd_sc_hd__o2bb2a_1 _29082_ (.A1_N(_00578_),
    .A2_N(_00580_),
    .B1(_18305_),
    .B2(_21618_),
    .X(_00582_));
 sky130_fd_sc_hd__nor2_1 _29083_ (.A(_00581_),
    .B(_00582_),
    .Y(_00583_));
 sky130_fd_sc_hd__o22ai_2 _29084_ (.A1(_24603_),
    .A2(_24599_),
    .B1(_24604_),
    .B2(_24608_),
    .Y(_00584_));
 sky130_fd_sc_hd__or2_1 _29085_ (.A(_00583_),
    .B(_00584_),
    .X(_00585_));
 sky130_fd_sc_hd__nand2_2 _29086_ (.A(_00584_),
    .B(_00583_),
    .Y(_00586_));
 sky130_fd_sc_hd__or4bb_1 _29087_ (.A(_00543_),
    .B(_00544_),
    .C_N(_00585_),
    .D_N(_00586_),
    .X(_00587_));
 sky130_fd_sc_hd__inv_2 _29088_ (.A(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__a2bb2oi_1 _29089_ (.A1_N(_00543_),
    .A2_N(_00544_),
    .B1(_00585_),
    .B2(_00586_),
    .Y(_00589_));
 sky130_fd_sc_hd__nor2_1 _29090_ (.A(_00588_),
    .B(_00589_),
    .Y(_00591_));
 sky130_fd_sc_hd__xnor2_2 _29091_ (.A(_00509_),
    .B(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__nor3_1 _29092_ (.A(net108),
    .B(_24727_),
    .C(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__o21a_1 _29093_ (.A1(net108),
    .A2(_24727_),
    .B1(_00592_),
    .X(_00594_));
 sky130_fd_sc_hd__o21a_1 _29094_ (.A1(_24540_),
    .A2(_24614_),
    .B1(_24612_),
    .X(_00595_));
 sky130_fd_sc_hd__o21ai_1 _29095_ (.A1(_00593_),
    .A2(_00594_),
    .B1(_00595_),
    .Y(_00596_));
 sky130_fd_sc_hd__inv_2 _29096_ (.A(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hd__nor3_1 _29097_ (.A(_00595_),
    .B(_00593_),
    .C(_00594_),
    .Y(_00598_));
 sky130_fd_sc_hd__o21a_2 _29098_ (.A1(_24729_),
    .A2(_24854_),
    .B1(_24850_),
    .X(_00599_));
 sky130_fd_sc_hd__a21oi_1 _29099_ (.A1(_07338_),
    .A2(_07580_),
    .B1(_07569_),
    .Y(_00600_));
 sky130_fd_sc_hd__o211a_1 _29100_ (.A1(_23995_),
    .A2(_07580_),
    .B1(_16525_),
    .C1(_16514_),
    .X(_00602_));
 sky130_fd_sc_hd__nand3_1 _29101_ (.A(_24638_),
    .B(_24640_),
    .C(_24637_),
    .Y(_00603_));
 sky130_fd_sc_hd__nor2_1 _29102_ (.A(_07316_),
    .B(_18359_),
    .Y(_00604_));
 sky130_fd_sc_hd__and2_1 _29103_ (.A(_18358_),
    .B(_21419_),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _29104_ (.A(_16525_),
    .B(_16514_),
    .Y(_00606_));
 sky130_fd_sc_hd__a21oi_2 _29105_ (.A1(_00606_),
    .A2(_07294_),
    .B1(_20528_),
    .Y(_00607_));
 sky130_fd_sc_hd__o21bai_1 _29106_ (.A1(_00604_),
    .A2(_00605_),
    .B1_N(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _29107_ (.A(_18359_),
    .B(_07316_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand3b_1 _29108_ (.A_N(_00604_),
    .B(_00609_),
    .C(_00607_),
    .Y(_00610_));
 sky130_fd_sc_hd__a21bo_1 _29109_ (.A1(_24631_),
    .A2(_18348_),
    .B1_N(_24632_),
    .X(_00611_));
 sky130_fd_sc_hd__clkbuf_2 _29110_ (.A(net358),
    .X(_00613_));
 sky130_fd_sc_hd__nor2_1 _29111_ (.A(_24628_),
    .B(_00613_),
    .Y(_00614_));
 sky130_fd_sc_hd__and2_1 _29112_ (.A(\delay_line[21][9] ),
    .B(net358),
    .X(_00615_));
 sky130_fd_sc_hd__nand2_2 _29113_ (.A(\delay_line[21][8] ),
    .B(_24628_),
    .Y(_00616_));
 sky130_fd_sc_hd__o21ai_1 _29114_ (.A1(_00614_),
    .A2(_00615_),
    .B1(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__or2_1 _29115_ (.A(_00613_),
    .B(_00616_),
    .X(_00618_));
 sky130_fd_sc_hd__a21o_1 _29116_ (.A1(_00617_),
    .A2(_00618_),
    .B1(_21412_),
    .X(_00619_));
 sky130_fd_sc_hd__o211ai_2 _29117_ (.A1(_00613_),
    .A2(_00616_),
    .B1(_21412_),
    .C1(_00617_),
    .Y(_00620_));
 sky130_fd_sc_hd__clkbuf_2 _29118_ (.A(_00620_),
    .X(_00621_));
 sky130_fd_sc_hd__nand3_1 _29119_ (.A(_00611_),
    .B(_00619_),
    .C(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__a21o_1 _29120_ (.A1(_00619_),
    .A2(_00621_),
    .B1(_00611_),
    .X(_00624_));
 sky130_fd_sc_hd__nand4_1 _29121_ (.A(_00608_),
    .B(_00610_),
    .C(_00622_),
    .D(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__and3_1 _29122_ (.A(_00611_),
    .B(_00619_),
    .C(_00620_),
    .X(_00626_));
 sky130_fd_sc_hd__a21oi_1 _29123_ (.A1(_00619_),
    .A2(_00621_),
    .B1(_00611_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _29124_ (.A(_00608_),
    .B(_00610_),
    .Y(_00628_));
 sky130_fd_sc_hd__o21ai_1 _29125_ (.A1(_00626_),
    .A2(_00627_),
    .B1(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand4_1 _29126_ (.A(_24637_),
    .B(_00603_),
    .C(_00625_),
    .D(_00629_),
    .Y(_00630_));
 sky130_fd_sc_hd__a22o_1 _29127_ (.A1(_24637_),
    .A2(_00603_),
    .B1(_00625_),
    .B2(_00629_),
    .X(_00631_));
 sky130_fd_sc_hd__a2bb2o_1 _29128_ (.A1_N(_00600_),
    .A2_N(_00602_),
    .B1(_00630_),
    .B2(_00631_),
    .X(_00632_));
 sky130_fd_sc_hd__or2_1 _29129_ (.A(_00600_),
    .B(_00602_),
    .X(_00633_));
 sky130_fd_sc_hd__nand3b_1 _29130_ (.A_N(_00633_),
    .B(_00630_),
    .C(_00631_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _29131_ (.A(_24645_),
    .B(_24647_),
    .Y(_00636_));
 sky130_fd_sc_hd__a21o_1 _29132_ (.A1(_00632_),
    .A2(_00635_),
    .B1(_00636_),
    .X(_00637_));
 sky130_fd_sc_hd__nand3_1 _29133_ (.A(_00632_),
    .B(_00635_),
    .C(_00636_),
    .Y(_00638_));
 sky130_fd_sc_hd__a32o_1 _29134_ (.A1(_24017_),
    .A2(_16492_),
    .A3(_07602_),
    .B1(_00637_),
    .B2(_00638_),
    .X(_00639_));
 sky130_fd_sc_hd__nand3_1 _29135_ (.A(_00637_),
    .B(_00638_),
    .C(_07613_),
    .Y(_00640_));
 sky130_fd_sc_hd__inv_2 _29136_ (.A(_24649_),
    .Y(_00641_));
 sky130_fd_sc_hd__o211a_1 _29137_ (.A1(_22994_),
    .A2(_22998_),
    .B1(_23001_),
    .C1(_22982_),
    .X(_00642_));
 sky130_fd_sc_hd__and3_1 _29138_ (.A(_00640_),
    .B(_00641_),
    .C(_00642_),
    .X(_00643_));
 sky130_fd_sc_hd__a22oi_2 _29139_ (.A1(_00642_),
    .A2(_00641_),
    .B1(_00639_),
    .B2(_00640_),
    .Y(_00644_));
 sky130_fd_sc_hd__a21oi_2 _29140_ (.A1(_00639_),
    .A2(_00643_),
    .B1(_00644_),
    .Y(_00646_));
 sky130_fd_sc_hd__and4b_1 _29141_ (.A_N(_23003_),
    .B(_21434_),
    .C(_21432_),
    .D(_21431_),
    .X(_00647_));
 sky130_fd_sc_hd__a22oi_4 _29142_ (.A1(_00647_),
    .A2(_00641_),
    .B1(_24650_),
    .B2(_24651_),
    .Y(_00648_));
 sky130_fd_sc_hd__xnor2_4 _29143_ (.A(_00646_),
    .B(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__nor2_1 _29144_ (.A(_16393_),
    .B(_16415_),
    .Y(_00650_));
 sky130_fd_sc_hd__a22oi_2 _29145_ (.A1(_01644_),
    .A2(_22964_),
    .B1(_00650_),
    .B2(_16448_),
    .Y(_00651_));
 sky130_fd_sc_hd__a22oi_2 _29146_ (.A1(_24661_),
    .A2(_22949_),
    .B1(_24659_),
    .B2(_18374_),
    .Y(_00652_));
 sky130_fd_sc_hd__nor2_1 _29147_ (.A(_24654_),
    .B(\delay_line[19][10] ),
    .Y(_00653_));
 sky130_fd_sc_hd__and2_1 _29148_ (.A(\delay_line[19][9] ),
    .B(\delay_line[19][10] ),
    .X(_00654_));
 sky130_fd_sc_hd__nand2_1 _29149_ (.A(_22948_),
    .B(_24654_),
    .Y(_00655_));
 sky130_fd_sc_hd__o21ai_1 _29150_ (.A1(_00653_),
    .A2(_00654_),
    .B1(_00655_),
    .Y(_00657_));
 sky130_fd_sc_hd__buf_1 _29151_ (.A(\delay_line[19][10] ),
    .X(_00658_));
 sky130_fd_sc_hd__or2_1 _29152_ (.A(_00658_),
    .B(_00655_),
    .X(_00659_));
 sky130_fd_sc_hd__buf_1 _29153_ (.A(_19402_),
    .X(_00660_));
 sky130_fd_sc_hd__a21o_1 _29154_ (.A1(_00657_),
    .A2(_00659_),
    .B1(_00660_),
    .X(_00661_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29155_ (.A(_00658_),
    .X(_00662_));
 sky130_fd_sc_hd__buf_1 _29156_ (.A(_00657_),
    .X(_00663_));
 sky130_fd_sc_hd__o211ai_1 _29157_ (.A1(_00662_),
    .A2(_00655_),
    .B1(_00660_),
    .C1(_00663_),
    .Y(_00664_));
 sky130_fd_sc_hd__nand3b_1 _29158_ (.A_N(_00652_),
    .B(_00661_),
    .C(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__buf_1 _29159_ (.A(_00665_),
    .X(_00666_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29160_ (.A(_00660_),
    .X(_00668_));
 sky130_fd_sc_hd__a21oi_1 _29161_ (.A1(_00663_),
    .A2(_00659_),
    .B1(_00668_),
    .Y(_00669_));
 sky130_fd_sc_hd__and3_1 _29162_ (.A(_00663_),
    .B(_00659_),
    .C(_00660_),
    .X(_00670_));
 sky130_fd_sc_hd__o21ai_2 _29163_ (.A1(_00669_),
    .A2(_00670_),
    .B1(_00652_),
    .Y(_00671_));
 sky130_fd_sc_hd__o21a_1 _29164_ (.A1(_16393_),
    .A2(_16415_),
    .B1(_07360_),
    .X(_00672_));
 sky130_fd_sc_hd__nand3_1 _29165_ (.A(_16371_),
    .B(_18371_),
    .C(_18372_),
    .Y(_00673_));
 sky130_fd_sc_hd__a21o_1 _29166_ (.A1(_18371_),
    .A2(_18372_),
    .B1(_16371_),
    .X(_00674_));
 sky130_fd_sc_hd__nand2_1 _29167_ (.A(_00673_),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__o21ai_1 _29168_ (.A1(_18377_),
    .A2(_00672_),
    .B1(_00675_),
    .Y(_00676_));
 sky130_fd_sc_hd__o2111ai_1 _29169_ (.A1(_01644_),
    .A2(_00650_),
    .B1(_19410_),
    .C1(_00673_),
    .D1(_00674_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _29170_ (.A(_00676_),
    .B(_00677_),
    .Y(_00679_));
 sky130_fd_sc_hd__a21oi_1 _29171_ (.A1(_00666_),
    .A2(_00671_),
    .B1(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__and3_1 _29172_ (.A(_00679_),
    .B(_00666_),
    .C(_00671_),
    .X(_00681_));
 sky130_fd_sc_hd__a21boi_1 _29173_ (.A1(_24669_),
    .A2(_24671_),
    .B1_N(_24665_),
    .Y(_00682_));
 sky130_fd_sc_hd__o21ai_2 _29174_ (.A1(_00680_),
    .A2(_00681_),
    .B1(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__a21o_1 _29175_ (.A1(_00666_),
    .A2(_00671_),
    .B1(_00679_),
    .X(_00684_));
 sky130_fd_sc_hd__nand3_1 _29176_ (.A(_00679_),
    .B(_00665_),
    .C(_00671_),
    .Y(_00685_));
 sky130_fd_sc_hd__nand3b_1 _29177_ (.A_N(_00682_),
    .B(_00684_),
    .C(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand3b_2 _29178_ (.A_N(_00651_),
    .B(_00683_),
    .C(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hd__a21bo_1 _29179_ (.A1(_00683_),
    .A2(_00686_),
    .B1_N(_00651_),
    .X(_00688_));
 sky130_fd_sc_hd__a22oi_2 _29180_ (.A1(_24680_),
    .A2(_24681_),
    .B1(_00687_),
    .B2(_00688_),
    .Y(_00690_));
 sky130_fd_sc_hd__nand4_2 _29181_ (.A(_24680_),
    .B(_24681_),
    .C(_00687_),
    .D(_00688_),
    .Y(_00691_));
 sky130_fd_sc_hd__nand2_1 _29182_ (.A(_00691_),
    .B(_07492_),
    .Y(_00692_));
 sky130_fd_sc_hd__or2_1 _29183_ (.A(_00690_),
    .B(_00692_),
    .X(_00693_));
 sky130_fd_sc_hd__a221o_1 _29184_ (.A1(_22942_),
    .A2(_22943_),
    .B1(_22966_),
    .B2(_22967_),
    .C1(_24683_),
    .X(_00694_));
 sky130_fd_sc_hd__a22o_1 _29185_ (.A1(_24680_),
    .A2(_24681_),
    .B1(_00687_),
    .B2(_00688_),
    .X(_00695_));
 sky130_fd_sc_hd__a21oi_1 _29186_ (.A1(_00691_),
    .A2(_00695_),
    .B1(_07492_),
    .Y(_00696_));
 sky130_fd_sc_hd__nor2_1 _29187_ (.A(_00694_),
    .B(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__and3_1 _29188_ (.A(_00695_),
    .B(_07481_),
    .C(_00691_),
    .X(_00698_));
 sky130_fd_sc_hd__o21ai_1 _29189_ (.A1(_00696_),
    .A2(_00698_),
    .B1(_00694_),
    .Y(_00699_));
 sky130_fd_sc_hd__a21bo_1 _29190_ (.A1(_00693_),
    .A2(_00697_),
    .B1_N(_00699_),
    .X(_00701_));
 sky130_fd_sc_hd__a221o_1 _29191_ (.A1(_20563_),
    .A2(_20565_),
    .B1(_21389_),
    .B2(_21390_),
    .C1(_24718_),
    .X(_00702_));
 sky130_fd_sc_hd__o22ai_2 _29192_ (.A1(_24683_),
    .A2(_00702_),
    .B1(_24685_),
    .B2(_24720_),
    .Y(_00703_));
 sky130_fd_sc_hd__and2b_1 _29193_ (.A_N(_00701_),
    .B(_00703_),
    .X(_00704_));
 sky130_fd_sc_hd__o221a_1 _29194_ (.A1(_24683_),
    .A2(_00702_),
    .B1(_24685_),
    .B2(_24720_),
    .C1(_00701_),
    .X(_00705_));
 sky130_fd_sc_hd__a31oi_2 _29195_ (.A1(_24709_),
    .A2(_24712_),
    .A3(_24714_),
    .B1(_24723_),
    .Y(_00706_));
 sky130_fd_sc_hd__and3_1 _29196_ (.A(_24712_),
    .B(_22937_),
    .C(_24709_),
    .X(_00707_));
 sky130_fd_sc_hd__nand2_1 _29197_ (.A(_21357_),
    .B(net374),
    .Y(_00708_));
 sky130_fd_sc_hd__or2_1 _29198_ (.A(net375),
    .B(_00708_),
    .X(_00709_));
 sky130_fd_sc_hd__o21ai_2 _29199_ (.A1(\delay_line[18][1] ),
    .A2(_21355_),
    .B1(_16327_),
    .Y(_00710_));
 sky130_fd_sc_hd__buf_2 _29200_ (.A(net373),
    .X(_00712_));
 sky130_fd_sc_hd__o211ai_4 _29201_ (.A1(_21362_),
    .A2(_00712_),
    .B1(_24694_),
    .C1(_19390_),
    .Y(_00713_));
 sky130_fd_sc_hd__a21o_1 _29202_ (.A1(_20542_),
    .A2(_00712_),
    .B1(_00713_),
    .X(_00714_));
 sky130_fd_sc_hd__and2_2 _29203_ (.A(\delay_line[18][6] ),
    .B(net373),
    .X(_00715_));
 sky130_fd_sc_hd__nor2_1 _29204_ (.A(_21362_),
    .B(_00712_),
    .Y(_00716_));
 sky130_fd_sc_hd__o21ai_2 _29205_ (.A1(_00715_),
    .A2(_00716_),
    .B1(_24695_),
    .Y(_00717_));
 sky130_fd_sc_hd__a22o_1 _29206_ (.A1(_00709_),
    .A2(_00710_),
    .B1(_00714_),
    .B2(_00717_),
    .X(_00718_));
 sky130_fd_sc_hd__o2111ai_4 _29207_ (.A1(_00713_),
    .A2(_00715_),
    .B1(_00710_),
    .C1(_00709_),
    .D1(_00717_),
    .Y(_00719_));
 sky130_fd_sc_hd__nand2_1 _29208_ (.A(_24696_),
    .B(_24700_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand3_2 _29209_ (.A(_00718_),
    .B(_00719_),
    .C(_00720_),
    .Y(_00721_));
 sky130_fd_sc_hd__a21o_1 _29210_ (.A1(_00718_),
    .A2(_00719_),
    .B1(_00720_),
    .X(_00723_));
 sky130_fd_sc_hd__o2111ai_4 _29211_ (.A1(_23940_),
    .A2(_07525_),
    .B1(_01677_),
    .C1(_00721_),
    .D1(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__and3_1 _29212_ (.A(_21355_),
    .B(_01677_),
    .C(_23852_),
    .X(_00725_));
 sky130_fd_sc_hd__o2bb2ai_1 _29213_ (.A1_N(_00723_),
    .A2_N(_00721_),
    .B1(_19393_),
    .B2(_00725_),
    .Y(_00726_));
 sky130_fd_sc_hd__o21ai_1 _29214_ (.A1(_23951_),
    .A2(_24707_),
    .B1(_24708_),
    .Y(_00727_));
 sky130_fd_sc_hd__a21oi_1 _29215_ (.A1(_00724_),
    .A2(_00726_),
    .B1(_00727_),
    .Y(_00728_));
 sky130_fd_sc_hd__and3_1 _29216_ (.A(_00727_),
    .B(_00724_),
    .C(_00726_),
    .X(_00729_));
 sky130_fd_sc_hd__nor2_1 _29217_ (.A(_00728_),
    .B(_00729_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _29218_ (.A(_00707_),
    .B(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__o22ai_1 _29219_ (.A1(_24690_),
    .A2(_24715_),
    .B1(_00728_),
    .B2(_00729_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand2_1 _29220_ (.A(_00731_),
    .B(_00732_),
    .Y(_00734_));
 sky130_fd_sc_hd__xnor2_1 _29221_ (.A(_00706_),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__o21ai_1 _29222_ (.A1(_00704_),
    .A2(_00705_),
    .B1(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__or3_1 _29223_ (.A(_00705_),
    .B(_00735_),
    .C(_00704_),
    .X(_00737_));
 sky130_fd_sc_hd__and2_2 _29224_ (.A(_00736_),
    .B(_00737_),
    .X(_00738_));
 sky130_fd_sc_hd__xnor2_4 _29225_ (.A(_00649_),
    .B(_00738_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand3_1 _29226_ (.A(_24791_),
    .B(_24794_),
    .C(_24789_),
    .Y(_00740_));
 sky130_fd_sc_hd__a21oi_1 _29227_ (.A1(_18407_),
    .A2(_19451_),
    .B1(_07184_),
    .Y(_00741_));
 sky130_fd_sc_hd__and3_2 _29228_ (.A(_07173_),
    .B(_18406_),
    .C(_19451_),
    .X(_00742_));
 sky130_fd_sc_hd__nor2_1 _29229_ (.A(net391),
    .B(\delay_line[14][6] ),
    .Y(_00743_));
 sky130_fd_sc_hd__and2_1 _29230_ (.A(net391),
    .B(\delay_line[14][6] ),
    .X(_00745_));
 sky130_fd_sc_hd__o21bai_1 _29231_ (.A1(_00743_),
    .A2(_00745_),
    .B1_N(\delay_line[14][10] ),
    .Y(_00746_));
 sky130_fd_sc_hd__a21oi_1 _29232_ (.A1(_18406_),
    .A2(_19450_),
    .B1(_24784_),
    .Y(_00747_));
 sky130_fd_sc_hd__nand2_1 _29233_ (.A(_19450_),
    .B(_20587_),
    .Y(_00748_));
 sky130_fd_sc_hd__clkbuf_2 _29234_ (.A(\delay_line[14][10] ),
    .X(_00749_));
 sky130_fd_sc_hd__nand3b_1 _29235_ (.A_N(_00743_),
    .B(_00748_),
    .C(_00749_),
    .Y(_00750_));
 sky130_fd_sc_hd__and3_1 _29236_ (.A(_00746_),
    .B(_00747_),
    .C(_00750_),
    .X(_00751_));
 sky130_fd_sc_hd__o2bb2a_1 _29237_ (.A1_N(_00750_),
    .A2_N(_00746_),
    .B1(_24782_),
    .B2(_24784_),
    .X(_00752_));
 sky130_fd_sc_hd__nor4_1 _29238_ (.A(_00741_),
    .B(_00742_),
    .C(_00751_),
    .D(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hd__o22a_1 _29239_ (.A1(_00741_),
    .A2(_00742_),
    .B1(_00751_),
    .B2(_00752_),
    .X(_00754_));
 sky130_fd_sc_hd__a211o_1 _29240_ (.A1(_24789_),
    .A2(_00740_),
    .B1(net258),
    .C1(_00754_),
    .X(_00756_));
 sky130_fd_sc_hd__o211ai_2 _29241_ (.A1(net258),
    .A2(_00754_),
    .B1(_24789_),
    .C1(_00740_),
    .Y(_00757_));
 sky130_fd_sc_hd__nand4_2 _29242_ (.A(_00756_),
    .B(_01776_),
    .C(_00757_),
    .D(_23050_),
    .Y(_00758_));
 sky130_fd_sc_hd__a32o_1 _29243_ (.A1(_01776_),
    .A2(_16843_),
    .A3(_18408_),
    .B1(_00757_),
    .B2(_00756_),
    .X(_00759_));
 sky130_fd_sc_hd__nand2_1 _29244_ (.A(_24799_),
    .B(_24801_),
    .Y(_00760_));
 sky130_fd_sc_hd__a21oi_2 _29245_ (.A1(_00758_),
    .A2(_00759_),
    .B1(_00760_),
    .Y(_00761_));
 sky130_fd_sc_hd__and3_1 _29246_ (.A(_00760_),
    .B(_00758_),
    .C(_00759_),
    .X(_00762_));
 sky130_fd_sc_hd__a21oi_2 _29247_ (.A1(_24781_),
    .A2(_24804_),
    .B1(_24803_),
    .Y(_00763_));
 sky130_fd_sc_hd__nor3_2 _29248_ (.A(_00761_),
    .B(_00762_),
    .C(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__o21a_1 _29249_ (.A1(_00761_),
    .A2(_00762_),
    .B1(_00763_),
    .X(_00765_));
 sky130_fd_sc_hd__a21oi_1 _29250_ (.A1(_24757_),
    .A2(_24758_),
    .B1(_24730_),
    .Y(_00767_));
 sky130_fd_sc_hd__a31oi_1 _29251_ (.A1(_24759_),
    .A2(_24760_),
    .A3(_24094_),
    .B1(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__clkbuf_2 _29252_ (.A(_07107_),
    .X(_00769_));
 sky130_fd_sc_hd__a21oi_1 _29253_ (.A1(_24744_),
    .A2(_24747_),
    .B1(_24748_),
    .Y(_00770_));
 sky130_fd_sc_hd__o21ai_1 _29254_ (.A1(_24733_),
    .A2(_00770_),
    .B1(_24749_),
    .Y(_00771_));
 sky130_fd_sc_hd__nor2_1 _29255_ (.A(_07074_),
    .B(_16689_),
    .Y(_00772_));
 sky130_fd_sc_hd__and3_1 _29256_ (.A(_16700_),
    .B(_16744_),
    .C(_07096_),
    .X(_00773_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29257_ (.A(\delay_line[15][11] ),
    .X(_00774_));
 sky130_fd_sc_hd__and2_1 _29258_ (.A(\delay_line[15][9] ),
    .B(_00774_),
    .X(_00775_));
 sky130_fd_sc_hd__o211ai_2 _29259_ (.A1(_23078_),
    .A2(_00774_),
    .B1(_24737_),
    .C1(_21452_),
    .Y(_00776_));
 sky130_fd_sc_hd__nor2_1 _29260_ (.A(_23078_),
    .B(_00774_),
    .Y(_00778_));
 sky130_fd_sc_hd__o21bai_2 _29261_ (.A1(_00775_),
    .A2(_00778_),
    .B1_N(_24734_),
    .Y(_00779_));
 sky130_fd_sc_hd__o211a_1 _29262_ (.A1(_00775_),
    .A2(_00776_),
    .B1(_19461_),
    .C1(_00779_),
    .X(_00780_));
 sky130_fd_sc_hd__buf_1 _29263_ (.A(_00774_),
    .X(_00781_));
 sky130_fd_sc_hd__a21o_1 _29264_ (.A1(_23076_),
    .A2(_00781_),
    .B1(_00776_),
    .X(_00782_));
 sky130_fd_sc_hd__a21o_1 _29265_ (.A1(_00782_),
    .A2(_00779_),
    .B1(_21458_),
    .X(_00783_));
 sky130_fd_sc_hd__a2bb2o_1 _29266_ (.A1_N(_24735_),
    .A2_N(_24738_),
    .B1(_18422_),
    .B2(_24742_),
    .X(_00784_));
 sky130_fd_sc_hd__nand3b_4 _29267_ (.A_N(_00780_),
    .B(_00783_),
    .C(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__a21oi_2 _29268_ (.A1(_00782_),
    .A2(_00779_),
    .B1(_21458_),
    .Y(_00786_));
 sky130_fd_sc_hd__o31a_1 _29269_ (.A1(_23082_),
    .A2(_24735_),
    .A3(_24741_),
    .B1(_24744_),
    .X(_00787_));
 sky130_fd_sc_hd__o21ai_4 _29270_ (.A1(_00780_),
    .A2(_00786_),
    .B1(_00787_),
    .Y(_00789_));
 sky130_fd_sc_hd__o211ai_2 _29271_ (.A1(_00772_),
    .A2(_00773_),
    .B1(_00785_),
    .C1(_00789_),
    .Y(_00790_));
 sky130_fd_sc_hd__a31o_1 _29272_ (.A1(_16711_),
    .A2(_16755_),
    .A3(_07096_),
    .B1(_00772_),
    .X(_00791_));
 sky130_fd_sc_hd__a21o_1 _29273_ (.A1(_00785_),
    .A2(_00789_),
    .B1(_00791_),
    .X(_00792_));
 sky130_fd_sc_hd__nand3_2 _29274_ (.A(_00771_),
    .B(_00790_),
    .C(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hd__o211a_1 _29275_ (.A1(_00772_),
    .A2(_00773_),
    .B1(_00785_),
    .C1(_00789_),
    .X(_00794_));
 sky130_fd_sc_hd__a21oi_1 _29276_ (.A1(_00785_),
    .A2(_00789_),
    .B1(_00791_),
    .Y(_00795_));
 sky130_fd_sc_hd__o21bai_4 _29277_ (.A1(_00794_),
    .A2(_00795_),
    .B1_N(_00771_),
    .Y(_00796_));
 sky130_fd_sc_hd__o2111ai_4 _29278_ (.A1(_24763_),
    .A2(_00769_),
    .B1(_01820_),
    .C1(_00793_),
    .D1(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hd__buf_1 _29279_ (.A(_16722_),
    .X(_00798_));
 sky130_fd_sc_hd__or3_1 _29280_ (.A(_07107_),
    .B(_00798_),
    .C(_24763_),
    .X(_00800_));
 sky130_fd_sc_hd__a22o_1 _29281_ (.A1(_01820_),
    .A2(_00800_),
    .B1(_00796_),
    .B2(_00793_),
    .X(_00801_));
 sky130_fd_sc_hd__nand3b_2 _29282_ (.A_N(_00768_),
    .B(_00797_),
    .C(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__buf_1 _29283_ (.A(_00793_),
    .X(_00803_));
 sky130_fd_sc_hd__o21ai_1 _29284_ (.A1(_00769_),
    .A2(_24763_),
    .B1(_01820_),
    .Y(_00804_));
 sky130_fd_sc_hd__a21o_1 _29285_ (.A1(_00796_),
    .A2(_00803_),
    .B1(_00804_),
    .X(_00805_));
 sky130_fd_sc_hd__o211ai_1 _29286_ (.A1(_07129_),
    .A2(_00798_),
    .B1(_00803_),
    .C1(_00796_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand3_1 _29287_ (.A(_00805_),
    .B(_00806_),
    .C(_00768_),
    .Y(_00807_));
 sky130_fd_sc_hd__nand3_1 _29288_ (.A(_00802_),
    .B(_00807_),
    .C(_24762_),
    .Y(_00808_));
 sky130_fd_sc_hd__clkbuf_2 _29289_ (.A(_00808_),
    .X(_00809_));
 sky130_fd_sc_hd__a21o_1 _29290_ (.A1(_00802_),
    .A2(_00807_),
    .B1(_24762_),
    .X(_00811_));
 sky130_fd_sc_hd__and4b_1 _29291_ (.A_N(_24769_),
    .B(_24761_),
    .C(_24764_),
    .D(_00811_),
    .X(_00812_));
 sky130_fd_sc_hd__a2bb2o_1 _29292_ (.A1_N(_24766_),
    .A2_N(_24769_),
    .B1(_00808_),
    .B2(_00811_),
    .X(_00813_));
 sky130_fd_sc_hd__a21bo_1 _29293_ (.A1(_00809_),
    .A2(_00812_),
    .B1_N(_00813_),
    .X(_00814_));
 sky130_fd_sc_hd__a21oi_1 _29294_ (.A1(_24771_),
    .A2(_24780_),
    .B1(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__and3_1 _29295_ (.A(_24771_),
    .B(_24780_),
    .C(_00814_),
    .X(_00816_));
 sky130_fd_sc_hd__nor4_1 _29296_ (.A(_00764_),
    .B(_00765_),
    .C(_00815_),
    .D(_00816_),
    .Y(_00817_));
 sky130_fd_sc_hd__o22a_1 _29297_ (.A1(_00764_),
    .A2(_00765_),
    .B1(_00815_),
    .B2(_00816_),
    .X(_00818_));
 sky130_fd_sc_hd__nor2_1 _29298_ (.A(net102),
    .B(_00818_),
    .Y(_00819_));
 sky130_fd_sc_hd__nor2_1 _29299_ (.A(_24847_),
    .B(_24846_),
    .Y(_00820_));
 sky130_fd_sc_hd__a21oi_1 _29300_ (.A1(_24823_),
    .A2(_24824_),
    .B1(_23030_),
    .Y(_00822_));
 sky130_fd_sc_hd__o21ai_1 _29301_ (.A1(_24812_),
    .A2(_00822_),
    .B1(_24828_),
    .Y(_00823_));
 sky130_fd_sc_hd__mux2_1 _29302_ (.A0(_24813_),
    .A1(_24817_),
    .S(_18400_),
    .X(_00824_));
 sky130_fd_sc_hd__and2_1 _29303_ (.A(net385),
    .B(net384),
    .X(_00825_));
 sky130_fd_sc_hd__clkbuf_2 _29304_ (.A(_00825_),
    .X(_00826_));
 sky130_fd_sc_hd__o21ai_1 _29305_ (.A1(_24816_),
    .A2(_21516_),
    .B1(_23016_),
    .Y(_00827_));
 sky130_fd_sc_hd__clkbuf_2 _29306_ (.A(net382),
    .X(_00828_));
 sky130_fd_sc_hd__nor2_1 _29307_ (.A(_24816_),
    .B(_21516_),
    .Y(_00829_));
 sky130_fd_sc_hd__o21bai_2 _29308_ (.A1(_00825_),
    .A2(_00829_),
    .B1_N(_23016_),
    .Y(_00830_));
 sky130_fd_sc_hd__o211a_1 _29309_ (.A1(_00826_),
    .A2(_00827_),
    .B1(_00828_),
    .C1(_00830_),
    .X(_00831_));
 sky130_fd_sc_hd__a21o_1 _29310_ (.A1(_20630_),
    .A2(_21516_),
    .B1(_00827_),
    .X(_00833_));
 sky130_fd_sc_hd__clkbuf_2 _29311_ (.A(_00828_),
    .X(_00834_));
 sky130_fd_sc_hd__a21oi_1 _29312_ (.A1(_00833_),
    .A2(_00830_),
    .B1(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__o21bai_1 _29313_ (.A1(_00831_),
    .A2(_00835_),
    .B1_N(_24822_),
    .Y(_00836_));
 sky130_fd_sc_hd__clkbuf_2 _29314_ (.A(_00827_),
    .X(_00837_));
 sky130_fd_sc_hd__o211ai_2 _29315_ (.A1(_00826_),
    .A2(_00837_),
    .B1(_00834_),
    .C1(_00830_),
    .Y(_00838_));
 sky130_fd_sc_hd__a21o_1 _29316_ (.A1(_00833_),
    .A2(_00830_),
    .B1(_00828_),
    .X(_00839_));
 sky130_fd_sc_hd__nand3_1 _29317_ (.A(_24823_),
    .B(_00838_),
    .C(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hd__nand3b_1 _29318_ (.A_N(_00824_),
    .B(_00836_),
    .C(_00840_),
    .Y(_00841_));
 sky130_fd_sc_hd__o21ai_1 _29319_ (.A1(_00831_),
    .A2(_00835_),
    .B1(_24822_),
    .Y(_00842_));
 sky130_fd_sc_hd__nand3b_1 _29320_ (.A_N(_24822_),
    .B(_00838_),
    .C(_00839_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand3_1 _29321_ (.A(_00842_),
    .B(_00824_),
    .C(_00844_),
    .Y(_00845_));
 sky130_fd_sc_hd__nand3_1 _29322_ (.A(_00823_),
    .B(_00841_),
    .C(_00845_),
    .Y(_00846_));
 sky130_fd_sc_hd__buf_1 _29323_ (.A(_00846_),
    .X(_00847_));
 sky130_fd_sc_hd__a21o_1 _29324_ (.A1(_00841_),
    .A2(_00845_),
    .B1(_00823_),
    .X(_00848_));
 sky130_fd_sc_hd__o211a_1 _29325_ (.A1(_24835_),
    .A2(_19441_),
    .B1(_01875_),
    .C1(_16612_),
    .X(_00849_));
 sky130_fd_sc_hd__o21a_1 _29326_ (.A1(_18400_),
    .A2(_19441_),
    .B1(_16601_),
    .X(_00850_));
 sky130_fd_sc_hd__nor2_1 _29327_ (.A(_01875_),
    .B(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__nor2_1 _29328_ (.A(_00849_),
    .B(_00851_),
    .Y(_00852_));
 sky130_fd_sc_hd__a21bo_1 _29329_ (.A1(_00847_),
    .A2(_00848_),
    .B1_N(_00852_),
    .X(_00853_));
 sky130_fd_sc_hd__o211ai_1 _29330_ (.A1(_00849_),
    .A2(_00851_),
    .B1(_00847_),
    .C1(_00848_),
    .Y(_00855_));
 sky130_fd_sc_hd__nand4_1 _29331_ (.A(_24839_),
    .B(_24840_),
    .C(_00853_),
    .D(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__o21ai_1 _29332_ (.A1(_24833_),
    .A2(_24832_),
    .B1(_24840_),
    .Y(_00857_));
 sky130_fd_sc_hd__nand3_1 _29333_ (.A(_00848_),
    .B(_00852_),
    .C(_00847_),
    .Y(_00858_));
 sky130_fd_sc_hd__a2bb2o_1 _29334_ (.A1_N(_00849_),
    .A2_N(_00851_),
    .B1(_00847_),
    .B2(_00848_),
    .X(_00859_));
 sky130_fd_sc_hd__nand3_1 _29335_ (.A(_00857_),
    .B(_00858_),
    .C(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__and3_1 _29336_ (.A(_00856_),
    .B(_00860_),
    .C(_24836_),
    .X(_00861_));
 sky130_fd_sc_hd__o2bb2a_1 _29337_ (.A1_N(_00856_),
    .A2_N(_00860_),
    .B1(_16645_),
    .B2(_21515_),
    .X(_00862_));
 sky130_fd_sc_hd__nor2_2 _29338_ (.A(_00861_),
    .B(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__o21ai_1 _29339_ (.A1(_24845_),
    .A2(_00820_),
    .B1(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__a311o_1 _29340_ (.A1(_24843_),
    .A2(_24840_),
    .A3(_24841_),
    .B1(_00820_),
    .C1(_00863_),
    .X(_00866_));
 sky130_fd_sc_hd__and3_1 _29341_ (.A(_00819_),
    .B(_00864_),
    .C(_00866_),
    .X(_00867_));
 sky130_fd_sc_hd__o2bb2a_1 _29342_ (.A1_N(_00866_),
    .A2_N(_00864_),
    .B1(net102),
    .B2(_00818_),
    .X(_00868_));
 sky130_fd_sc_hd__nand2_1 _29343_ (.A(_24811_),
    .B(_24848_),
    .Y(_00869_));
 sky130_fd_sc_hd__o211ai_2 _29344_ (.A1(_00867_),
    .A2(_00868_),
    .B1(_24808_),
    .C1(_00869_),
    .Y(_00870_));
 sky130_fd_sc_hd__a211o_2 _29345_ (.A1(_24808_),
    .A2(_00869_),
    .B1(_00867_),
    .C1(_00868_),
    .X(_00871_));
 sky130_fd_sc_hd__nand2_4 _29346_ (.A(_00870_),
    .B(_00871_),
    .Y(_00872_));
 sky130_fd_sc_hd__xnor2_4 _29347_ (.A(_00739_),
    .B(_00872_),
    .Y(_00873_));
 sky130_fd_sc_hd__xnor2_1 _29348_ (.A(_00599_),
    .B(_00873_),
    .Y(_00874_));
 sky130_fd_sc_hd__nor3_1 _29349_ (.A(_00597_),
    .B(_00598_),
    .C(_00874_),
    .Y(_00875_));
 sky130_fd_sc_hd__o21a_1 _29350_ (.A1(_00597_),
    .A2(_00598_),
    .B1(_00874_),
    .X(_00877_));
 sky130_fd_sc_hd__a21oi_1 _29351_ (.A1(_24621_),
    .A2(_24858_),
    .B1(_24857_),
    .Y(_00878_));
 sky130_fd_sc_hd__o21ai_1 _29352_ (.A1(_00875_),
    .A2(_00877_),
    .B1(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hd__or3_1 _29353_ (.A(_00878_),
    .B(_00875_),
    .C(_00877_),
    .X(_00880_));
 sky130_fd_sc_hd__nand2_1 _29354_ (.A(_00879_),
    .B(_00880_),
    .Y(_00881_));
 sky130_fd_sc_hd__o21ai_2 _29355_ (.A1(_23221_),
    .A2(_24473_),
    .B1(_24472_),
    .Y(_00882_));
 sky130_fd_sc_hd__nor2_1 _29356_ (.A(_24453_),
    .B(net316),
    .Y(_00883_));
 sky130_fd_sc_hd__buf_1 _29357_ (.A(\delay_line[31][10] ),
    .X(_00884_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29358_ (.A(net316),
    .X(_00885_));
 sky130_fd_sc_hd__nand2_1 _29359_ (.A(_00884_),
    .B(_00885_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand3b_1 _29360_ (.A_N(_00883_),
    .B(_00886_),
    .C(_23213_),
    .Y(_00888_));
 sky130_fd_sc_hd__and2_1 _29361_ (.A(_24453_),
    .B(net316),
    .X(_00889_));
 sky130_fd_sc_hd__o21ai_1 _29362_ (.A1(_00883_),
    .A2(_00889_),
    .B1(_23207_),
    .Y(_00890_));
 sky130_fd_sc_hd__o21ai_1 _29363_ (.A1(_21262_),
    .A2(_24454_),
    .B1(_24455_),
    .Y(_00891_));
 sky130_fd_sc_hd__a21oi_1 _29364_ (.A1(_00888_),
    .A2(_00890_),
    .B1(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__and3_1 _29365_ (.A(_24460_),
    .B(_24456_),
    .C(_24459_),
    .X(_00893_));
 sky130_fd_sc_hd__nand3_1 _29366_ (.A(_00888_),
    .B(_00890_),
    .C(_00891_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand3b_1 _29367_ (.A_N(_00892_),
    .B(_00893_),
    .C(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__and3_1 _29368_ (.A(_00888_),
    .B(_00890_),
    .C(_00891_),
    .X(_00896_));
 sky130_fd_sc_hd__o21ai_1 _29369_ (.A1(_00896_),
    .A2(_00892_),
    .B1(_24463_),
    .Y(_00897_));
 sky130_fd_sc_hd__or2_1 _29370_ (.A(_20307_),
    .B(_06249_),
    .X(_00899_));
 sky130_fd_sc_hd__nand2_1 _29371_ (.A(_06260_),
    .B(_20307_),
    .Y(_00900_));
 sky130_fd_sc_hd__and3_1 _29372_ (.A(_00899_),
    .B(_24445_),
    .C(_00900_),
    .X(_00901_));
 sky130_fd_sc_hd__o2bb2a_1 _29373_ (.A1_N(_00900_),
    .A2_N(_00899_),
    .B1(_00963_),
    .B2(_24447_),
    .X(_00902_));
 sky130_fd_sc_hd__nor2_1 _29374_ (.A(_00901_),
    .B(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__a21o_1 _29375_ (.A1(_00895_),
    .A2(_00897_),
    .B1(_00903_),
    .X(_00904_));
 sky130_fd_sc_hd__nand3_1 _29376_ (.A(_00895_),
    .B(_00897_),
    .C(_00903_),
    .Y(_00905_));
 sky130_fd_sc_hd__o211ai_2 _29377_ (.A1(_24464_),
    .A2(net233),
    .B1(_00904_),
    .C1(_00905_),
    .Y(_00906_));
 sky130_fd_sc_hd__a211o_1 _29378_ (.A1(_00904_),
    .A2(_00905_),
    .B1(_24464_),
    .C1(net233),
    .X(_00907_));
 sky130_fd_sc_hd__nand2_1 _29379_ (.A(_00906_),
    .B(_00907_),
    .Y(_00908_));
 sky130_fd_sc_hd__or2_1 _29380_ (.A(_24449_),
    .B(_00908_),
    .X(_00909_));
 sky130_fd_sc_hd__nand2_1 _29381_ (.A(_24449_),
    .B(_00908_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand2_2 _29382_ (.A(_00909_),
    .B(_00910_),
    .Y(_00911_));
 sky130_fd_sc_hd__xnor2_4 _29383_ (.A(_00882_),
    .B(_00911_),
    .Y(_00912_));
 sky130_fd_sc_hd__o22ai_4 _29384_ (.A1(_23222_),
    .A2(_24473_),
    .B1(_24476_),
    .B2(_24481_),
    .Y(_00913_));
 sky130_fd_sc_hd__xnor2_4 _29385_ (.A(_00912_),
    .B(_00913_),
    .Y(_00914_));
 sky130_fd_sc_hd__clkbuf_2 _29386_ (.A(\delay_line[29][7] ),
    .X(_00915_));
 sky130_fd_sc_hd__and3_1 _29387_ (.A(_24433_),
    .B(_18451_),
    .C(_00915_),
    .X(_00916_));
 sky130_fd_sc_hd__nor2b_1 _29388_ (.A(_20332_),
    .B_N(net321),
    .Y(_00917_));
 sky130_fd_sc_hd__and2b_1 _29389_ (.A_N(net321),
    .B(_20332_),
    .X(_00918_));
 sky130_fd_sc_hd__nor2_1 _29390_ (.A(_00917_),
    .B(_00918_),
    .Y(_00920_));
 sky130_fd_sc_hd__o21a_1 _29391_ (.A1(_24431_),
    .A2(_00916_),
    .B1(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__a311oi_2 _29392_ (.A1(_24433_),
    .A2(_18451_),
    .A3(_00915_),
    .B1(_00920_),
    .C1(_24431_),
    .Y(_00922_));
 sky130_fd_sc_hd__or4_1 _29393_ (.A(_21299_),
    .B(_24431_),
    .C(_24432_),
    .D(_23235_),
    .X(_00923_));
 sky130_fd_sc_hd__o211a_1 _29394_ (.A1(_00921_),
    .A2(_00922_),
    .B1(_24438_),
    .C1(_00923_),
    .X(_00924_));
 sky130_fd_sc_hd__a211oi_1 _29395_ (.A1(_24438_),
    .A2(_00923_),
    .B1(_00921_),
    .C1(_00922_),
    .Y(_00925_));
 sky130_fd_sc_hd__inv_2 _29396_ (.A(_24421_),
    .Y(_00926_));
 sky130_fd_sc_hd__nand2_2 _29397_ (.A(_24415_),
    .B(_24417_),
    .Y(_00927_));
 sky130_fd_sc_hd__o2bb2a_2 _29398_ (.A1_N(_01040_),
    .A2_N(_23257_),
    .B1(_19329_),
    .B2(_24405_),
    .X(_00928_));
 sky130_fd_sc_hd__a211oi_2 _29399_ (.A1(_23250_),
    .A2(_23254_),
    .B1(_24396_),
    .C1(_24397_),
    .Y(_00929_));
 sky130_fd_sc_hd__and4_2 _29400_ (.A(_24404_),
    .B(_24406_),
    .C(_24400_),
    .D(_24401_),
    .X(_00931_));
 sky130_fd_sc_hd__inv_2 _29401_ (.A(\delay_line[30][11] ),
    .Y(_00932_));
 sky130_fd_sc_hd__nor2_1 _29402_ (.A(_19335_),
    .B(_23269_),
    .Y(_00933_));
 sky130_fd_sc_hd__and2_1 _29403_ (.A(_19335_),
    .B(_21307_),
    .X(_00934_));
 sky130_fd_sc_hd__or3_1 _29404_ (.A(_00932_),
    .B(_00933_),
    .C(_00934_),
    .X(_00935_));
 sky130_fd_sc_hd__o21ai_1 _29405_ (.A1(_00933_),
    .A2(_00934_),
    .B1(_00932_),
    .Y(_00936_));
 sky130_fd_sc_hd__and3_1 _29406_ (.A(_00935_),
    .B(_00936_),
    .C(_24396_),
    .X(_00937_));
 sky130_fd_sc_hd__a21oi_2 _29407_ (.A1(_00935_),
    .A2(_00936_),
    .B1(_24396_),
    .Y(_00938_));
 sky130_fd_sc_hd__nor2_1 _29408_ (.A(_00937_),
    .B(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29409_ (.A(_20348_),
    .X(_00940_));
 sky130_fd_sc_hd__o21ai_2 _29410_ (.A1(_00940_),
    .A2(_23268_),
    .B1(_06315_),
    .Y(_00942_));
 sky130_fd_sc_hd__or3_2 _29411_ (.A(_06304_),
    .B(_00940_),
    .C(_23268_),
    .X(_00943_));
 sky130_fd_sc_hd__a2bb2o_1 _29412_ (.A1_N(_20343_),
    .A2_N(_01018_),
    .B1(_00942_),
    .B2(_00943_),
    .X(_00944_));
 sky130_fd_sc_hd__nand3_1 _29413_ (.A(_00943_),
    .B(_00942_),
    .C(_20346_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand3_2 _29414_ (.A(_00939_),
    .B(_00944_),
    .C(_00945_),
    .Y(_00946_));
 sky130_fd_sc_hd__nand2_1 _29415_ (.A(_00945_),
    .B(_00944_),
    .Y(_00947_));
 sky130_fd_sc_hd__o21ai_2 _29416_ (.A1(_00937_),
    .A2(_00938_),
    .B1(_00947_),
    .Y(_00948_));
 sky130_fd_sc_hd__o211ai_4 _29417_ (.A1(_00929_),
    .A2(_00931_),
    .B1(_00946_),
    .C1(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__a221o_1 _29418_ (.A1(_24399_),
    .A2(_24398_),
    .B1(_00946_),
    .B2(_00948_),
    .C1(_00931_),
    .X(_00950_));
 sky130_fd_sc_hd__nand2_2 _29419_ (.A(_00949_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__xor2_4 _29420_ (.A(_00928_),
    .B(_00951_),
    .X(_00953_));
 sky130_fd_sc_hd__xnor2_2 _29421_ (.A(_00927_),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__nand2_1 _29422_ (.A(_24428_),
    .B(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__a21oi_1 _29423_ (.A1(_24422_),
    .A2(_24428_),
    .B1(_00954_),
    .Y(_00956_));
 sky130_fd_sc_hd__and3_1 _29424_ (.A(_24422_),
    .B(_24428_),
    .C(_00954_),
    .X(_00957_));
 sky130_fd_sc_hd__o22a_1 _29425_ (.A1(_24418_),
    .A2(_24419_),
    .B1(_00956_),
    .B2(_00957_),
    .X(_00958_));
 sky130_fd_sc_hd__a21oi_1 _29426_ (.A1(_00926_),
    .A2(_00955_),
    .B1(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__or3b_2 _29427_ (.A(_00924_),
    .B(_00925_),
    .C_N(_00959_),
    .X(_00960_));
 sky130_fd_sc_hd__o21bai_1 _29428_ (.A1(_00924_),
    .A2(_00925_),
    .B1_N(_00959_),
    .Y(_00961_));
 sky130_fd_sc_hd__nand2_2 _29429_ (.A(_00960_),
    .B(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__xnor2_4 _29430_ (.A(_00914_),
    .B(_00962_),
    .Y(_00964_));
 sky130_fd_sc_hd__nor2_1 _29431_ (.A(_23158_),
    .B(net330),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _29432_ (.A(_23158_),
    .B(net330),
    .Y(_00966_));
 sky130_fd_sc_hd__nand3b_2 _29433_ (.A_N(_00965_),
    .B(_24363_),
    .C(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__and2_1 _29434_ (.A(\delay_line[27][9] ),
    .B(\delay_line[27][11] ),
    .X(_00968_));
 sky130_fd_sc_hd__o21ai_2 _29435_ (.A1(_00968_),
    .A2(_00965_),
    .B1(_24361_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand3_1 _29436_ (.A(_24362_),
    .B(_00967_),
    .C(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__clkbuf_2 _29437_ (.A(net330),
    .X(_00971_));
 sky130_fd_sc_hd__nor2_1 _29438_ (.A(_24359_),
    .B(_24363_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand4_1 _29439_ (.A(_20373_),
    .B(_23158_),
    .C(_00971_),
    .D(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__a21oi_1 _29440_ (.A1(_00970_),
    .A2(_00973_),
    .B1(_18499_),
    .Y(_00975_));
 sky130_fd_sc_hd__and3_1 _29441_ (.A(_18498_),
    .B(_00970_),
    .C(_00973_),
    .X(_00976_));
 sky130_fd_sc_hd__o221ai_2 _29442_ (.A1(_23162_),
    .A2(_24366_),
    .B1(_00975_),
    .B2(_00976_),
    .C1(_24370_),
    .Y(_00977_));
 sky130_fd_sc_hd__nor2_1 _29443_ (.A(_00976_),
    .B(_00975_),
    .Y(_00978_));
 sky130_fd_sc_hd__a31o_1 _29444_ (.A1(_24368_),
    .A2(_16119_),
    .A3(_16086_),
    .B1(_24367_),
    .X(_00979_));
 sky130_fd_sc_hd__nand2_1 _29445_ (.A(_00978_),
    .B(_00979_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand3b_1 _29446_ (.A_N(_16108_),
    .B(_00977_),
    .C(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__a21bo_1 _29447_ (.A1(_00977_),
    .A2(_00980_),
    .B1_N(_16097_),
    .X(_00982_));
 sky130_fd_sc_hd__nand2_1 _29448_ (.A(_00981_),
    .B(_00982_),
    .Y(_00983_));
 sky130_fd_sc_hd__and3_1 _29449_ (.A(_24374_),
    .B(_24375_),
    .C(_00983_),
    .X(_00984_));
 sky130_fd_sc_hd__a21o_1 _29450_ (.A1(_24374_),
    .A2(_24375_),
    .B1(_00983_),
    .X(_00986_));
 sky130_fd_sc_hd__inv_2 _29451_ (.A(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__nor4_1 _29452_ (.A(_23165_),
    .B(_00984_),
    .C(_24377_),
    .D(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__o22a_1 _29453_ (.A1(_23165_),
    .A2(_24377_),
    .B1(_00987_),
    .B2(_00984_),
    .X(_00989_));
 sky130_fd_sc_hd__or2_1 _29454_ (.A(_23168_),
    .B(_23167_),
    .X(_00990_));
 sky130_fd_sc_hd__a2bb2oi_1 _29455_ (.A1_N(_24377_),
    .A2_N(_00990_),
    .B1(_24379_),
    .B2(_24382_),
    .Y(_00991_));
 sky130_fd_sc_hd__nor3_1 _29456_ (.A(net135),
    .B(_00989_),
    .C(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__o21a_1 _29457_ (.A1(net135),
    .A2(_00989_),
    .B1(_00991_),
    .X(_00993_));
 sky130_fd_sc_hd__buf_1 _29458_ (.A(\delay_line[26][10] ),
    .X(_00994_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29459_ (.A(_00994_),
    .X(_00995_));
 sky130_fd_sc_hd__o21a_1 _29460_ (.A1(_18486_),
    .A2(_24338_),
    .B1(_01161_),
    .X(_00997_));
 sky130_fd_sc_hd__buf_1 _29461_ (.A(\delay_line[26][6] ),
    .X(_00998_));
 sky130_fd_sc_hd__nor2_1 _29462_ (.A(net338),
    .B(_00998_),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_1 _29463_ (.A(_24338_),
    .B(_00998_),
    .Y(_01000_));
 sky130_fd_sc_hd__nand3b_2 _29464_ (.A_N(_00999_),
    .B(_01000_),
    .C(net339),
    .Y(_01001_));
 sky130_fd_sc_hd__and2_1 _29465_ (.A(net338),
    .B(_00998_),
    .X(_01002_));
 sky130_fd_sc_hd__o21ai_2 _29466_ (.A1(_00999_),
    .A2(_01002_),
    .B1(_06469_),
    .Y(_01003_));
 sky130_fd_sc_hd__o211a_1 _29467_ (.A1(_24340_),
    .A2(_00997_),
    .B1(_01001_),
    .C1(_01003_),
    .X(_01004_));
 sky130_fd_sc_hd__a21o_1 _29468_ (.A1(_19271_),
    .A2(_19264_),
    .B1(_00997_),
    .X(_01005_));
 sky130_fd_sc_hd__a21oi_1 _29469_ (.A1(_01001_),
    .A2(_01003_),
    .B1(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__o21ai_1 _29470_ (.A1(_23132_),
    .A2(_24351_),
    .B1(_24344_),
    .Y(_01008_));
 sky130_fd_sc_hd__or3_1 _29471_ (.A(_01004_),
    .B(_01006_),
    .C(_01008_),
    .X(_01009_));
 sky130_fd_sc_hd__o21ai_1 _29472_ (.A1(_01004_),
    .A2(_01006_),
    .B1(_01008_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand3b_1 _29473_ (.A_N(_00995_),
    .B(_01009_),
    .C(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__a21bo_1 _29474_ (.A1(_01009_),
    .A2(_01010_),
    .B1_N(_00995_),
    .X(_01012_));
 sky130_fd_sc_hd__o41ai_2 _29475_ (.A1(_23134_),
    .A2(_23135_),
    .A3(_24350_),
    .A4(_24351_),
    .B1(_24354_),
    .Y(_01013_));
 sky130_fd_sc_hd__a21o_1 _29476_ (.A1(_01011_),
    .A2(_01012_),
    .B1(_01013_),
    .X(_01014_));
 sky130_fd_sc_hd__nand3_2 _29477_ (.A(_01013_),
    .B(_01011_),
    .C(_01012_),
    .Y(_01015_));
 sky130_fd_sc_hd__a21oi_1 _29478_ (.A1(_24353_),
    .A2(_24354_),
    .B1(_24335_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand3_1 _29479_ (.A(_24335_),
    .B(_24353_),
    .C(_24354_),
    .Y(_01017_));
 sky130_fd_sc_hd__o21ai_2 _29480_ (.A1(_01016_),
    .A2(_23145_),
    .B1(_01017_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand3_1 _29481_ (.A(_01014_),
    .B(_01015_),
    .C(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__a21o_1 _29482_ (.A1(_01014_),
    .A2(_01015_),
    .B1(_01019_),
    .X(_01021_));
 sky130_fd_sc_hd__nand2_1 _29483_ (.A(_01020_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__o21ai_1 _29484_ (.A1(net107),
    .A2(_00993_),
    .B1(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__or3_1 _29485_ (.A(_01022_),
    .B(net107),
    .C(_00993_),
    .X(_01024_));
 sky130_fd_sc_hd__nand2_1 _29486_ (.A(_01023_),
    .B(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__o21ba_1 _29487_ (.A1(_20428_),
    .A2(_24320_),
    .B1_N(_24321_),
    .X(_01026_));
 sky130_fd_sc_hd__and3_1 _29488_ (.A(_24312_),
    .B(_24313_),
    .C(_24315_),
    .X(_01027_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29489_ (.A(_24311_),
    .X(_01028_));
 sky130_fd_sc_hd__and3_1 _29490_ (.A(_01028_),
    .B(_23178_),
    .C(_23177_),
    .X(_01030_));
 sky130_fd_sc_hd__clkbuf_2 _29491_ (.A(\delay_line[28][10] ),
    .X(_01031_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29492_ (.A(net326),
    .X(_01032_));
 sky130_fd_sc_hd__nand3_1 _29493_ (.A(_23179_),
    .B(_01031_),
    .C(net326),
    .Y(_01033_));
 sky130_fd_sc_hd__or3_2 _29494_ (.A(\delay_line[28][11] ),
    .B(_24311_),
    .C(_23179_),
    .X(_01034_));
 sky130_fd_sc_hd__o2111ai_2 _29495_ (.A1(_01031_),
    .A2(_01032_),
    .B1(_01033_),
    .C1(_19304_),
    .D1(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__o21a_1 _29496_ (.A1(_01031_),
    .A2(_01032_),
    .B1(_01033_),
    .X(_01036_));
 sky130_fd_sc_hd__a21o_1 _29497_ (.A1(_01034_),
    .A2(_01036_),
    .B1(_19304_),
    .X(_01037_));
 sky130_fd_sc_hd__o211a_1 _29498_ (.A1(_01027_),
    .A2(_01030_),
    .B1(_01035_),
    .C1(_01037_),
    .X(_01038_));
 sky130_fd_sc_hd__a211oi_1 _29499_ (.A1(_01035_),
    .A2(_01037_),
    .B1(_01027_),
    .C1(_01030_),
    .Y(_01039_));
 sky130_fd_sc_hd__nor3b_2 _29500_ (.A(_01038_),
    .B(_01039_),
    .C_N(_24315_),
    .Y(_01041_));
 sky130_fd_sc_hd__o21ba_1 _29501_ (.A1(_01038_),
    .A2(_01039_),
    .B1_N(_24315_),
    .X(_01042_));
 sky130_fd_sc_hd__nor3_1 _29502_ (.A(_01026_),
    .B(_01041_),
    .C(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__o21a_1 _29503_ (.A1(_01041_),
    .A2(_01042_),
    .B1(_01026_),
    .X(_01044_));
 sky130_fd_sc_hd__nor3_1 _29504_ (.A(_24327_),
    .B(net206),
    .C(_01044_),
    .Y(_01045_));
 sky130_fd_sc_hd__o21a_1 _29505_ (.A1(net206),
    .A2(_01044_),
    .B1(_24327_),
    .X(_01046_));
 sky130_fd_sc_hd__or2_1 _29506_ (.A(_01045_),
    .B(_01046_),
    .X(_01047_));
 sky130_fd_sc_hd__a21oi_1 _29507_ (.A1(_24333_),
    .A2(_24331_),
    .B1(_24329_),
    .Y(_01048_));
 sky130_fd_sc_hd__xnor2_1 _29508_ (.A(_01047_),
    .B(_01048_),
    .Y(_01049_));
 sky130_fd_sc_hd__nand2_1 _29509_ (.A(_01025_),
    .B(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__or2_1 _29510_ (.A(_01025_),
    .B(_01049_),
    .X(_01052_));
 sky130_fd_sc_hd__nand2_2 _29511_ (.A(_01050_),
    .B(_01052_),
    .Y(_01053_));
 sky130_fd_sc_hd__and3_1 _29512_ (.A(_24384_),
    .B(_24387_),
    .C(_01053_),
    .X(_01054_));
 sky130_fd_sc_hd__a21oi_4 _29513_ (.A1(_24384_),
    .A2(_24387_),
    .B1(_01053_),
    .Y(_01055_));
 sky130_fd_sc_hd__nor2_2 _29514_ (.A(_01054_),
    .B(_01055_),
    .Y(_01056_));
 sky130_fd_sc_hd__xnor2_4 _29515_ (.A(_00964_),
    .B(_01056_),
    .Y(_01057_));
 sky130_fd_sc_hd__nor3_1 _29516_ (.A(_24617_),
    .B(_24619_),
    .C(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__o21a_1 _29517_ (.A1(_24617_),
    .A2(_24619_),
    .B1(_01057_),
    .X(_01059_));
 sky130_fd_sc_hd__nor2_1 _29518_ (.A(_01058_),
    .B(_01059_),
    .Y(_01060_));
 sky130_fd_sc_hd__or2_4 _29519_ (.A(_24392_),
    .B(_24486_),
    .X(_01061_));
 sky130_fd_sc_hd__xor2_1 _29520_ (.A(_01060_),
    .B(_01061_),
    .X(_01063_));
 sky130_fd_sc_hd__xnor2_1 _29521_ (.A(_00881_),
    .B(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__xor2_1 _29522_ (.A(_00463_),
    .B(_01064_),
    .X(_01065_));
 sky130_fd_sc_hd__a21oi_2 _29523_ (.A1(_25011_),
    .A2(_25118_),
    .B1(_25010_),
    .Y(_01066_));
 sky130_fd_sc_hd__a21oi_1 _29524_ (.A1(_24489_),
    .A2(_24492_),
    .B1(_24488_),
    .Y(_01067_));
 sky130_fd_sc_hd__nor2_1 _29525_ (.A(_24944_),
    .B(_24945_),
    .Y(_01068_));
 sky130_fd_sc_hd__nor2_1 _29526_ (.A(_24988_),
    .B(_24994_),
    .Y(_01069_));
 sky130_fd_sc_hd__or2b_2 _29527_ (.A(_24483_),
    .B_N(_24441_),
    .X(_01070_));
 sky130_fd_sc_hd__nor2_1 _29528_ (.A(_24872_),
    .B(_24903_),
    .Y(_01071_));
 sky130_fd_sc_hd__buf_1 _29529_ (.A(\delay_line[34][8] ),
    .X(_01072_));
 sky130_fd_sc_hd__or2_1 _29530_ (.A(_20741_),
    .B(_01072_),
    .X(_01074_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29531_ (.A(_20741_),
    .X(_01075_));
 sky130_fd_sc_hd__nand2_1 _29532_ (.A(_01075_),
    .B(_01072_),
    .Y(_01076_));
 sky130_fd_sc_hd__nor2_1 _29533_ (.A(_23312_),
    .B(net306),
    .Y(_01077_));
 sky130_fd_sc_hd__buf_1 _29534_ (.A(_23312_),
    .X(_01078_));
 sky130_fd_sc_hd__buf_1 _29535_ (.A(net306),
    .X(_01079_));
 sky130_fd_sc_hd__nand2_1 _29536_ (.A(_01078_),
    .B(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand3b_1 _29537_ (.A_N(_01077_),
    .B(_24883_),
    .C(_01080_),
    .Y(_01081_));
 sky130_fd_sc_hd__and2_1 _29538_ (.A(_23312_),
    .B(net306),
    .X(_01082_));
 sky130_fd_sc_hd__o21ai_1 _29539_ (.A1(_01082_),
    .A2(_01077_),
    .B1(_24881_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand4_1 _29540_ (.A(_01074_),
    .B(_01076_),
    .C(_01081_),
    .D(_01083_),
    .Y(_01085_));
 sky130_fd_sc_hd__a22o_1 _29541_ (.A1(_01074_),
    .A2(_01076_),
    .B1(_01081_),
    .B2(_01083_),
    .X(_01086_));
 sky130_fd_sc_hd__nand2_1 _29542_ (.A(_01085_),
    .B(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__a21boi_2 _29543_ (.A1(_24884_),
    .A2(_24888_),
    .B1_N(_24882_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand2_1 _29544_ (.A(_01087_),
    .B(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand3b_1 _29545_ (.A_N(_01088_),
    .B(_01085_),
    .C(_01086_),
    .Y(_01090_));
 sky130_fd_sc_hd__a21boi_1 _29546_ (.A1(_24874_),
    .A2(_01075_),
    .B1_N(_17812_),
    .Y(_01091_));
 sky130_fd_sc_hd__and3b_1 _29547_ (.A_N(_17812_),
    .B(_24874_),
    .C(_01075_),
    .X(_01092_));
 sky130_fd_sc_hd__nor2_1 _29548_ (.A(_01091_),
    .B(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__a21oi_1 _29549_ (.A1(_01089_),
    .A2(_01090_),
    .B1(_01093_),
    .Y(_01094_));
 sky130_fd_sc_hd__and3_1 _29550_ (.A(_01089_),
    .B(_01090_),
    .C(_01093_),
    .X(_01096_));
 sky130_fd_sc_hd__o211a_1 _29551_ (.A1(_01094_),
    .A2(_01096_),
    .B1(_24892_),
    .C1(_24895_),
    .X(_01097_));
 sky130_fd_sc_hd__a211oi_2 _29552_ (.A1(_24892_),
    .A2(_24895_),
    .B1(_01094_),
    .C1(_01096_),
    .Y(_01098_));
 sky130_fd_sc_hd__nor2_1 _29553_ (.A(_01097_),
    .B(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__xnor2_1 _29554_ (.A(_24878_),
    .B(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hd__o31a_1 _29555_ (.A1(_02260_),
    .A2(_21097_),
    .A3(_24898_),
    .B1(_24899_),
    .X(_01101_));
 sky130_fd_sc_hd__nand2_1 _29556_ (.A(_01100_),
    .B(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__a21o_1 _29557_ (.A1(_24899_),
    .A2(_24900_),
    .B1(_01100_),
    .X(_01103_));
 sky130_fd_sc_hd__and2_1 _29558_ (.A(_01102_),
    .B(_01103_),
    .X(_01104_));
 sky130_fd_sc_hd__a211o_1 _29559_ (.A1(_24907_),
    .A2(_24904_),
    .B1(_01071_),
    .C1(_01104_),
    .X(_01105_));
 sky130_fd_sc_hd__a21o_1 _29560_ (.A1(_24904_),
    .A2(_24907_),
    .B1(_01071_),
    .X(_01107_));
 sky130_fd_sc_hd__nand2_1 _29561_ (.A(_01107_),
    .B(_01104_),
    .Y(_01108_));
 sky130_fd_sc_hd__and2_1 _29562_ (.A(_01105_),
    .B(_01108_),
    .X(_01109_));
 sky130_fd_sc_hd__a21bo_1 _29563_ (.A1(_24982_),
    .A2(_23387_),
    .B1_N(_24981_),
    .X(_01110_));
 sky130_fd_sc_hd__buf_1 _29564_ (.A(\delay_line[32][11] ),
    .X(_01111_));
 sky130_fd_sc_hd__nor2_1 _29565_ (.A(_24956_),
    .B(_01111_),
    .Y(_01112_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29566_ (.A(\delay_line[32][11] ),
    .X(_01113_));
 sky130_fd_sc_hd__nand2_1 _29567_ (.A(_24956_),
    .B(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__clkbuf_2 _29568_ (.A(_23389_),
    .X(_01115_));
 sky130_fd_sc_hd__nand3b_1 _29569_ (.A_N(_01112_),
    .B(_01114_),
    .C(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__and2_1 _29570_ (.A(_24956_),
    .B(_01111_),
    .X(_01118_));
 sky130_fd_sc_hd__inv_2 _29571_ (.A(_24954_),
    .Y(_01119_));
 sky130_fd_sc_hd__o21ai_1 _29572_ (.A1(_01112_),
    .A2(_01118_),
    .B1(_01119_),
    .Y(_01120_));
 sky130_fd_sc_hd__buf_1 _29573_ (.A(_21113_),
    .X(_01121_));
 sky130_fd_sc_hd__o21ai_1 _29574_ (.A1(_01121_),
    .A2(_24955_),
    .B1(_24957_),
    .Y(_01122_));
 sky130_fd_sc_hd__nand3_1 _29575_ (.A(_01116_),
    .B(_01120_),
    .C(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__a21o_1 _29576_ (.A1(_01116_),
    .A2(_01120_),
    .B1(_01122_),
    .X(_01124_));
 sky130_fd_sc_hd__a21o_1 _29577_ (.A1(_01123_),
    .A2(_01124_),
    .B1(_01121_),
    .X(_01125_));
 sky130_fd_sc_hd__nand3_1 _29578_ (.A(_01121_),
    .B(_01123_),
    .C(_01124_),
    .Y(_01126_));
 sky130_fd_sc_hd__a21oi_1 _29579_ (.A1(_24966_),
    .A2(_21126_),
    .B1(_24965_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand3_1 _29580_ (.A(_01125_),
    .B(_01126_),
    .C(_01127_),
    .Y(_01129_));
 sky130_fd_sc_hd__a21o_1 _29581_ (.A1(_01125_),
    .A2(_01126_),
    .B1(_01127_),
    .X(_01130_));
 sky130_fd_sc_hd__and2_1 _29582_ (.A(_05249_),
    .B(_18667_),
    .X(_01131_));
 sky130_fd_sc_hd__buf_1 _29583_ (.A(_18667_),
    .X(_01132_));
 sky130_fd_sc_hd__nor2_1 _29584_ (.A(_01132_),
    .B(_05260_),
    .Y(_01133_));
 sky130_fd_sc_hd__nor2_1 _29585_ (.A(_01131_),
    .B(_01133_),
    .Y(_01134_));
 sky130_fd_sc_hd__xnor2_1 _29586_ (.A(_24949_),
    .B(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand3_2 _29587_ (.A(_01129_),
    .B(_01130_),
    .C(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__a21o_1 _29588_ (.A1(_01129_),
    .A2(_01130_),
    .B1(_01135_),
    .X(_01137_));
 sky130_fd_sc_hd__a21o_1 _29589_ (.A1(_24977_),
    .A2(_24979_),
    .B1(_24975_),
    .X(_01138_));
 sky130_fd_sc_hd__a21oi_1 _29590_ (.A1(_01136_),
    .A2(_01137_),
    .B1(_01138_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand3_1 _29591_ (.A(_01138_),
    .B(_01136_),
    .C(_01137_),
    .Y(_01141_));
 sky130_fd_sc_hd__nand3b_2 _29592_ (.A_N(_01140_),
    .B(_01141_),
    .C(_24951_),
    .Y(_01142_));
 sky130_fd_sc_hd__and3_1 _29593_ (.A(_01138_),
    .B(_01136_),
    .C(_01137_),
    .X(_01143_));
 sky130_fd_sc_hd__o21bai_1 _29594_ (.A1(_01140_),
    .A2(_01143_),
    .B1_N(_24951_),
    .Y(_01144_));
 sky130_fd_sc_hd__and3_1 _29595_ (.A(_01110_),
    .B(_01142_),
    .C(_01144_),
    .X(_01145_));
 sky130_fd_sc_hd__clkbuf_2 _29596_ (.A(_01145_),
    .X(_01146_));
 sky130_fd_sc_hd__a21oi_1 _29597_ (.A1(_01142_),
    .A2(_01144_),
    .B1(_01110_),
    .Y(_01147_));
 sky130_fd_sc_hd__inv_2 _29598_ (.A(_24986_),
    .Y(_01148_));
 sky130_fd_sc_hd__or4bb_1 _29599_ (.A(_01146_),
    .B(_01147_),
    .C_N(_24947_),
    .D_N(_01148_),
    .X(_01149_));
 sky130_fd_sc_hd__buf_1 _29600_ (.A(_01148_),
    .X(_01151_));
 sky130_fd_sc_hd__a2bb2o_1 _29601_ (.A1_N(_01146_),
    .A2_N(_01147_),
    .B1(_24947_),
    .B2(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__nand2_1 _29602_ (.A(_01149_),
    .B(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__and4_1 _29603_ (.A(_23407_),
    .B(_21140_),
    .C(_21139_),
    .D(_21138_),
    .X(_01154_));
 sky130_fd_sc_hd__a22oi_2 _29604_ (.A1(_01154_),
    .A2(_01151_),
    .B1(_24993_),
    .B2(_24987_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _29605_ (.A(_01153_),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hd__inv_2 _29606_ (.A(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__nor2_1 _29607_ (.A(_23376_),
    .B(_24942_),
    .Y(_01158_));
 sky130_fd_sc_hd__a2111oi_4 _29608_ (.A1(_17824_),
    .A2(_24918_),
    .B1(_23367_),
    .C1(_00568_),
    .D1(_24916_),
    .Y(_01159_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29609_ (.A(_24913_),
    .X(_01160_));
 sky130_fd_sc_hd__and3_1 _29610_ (.A(_02172_),
    .B(_17824_),
    .C(_01160_),
    .X(_01162_));
 sky130_fd_sc_hd__inv_2 _29611_ (.A(\delay_line[33][11] ),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _29612_ (.A(_20671_),
    .B(_19576_),
    .Y(_01164_));
 sky130_fd_sc_hd__nand2_1 _29613_ (.A(_19573_),
    .B(_20666_),
    .Y(_01165_));
 sky130_fd_sc_hd__nand3_1 _29614_ (.A(_01163_),
    .B(_01164_),
    .C(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__a21o_1 _29615_ (.A1(_01164_),
    .A2(_01165_),
    .B1(_01163_),
    .X(_01167_));
 sky130_fd_sc_hd__a21oi_1 _29616_ (.A1(_01166_),
    .A2(_01167_),
    .B1(_24926_),
    .Y(_01168_));
 sky130_fd_sc_hd__a21oi_1 _29617_ (.A1(_19574_),
    .A2(_23352_),
    .B1(_23366_),
    .Y(_01169_));
 sky130_fd_sc_hd__or2b_1 _29618_ (.A(_02150_),
    .B_N(\delay_line[33][4] ),
    .X(_01170_));
 sky130_fd_sc_hd__a31o_1 _29619_ (.A1(_23366_),
    .A2(_24913_),
    .A3(_19574_),
    .B1(_01170_),
    .X(_01171_));
 sky130_fd_sc_hd__and3_1 _29620_ (.A(_23366_),
    .B(_19574_),
    .C(_23352_),
    .X(_01173_));
 sky130_fd_sc_hd__o21ai_1 _29621_ (.A1(_01173_),
    .A2(_01169_),
    .B1(_01170_),
    .Y(_01174_));
 sky130_fd_sc_hd__o21ai_1 _29622_ (.A1(_01169_),
    .A2(_01171_),
    .B1(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__and3_1 _29623_ (.A(_01167_),
    .B(_24926_),
    .C(_01166_),
    .X(_01176_));
 sky130_fd_sc_hd__nor3_1 _29624_ (.A(_01168_),
    .B(_01175_),
    .C(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__o21a_1 _29625_ (.A1(_01176_),
    .A2(_01168_),
    .B1(_01175_),
    .X(_01178_));
 sky130_fd_sc_hd__o221ai_4 _29626_ (.A1(_24934_),
    .A2(_24933_),
    .B1(net232),
    .B2(_01178_),
    .C1(_24928_),
    .Y(_01179_));
 sky130_fd_sc_hd__nor2_1 _29627_ (.A(net232),
    .B(_01178_),
    .Y(_01180_));
 sky130_fd_sc_hd__a31o_1 _29628_ (.A1(_24917_),
    .A2(_24920_),
    .A3(_24929_),
    .B1(_24932_),
    .X(_01181_));
 sky130_fd_sc_hd__nand2_1 _29629_ (.A(_01180_),
    .B(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__o211a_1 _29630_ (.A1(_01159_),
    .A2(_01162_),
    .B1(_01179_),
    .C1(_01182_),
    .X(_01184_));
 sky130_fd_sc_hd__clkbuf_2 _29631_ (.A(_01182_),
    .X(_01185_));
 sky130_fd_sc_hd__a31o_1 _29632_ (.A1(_02172_),
    .A2(_17824_),
    .A3(_01160_),
    .B1(_01159_),
    .X(_01186_));
 sky130_fd_sc_hd__a21oi_1 _29633_ (.A1(_01179_),
    .A2(_01185_),
    .B1(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _29634_ (.A(_00579_),
    .B(_02183_),
    .Y(_01188_));
 sky130_fd_sc_hd__a21oi_1 _29635_ (.A1(_24931_),
    .A2(_24935_),
    .B1(_24936_),
    .Y(_01189_));
 sky130_fd_sc_hd__o31ai_2 _29636_ (.A1(_23367_),
    .A2(_01188_),
    .A3(_01189_),
    .B1(_24938_),
    .Y(_01190_));
 sky130_fd_sc_hd__o21bai_2 _29637_ (.A1(_01184_),
    .A2(_01187_),
    .B1_N(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__o211ai_4 _29638_ (.A1(_01159_),
    .A2(_01162_),
    .B1(_01179_),
    .C1(_01185_),
    .Y(_01192_));
 sky130_fd_sc_hd__a21o_1 _29639_ (.A1(_01179_),
    .A2(_01185_),
    .B1(_01186_),
    .X(_01193_));
 sky130_fd_sc_hd__nand3_2 _29640_ (.A(_01192_),
    .B(_01193_),
    .C(_01190_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand3_1 _29641_ (.A(_01158_),
    .B(_01191_),
    .C(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__a2bb2o_1 _29642_ (.A1_N(_23376_),
    .A2_N(_24942_),
    .B1(_01191_),
    .B2(_01195_),
    .X(_01197_));
 sky130_fd_sc_hd__and2_1 _29643_ (.A(_01196_),
    .B(_01197_),
    .X(_01198_));
 sky130_fd_sc_hd__o22ai_4 _29644_ (.A1(_24911_),
    .A2(_24942_),
    .B1(_24943_),
    .B2(_24910_),
    .Y(_01199_));
 sky130_fd_sc_hd__xor2_1 _29645_ (.A(_01198_),
    .B(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__nand2_1 _29646_ (.A(_01155_),
    .B(_01153_),
    .Y(_01201_));
 sky130_fd_sc_hd__and3_1 _29647_ (.A(_01157_),
    .B(_01200_),
    .C(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__a21oi_1 _29648_ (.A1(_01201_),
    .A2(_01157_),
    .B1(_01200_),
    .Y(_01203_));
 sky130_fd_sc_hd__nor2_1 _29649_ (.A(_01202_),
    .B(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__xnor2_1 _29650_ (.A(_01109_),
    .B(_01204_),
    .Y(_01206_));
 sky130_fd_sc_hd__and3_1 _29651_ (.A(_24440_),
    .B(_01070_),
    .C(_01206_),
    .X(_01207_));
 sky130_fd_sc_hd__a21oi_1 _29652_ (.A1(_24440_),
    .A2(_01070_),
    .B1(_01206_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _29653_ (.A(_01207_),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__a211oi_1 _29654_ (.A1(_01068_),
    .A2(_01069_),
    .B1(_24999_),
    .C1(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__o21a_1 _29655_ (.A1(_24997_),
    .A2(_24999_),
    .B1(_01209_),
    .X(_01211_));
 sky130_fd_sc_hd__a211o_1 _29656_ (.A1(_25003_),
    .A2(_25005_),
    .B1(_01210_),
    .C1(_01211_),
    .X(_01212_));
 sky130_fd_sc_hd__o211ai_2 _29657_ (.A1(_01210_),
    .A2(_01211_),
    .B1(_25003_),
    .C1(_25005_),
    .Y(_01213_));
 sky130_fd_sc_hd__nand2_1 _29658_ (.A(_01212_),
    .B(_01213_),
    .Y(_01214_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29659_ (.A(\delay_line[38][8] ),
    .X(_01215_));
 sky130_fd_sc_hd__nand4_2 _29660_ (.A(_21003_),
    .B(_01215_),
    .C(_23433_),
    .D(_25034_),
    .Y(_01217_));
 sky130_fd_sc_hd__and3_1 _29661_ (.A(_23429_),
    .B(net286),
    .C(_25033_),
    .X(_01218_));
 sky130_fd_sc_hd__nor2_1 _29662_ (.A(_01215_),
    .B(\delay_line[38][11] ),
    .Y(_01219_));
 sky130_fd_sc_hd__and2_1 _29663_ (.A(_01215_),
    .B(\delay_line[38][11] ),
    .X(_01220_));
 sky130_fd_sc_hd__nor2_1 _29664_ (.A(_01219_),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__o21a_1 _29665_ (.A1(_25032_),
    .A2(_01218_),
    .B1(_01221_),
    .X(_01222_));
 sky130_fd_sc_hd__clkbuf_2 _29666_ (.A(\delay_line[38][9] ),
    .X(_01223_));
 sky130_fd_sc_hd__clkbuf_2 _29667_ (.A(_01221_),
    .X(_01224_));
 sky130_fd_sc_hd__a311oi_4 _29668_ (.A1(_23429_),
    .A2(_01223_),
    .A3(_25034_),
    .B1(_01224_),
    .C1(_25032_),
    .Y(_01225_));
 sky130_fd_sc_hd__a211oi_2 _29669_ (.A1(_25041_),
    .A2(_01217_),
    .B1(_01222_),
    .C1(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__inv_2 _29670_ (.A(_01226_),
    .Y(_01228_));
 sky130_fd_sc_hd__o211ai_2 _29671_ (.A1(_01225_),
    .A2(_01222_),
    .B1(_01217_),
    .C1(_25041_),
    .Y(_01229_));
 sky130_fd_sc_hd__o21ba_1 _29672_ (.A1(_23452_),
    .A2(_23453_),
    .B1_N(_25023_),
    .X(_01230_));
 sky130_fd_sc_hd__buf_1 _29673_ (.A(\delay_line[39][10] ),
    .X(_01231_));
 sky130_fd_sc_hd__nand2_1 _29674_ (.A(_23443_),
    .B(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__buf_1 _29675_ (.A(\delay_line[39][11] ),
    .X(_01233_));
 sky130_fd_sc_hd__nor2_1 _29676_ (.A(_01231_),
    .B(_01233_),
    .Y(_01234_));
 sky130_fd_sc_hd__and2_1 _29677_ (.A(_01231_),
    .B(\delay_line[39][11] ),
    .X(_01235_));
 sky130_fd_sc_hd__or3_1 _29678_ (.A(_23446_),
    .B(_01234_),
    .C(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__o21ai_1 _29679_ (.A1(_01234_),
    .A2(_01235_),
    .B1(_23446_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_2 _29680_ (.A(_01236_),
    .B(_01237_),
    .Y(_01239_));
 sky130_fd_sc_hd__a21oi_2 _29681_ (.A1(_01232_),
    .A2(_25015_),
    .B1(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__a311oi_4 _29682_ (.A1(_25013_),
    .A2(_01232_),
    .A3(_01239_),
    .B1(_23445_),
    .C1(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__and3_1 _29683_ (.A(_01232_),
    .B(_25015_),
    .C(_01239_),
    .X(_01242_));
 sky130_fd_sc_hd__o21a_1 _29684_ (.A1(_01240_),
    .A2(_01242_),
    .B1(_23445_),
    .X(_01243_));
 sky130_fd_sc_hd__nor2_1 _29685_ (.A(_01241_),
    .B(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__or2_1 _29686_ (.A(_25019_),
    .B(_01244_),
    .X(_01245_));
 sky130_fd_sc_hd__o21a_1 _29687_ (.A1(_25019_),
    .A2(_25020_),
    .B1(_01244_),
    .X(_01246_));
 sky130_fd_sc_hd__o21ba_1 _29688_ (.A1(_25020_),
    .A2(_01245_),
    .B1_N(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__nor3_1 _29689_ (.A(_01230_),
    .B(_25026_),
    .C(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__o21a_1 _29690_ (.A1(_01230_),
    .A2(_25026_),
    .B1(_01247_),
    .X(_01250_));
 sky130_fd_sc_hd__nor2_1 _29691_ (.A(_01248_),
    .B(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__a21o_1 _29692_ (.A1(_01228_),
    .A2(_01229_),
    .B1(_01251_),
    .X(_01252_));
 sky130_fd_sc_hd__nand3_1 _29693_ (.A(_01251_),
    .B(_01229_),
    .C(_01228_),
    .Y(_01253_));
 sky130_fd_sc_hd__buf_1 _29694_ (.A(\delay_line[40][10] ),
    .X(_01254_));
 sky130_fd_sc_hd__a21oi_1 _29695_ (.A1(_25045_),
    .A2(_01254_),
    .B1(\delay_line[40][11] ),
    .Y(_01255_));
 sky130_fd_sc_hd__and3_1 _29696_ (.A(_25045_),
    .B(\delay_line[40][10] ),
    .C(\delay_line[40][11] ),
    .X(_01256_));
 sky130_fd_sc_hd__nor3_2 _29697_ (.A(_21017_),
    .B(_01255_),
    .C(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__o21a_1 _29698_ (.A1(_01255_),
    .A2(_01256_),
    .B1(_21017_),
    .X(_01258_));
 sky130_fd_sc_hd__o211a_1 _29699_ (.A1(_01257_),
    .A2(_01258_),
    .B1(_25047_),
    .C1(_25050_),
    .X(_01259_));
 sky130_fd_sc_hd__a211oi_2 _29700_ (.A1(_25047_),
    .A2(_25050_),
    .B1(_01257_),
    .C1(_01258_),
    .Y(_01261_));
 sky130_fd_sc_hd__o21bai_1 _29701_ (.A1(_25054_),
    .A2(_25056_),
    .B1_N(_25053_),
    .Y(_01262_));
 sky130_fd_sc_hd__or3_1 _29702_ (.A(_01259_),
    .B(_01261_),
    .C(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__o21ai_1 _29703_ (.A1(_01259_),
    .A2(_01261_),
    .B1(_01262_),
    .Y(_01264_));
 sky130_fd_sc_hd__nand2_1 _29704_ (.A(_01263_),
    .B(_01264_),
    .Y(_01265_));
 sky130_fd_sc_hd__a21oi_2 _29705_ (.A1(_01252_),
    .A2(_01253_),
    .B1(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__and3_1 _29706_ (.A(_01252_),
    .B(_01253_),
    .C(_01265_),
    .X(_01267_));
 sky130_fd_sc_hd__or2_2 _29707_ (.A(_01266_),
    .B(_01267_),
    .X(_01268_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29708_ (.A(\delay_line[37][10] ),
    .X(_01269_));
 sky130_fd_sc_hd__a22oi_1 _29709_ (.A1(_01269_),
    .A2(net279),
    .B1(_25074_),
    .B2(_25075_),
    .Y(_01270_));
 sky130_fd_sc_hd__xnor2_1 _29710_ (.A(_23521_),
    .B(\delay_line[37][11] ),
    .Y(_01272_));
 sky130_fd_sc_hd__a21bo_1 _29711_ (.A1(_25068_),
    .A2(_25067_),
    .B1_N(_25066_),
    .X(_01273_));
 sky130_fd_sc_hd__xor2_1 _29712_ (.A(_01272_),
    .B(_01273_),
    .X(_01274_));
 sky130_fd_sc_hd__and2b_1 _29713_ (.A_N(_01270_),
    .B(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__a221oi_1 _29714_ (.A1(_01269_),
    .A2(net279),
    .B1(_25074_),
    .B2(_25075_),
    .C1(_01274_),
    .Y(_01276_));
 sky130_fd_sc_hd__or2_1 _29715_ (.A(_01275_),
    .B(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__or2b_1 _29716_ (.A(_25077_),
    .B_N(\delay_line[36][8] ),
    .X(_01278_));
 sky130_fd_sc_hd__or2b_1 _29717_ (.A(\delay_line[36][8] ),
    .B_N(_25077_),
    .X(_01279_));
 sky130_fd_sc_hd__and3b_1 _29718_ (.A_N(_21046_),
    .B(\delay_line[36][6] ),
    .C(_25081_),
    .X(_01280_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29719_ (.A(_25079_),
    .X(_01281_));
 sky130_fd_sc_hd__o2bb2a_1 _29720_ (.A1_N(_01278_),
    .A2_N(_01279_),
    .B1(_01280_),
    .B2(_01281_),
    .X(_01283_));
 sky130_fd_sc_hd__a21oi_1 _29721_ (.A1(_23484_),
    .A2(_25081_),
    .B1(_01281_),
    .Y(_01284_));
 sky130_fd_sc_hd__and3_1 _29722_ (.A(_01284_),
    .B(_01279_),
    .C(_01278_),
    .X(_01285_));
 sky130_fd_sc_hd__and3_1 _29723_ (.A(net297),
    .B(_21048_),
    .C(_23486_),
    .X(_01286_));
 sky130_fd_sc_hd__or4_1 _29724_ (.A(_25086_),
    .B(_01283_),
    .C(_01285_),
    .D(_01286_),
    .X(_01287_));
 sky130_fd_sc_hd__o22ai_4 _29725_ (.A1(_01283_),
    .A2(_01285_),
    .B1(_01286_),
    .B2(_25086_),
    .Y(_01288_));
 sky130_fd_sc_hd__nor3_1 _29726_ (.A(_19697_),
    .B(_25100_),
    .C(_25102_),
    .Y(_01289_));
 sky130_fd_sc_hd__clkbuf_2 _29727_ (.A(_25091_),
    .X(_01290_));
 sky130_fd_sc_hd__nor2_1 _29728_ (.A(_25091_),
    .B(\delay_line[35][11] ),
    .Y(_01291_));
 sky130_fd_sc_hd__and2_1 _29729_ (.A(\delay_line[35][10] ),
    .B(\delay_line[35][11] ),
    .X(_01292_));
 sky130_fd_sc_hd__or3b_1 _29730_ (.A(_01291_),
    .B(_01292_),
    .C_N(_23496_),
    .X(_01294_));
 sky130_fd_sc_hd__o21bai_2 _29731_ (.A1(_01291_),
    .A2(_01292_),
    .B1_N(_23496_),
    .Y(_01295_));
 sky130_fd_sc_hd__nor3b_1 _29732_ (.A(_25092_),
    .B(_25093_),
    .C_N(_23503_),
    .Y(_01296_));
 sky130_fd_sc_hd__a221oi_1 _29733_ (.A1(_25098_),
    .A2(_01290_),
    .B1(_01294_),
    .B2(_01295_),
    .C1(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__o211ai_2 _29734_ (.A1(_25093_),
    .A2(net278),
    .B1(_01294_),
    .C1(_01295_),
    .Y(_01298_));
 sky130_fd_sc_hd__and3b_1 _29735_ (.A_N(_01297_),
    .B(_25097_),
    .C(_01298_),
    .X(_01299_));
 sky130_fd_sc_hd__o211a_1 _29736_ (.A1(_25093_),
    .A2(net278),
    .B1(_01294_),
    .C1(_01295_),
    .X(_01300_));
 sky130_fd_sc_hd__o21bai_1 _29737_ (.A1(_01300_),
    .A2(_01297_),
    .B1_N(_25097_),
    .Y(_01301_));
 sky130_fd_sc_hd__or2b_1 _29738_ (.A(_01299_),
    .B_N(_01301_),
    .X(_01302_));
 sky130_fd_sc_hd__xor2_1 _29739_ (.A(_20833_),
    .B(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__o21a_1 _29740_ (.A1(_25100_),
    .A2(_01289_),
    .B1(_01303_),
    .X(_01305_));
 sky130_fd_sc_hd__a211oi_1 _29741_ (.A1(_18549_),
    .A2(_25101_),
    .B1(_01303_),
    .C1(_25100_),
    .Y(_01306_));
 sky130_fd_sc_hd__or2_1 _29742_ (.A(_01305_),
    .B(_01306_),
    .X(_01307_));
 sky130_fd_sc_hd__inv_2 _29743_ (.A(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__o21ai_2 _29744_ (.A1(_25109_),
    .A2(_25110_),
    .B1(_25105_),
    .Y(_01309_));
 sky130_fd_sc_hd__xor2_1 _29745_ (.A(_01308_),
    .B(_01309_),
    .X(_01310_));
 sky130_fd_sc_hd__a21oi_1 _29746_ (.A1(_01287_),
    .A2(_01288_),
    .B1(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__and3_1 _29747_ (.A(_01310_),
    .B(_01288_),
    .C(_01287_),
    .X(_01312_));
 sky130_fd_sc_hd__or2_1 _29748_ (.A(_01311_),
    .B(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__or2_1 _29749_ (.A(_01277_),
    .B(_01313_),
    .X(_01314_));
 sky130_fd_sc_hd__nand2_1 _29750_ (.A(_01277_),
    .B(_01313_),
    .Y(_01316_));
 sky130_fd_sc_hd__a22oi_1 _29751_ (.A1(_25087_),
    .A2(_25088_),
    .B1(_25108_),
    .B2(_25111_),
    .Y(_01317_));
 sky130_fd_sc_hd__o21ai_1 _29752_ (.A1(_01317_),
    .A2(_25076_),
    .B1(_25112_),
    .Y(_01318_));
 sky130_fd_sc_hd__a21oi_1 _29753_ (.A1(_01314_),
    .A2(_01316_),
    .B1(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hd__nand3_1 _29754_ (.A(_01318_),
    .B(_01314_),
    .C(_01316_),
    .Y(_01320_));
 sky130_fd_sc_hd__and2b_1 _29755_ (.A_N(_01319_),
    .B(_01320_),
    .X(_01321_));
 sky130_fd_sc_hd__xnor2_4 _29756_ (.A(_01268_),
    .B(_01321_),
    .Y(_01322_));
 sky130_fd_sc_hd__xor2_1 _29757_ (.A(_01214_),
    .B(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__or2_2 _29758_ (.A(_01067_),
    .B(_01323_),
    .X(_01324_));
 sky130_fd_sc_hd__nand2_1 _29759_ (.A(_01323_),
    .B(_01067_),
    .Y(_01325_));
 sky130_fd_sc_hd__nand2_1 _29760_ (.A(_01324_),
    .B(_01325_),
    .Y(_01327_));
 sky130_fd_sc_hd__or2_1 _29761_ (.A(_01066_),
    .B(_01327_),
    .X(_01328_));
 sky130_fd_sc_hd__nand2_1 _29762_ (.A(_01327_),
    .B(_01066_),
    .Y(_01329_));
 sky130_fd_sc_hd__and2_1 _29763_ (.A(_01328_),
    .B(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__xor2_1 _29764_ (.A(_01065_),
    .B(_01330_),
    .X(_01331_));
 sky130_fd_sc_hd__a21oi_2 _29765_ (.A1(_24865_),
    .A2(_25126_),
    .B1(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__and3_1 _29766_ (.A(_24865_),
    .B(_25126_),
    .C(_01331_),
    .X(_01333_));
 sky130_fd_sc_hd__nor2_1 _29767_ (.A(_01332_),
    .B(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__nand3_1 _29768_ (.A(_00460_),
    .B(_00462_),
    .C(_01334_),
    .Y(_01335_));
 sky130_fd_sc_hd__a21boi_1 _29769_ (.A1(_00453_),
    .A2(_00456_),
    .B1_N(_00459_),
    .Y(_01336_));
 sky130_fd_sc_hd__o211a_1 _29770_ (.A1(_25207_),
    .A2(_00461_),
    .B1(_00453_),
    .C1(_00456_),
    .X(_01338_));
 sky130_fd_sc_hd__o22ai_2 _29771_ (.A1(_01332_),
    .A2(_01333_),
    .B1(_01336_),
    .B2(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__nand3_1 _29772_ (.A(_25286_),
    .B(_01335_),
    .C(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29773_ (.A(_01340_),
    .X(_01341_));
 sky130_fd_sc_hd__nand2_1 _29774_ (.A(_01335_),
    .B(_01339_),
    .Y(_01342_));
 sky130_fd_sc_hd__a2bb2oi_1 _29775_ (.A1_N(_25129_),
    .A2_N(_24309_),
    .B1(_24307_),
    .B2(_25141_),
    .Y(_01343_));
 sky130_fd_sc_hd__nand2_1 _29776_ (.A(_01342_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__nand3_1 _29777_ (.A(_25285_),
    .B(_01341_),
    .C(_01344_),
    .Y(_01345_));
 sky130_fd_sc_hd__a21o_1 _29778_ (.A1(_01341_),
    .A2(_01344_),
    .B1(_25285_),
    .X(_01346_));
 sky130_fd_sc_hd__nand3_2 _29779_ (.A(_25206_),
    .B(_01345_),
    .C(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__o22ai_4 _29780_ (.A1(_25131_),
    .A2(_25135_),
    .B1(_25154_),
    .B2(_25148_),
    .Y(_01349_));
 sky130_fd_sc_hd__a22o_1 _29781_ (.A1(_25283_),
    .A2(_25284_),
    .B1(_01340_),
    .B2(_01344_),
    .X(_01350_));
 sky130_fd_sc_hd__nand4_2 _29782_ (.A(_25283_),
    .B(_25284_),
    .C(_01341_),
    .D(_01344_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand3_1 _29783_ (.A(_01349_),
    .B(_01350_),
    .C(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__o2111ai_4 _29784_ (.A1(_22205_),
    .A2(_20967_),
    .B1(_25160_),
    .C1(_25165_),
    .D1(_25166_),
    .Y(_01353_));
 sky130_fd_sc_hd__o211a_1 _29785_ (.A1(_20965_),
    .A2(_20946_),
    .B1(_25238_),
    .C1(_25159_),
    .X(_01354_));
 sky130_fd_sc_hd__o21bai_2 _29786_ (.A1(_04898_),
    .A2(_04909_),
    .B1_N(_19811_),
    .Y(_01355_));
 sky130_fd_sc_hd__or3b_2 _29787_ (.A(_04898_),
    .B(_04909_),
    .C_N(_19811_),
    .X(_01356_));
 sky130_fd_sc_hd__a21o_1 _29788_ (.A1(_04953_),
    .A2(_04931_),
    .B1(_25164_),
    .X(_01357_));
 sky130_fd_sc_hd__a21oi_1 _29789_ (.A1(_01355_),
    .A2(_01356_),
    .B1(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__and3_1 _29790_ (.A(_01357_),
    .B(_01355_),
    .C(_01356_),
    .X(_01360_));
 sky130_fd_sc_hd__nor2_1 _29791_ (.A(_01358_),
    .B(_01360_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2_1 _29792_ (.A(_01354_),
    .B(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__o211a_2 _29793_ (.A1(_20965_),
    .A2(_20946_),
    .B1(_23593_),
    .C1(_01361_),
    .X(_01363_));
 sky130_fd_sc_hd__nor3_2 _29794_ (.A(_01362_),
    .B(_25165_),
    .C(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__nand2_1 _29795_ (.A(_04931_),
    .B(_22177_),
    .Y(_01365_));
 sky130_fd_sc_hd__o32a_1 _29796_ (.A1(_01365_),
    .A2(_25164_),
    .A3(_25163_),
    .B1(_01363_),
    .B2(_01362_),
    .X(_01366_));
 sky130_fd_sc_hd__o21a_1 _29797_ (.A1(_23705_),
    .A2(_23732_),
    .B1(_23734_),
    .X(_01367_));
 sky130_fd_sc_hd__o21ai_1 _29798_ (.A1(_01364_),
    .A2(_01366_),
    .B1(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__or3_1 _29799_ (.A(_01364_),
    .B(_01366_),
    .C(_01367_),
    .X(_01369_));
 sky130_fd_sc_hd__nand2_1 _29800_ (.A(_01368_),
    .B(_01369_),
    .Y(_01371_));
 sky130_fd_sc_hd__xor2_2 _29801_ (.A(_01353_),
    .B(_01371_),
    .X(_01372_));
 sky130_fd_sc_hd__o21a_1 _29802_ (.A1(_25169_),
    .A2(_25173_),
    .B1(_01372_),
    .X(_01373_));
 sky130_fd_sc_hd__a211oi_1 _29803_ (.A1(net259),
    .A2(_25171_),
    .B1(_25169_),
    .C1(_01372_),
    .Y(_01374_));
 sky130_fd_sc_hd__or2_1 _29804_ (.A(_01373_),
    .B(_01374_),
    .X(_01375_));
 sky130_fd_sc_hd__nand3_1 _29805_ (.A(_22807_),
    .B(_23737_),
    .C(_23738_),
    .Y(_01376_));
 sky130_fd_sc_hd__a21oi_1 _29806_ (.A1(_01376_),
    .A2(_23677_),
    .B1(_23740_),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _29807_ (.A(_01375_),
    .B(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__and2_1 _29808_ (.A(_01377_),
    .B(_01375_),
    .X(_01379_));
 sky130_fd_sc_hd__nor2_1 _29809_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__nand2_1 _29810_ (.A(_23643_),
    .B(_23645_),
    .Y(_01382_));
 sky130_fd_sc_hd__nor2_1 _29811_ (.A(_25173_),
    .B(_25174_),
    .Y(_01383_));
 sky130_fd_sc_hd__and3_1 _29812_ (.A(_01380_),
    .B(_01382_),
    .C(_01383_),
    .X(_01384_));
 sky130_fd_sc_hd__a21oi_1 _29813_ (.A1(_01382_),
    .A2(_01383_),
    .B1(_01380_),
    .Y(_01385_));
 sky130_fd_sc_hd__nor2_2 _29814_ (.A(_01384_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand3_1 _29815_ (.A(_01347_),
    .B(_01352_),
    .C(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__a21o_1 _29816_ (.A1(_01347_),
    .A2(_01352_),
    .B1(_01386_),
    .X(_01388_));
 sky130_fd_sc_hd__a21boi_1 _29817_ (.A1(_25186_),
    .A2(_25157_),
    .B1_N(_25152_),
    .Y(_01389_));
 sky130_fd_sc_hd__a21o_1 _29818_ (.A1(_01387_),
    .A2(_01388_),
    .B1(_01389_),
    .X(_01390_));
 sky130_fd_sc_hd__nand3_1 _29819_ (.A(_01387_),
    .B(_01388_),
    .C(_01389_),
    .Y(_01391_));
 sky130_fd_sc_hd__a21oi_1 _29820_ (.A1(_23647_),
    .A2(_25179_),
    .B1(_25178_),
    .Y(_01393_));
 sky130_fd_sc_hd__inv_2 _29821_ (.A(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__and3_1 _29822_ (.A(_01390_),
    .B(_01391_),
    .C(_01394_),
    .X(_01395_));
 sky130_fd_sc_hd__a32o_1 _29823_ (.A1(_23674_),
    .A2(_25182_),
    .A3(_25184_),
    .B1(_25190_),
    .B2(_25192_),
    .X(_01396_));
 sky130_fd_sc_hd__a21o_1 _29824_ (.A1(_01390_),
    .A2(_01391_),
    .B1(_01394_),
    .X(_01397_));
 sky130_fd_sc_hd__nand2_1 _29825_ (.A(_01396_),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand3_1 _29826_ (.A(_01390_),
    .B(_01391_),
    .C(_01394_),
    .Y(_01399_));
 sky130_fd_sc_hd__a21oi_2 _29827_ (.A1(_01397_),
    .A2(_01399_),
    .B1(_01396_),
    .Y(_01400_));
 sky130_fd_sc_hd__o21ba_1 _29828_ (.A1(_01395_),
    .A2(_01398_),
    .B1_N(_01400_),
    .X(_01401_));
 sky130_fd_sc_hd__xnor2_2 _29829_ (.A(_25205_),
    .B(_01401_),
    .Y(_00005_));
 sky130_fd_sc_hd__o211a_1 _29830_ (.A1(_24309_),
    .A2(_25129_),
    .B1(_25142_),
    .C1(_01342_),
    .X(_01403_));
 sky130_fd_sc_hd__o21ai_1 _29831_ (.A1(_25285_),
    .A2(_01403_),
    .B1(_01341_),
    .Y(_01404_));
 sky130_fd_sc_hd__and2b_1 _29832_ (.A_N(_25235_),
    .B(_25275_),
    .X(_01405_));
 sky130_fd_sc_hd__a21o_1 _29833_ (.A1(_25212_),
    .A2(_25234_),
    .B1(_01405_),
    .X(_01406_));
 sky130_fd_sc_hd__and2b_1 _29834_ (.A_N(_25249_),
    .B(_23719_),
    .X(_01407_));
 sky130_fd_sc_hd__a311o_1 _29835_ (.A1(_25247_),
    .A2(_25251_),
    .A3(_25255_),
    .B1(_01407_),
    .C1(_25252_),
    .X(_01408_));
 sky130_fd_sc_hd__buf_1 _29836_ (.A(_25249_),
    .X(_01409_));
 sky130_fd_sc_hd__or3b_1 _29837_ (.A(_01409_),
    .B(_25253_),
    .C_N(_25236_),
    .X(_01410_));
 sky130_fd_sc_hd__a21oi_1 _29838_ (.A1(_01408_),
    .A2(_01410_),
    .B1(_23721_),
    .Y(_01411_));
 sky130_fd_sc_hd__and3_1 _29839_ (.A(_23721_),
    .B(_01408_),
    .C(_01410_),
    .X(_01412_));
 sky130_fd_sc_hd__a21oi_1 _29840_ (.A1(_25258_),
    .A2(_25268_),
    .B1(_25267_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_1 _29841_ (.A(_25249_),
    .B(\delay_line[17][12] ),
    .Y(_01415_));
 sky130_fd_sc_hd__and2_1 _29842_ (.A(_25249_),
    .B(\delay_line[17][12] ),
    .X(_01416_));
 sky130_fd_sc_hd__nor2_1 _29843_ (.A(_19813_),
    .B(_18799_),
    .Y(_01417_));
 sky130_fd_sc_hd__and2_1 _29844_ (.A(_18799_),
    .B(_19813_),
    .X(_01418_));
 sky130_fd_sc_hd__o22a_1 _29845_ (.A1(_01415_),
    .A2(_01416_),
    .B1(_01417_),
    .B2(_01418_),
    .X(_01419_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29846_ (.A(_01415_),
    .X(_01420_));
 sky130_fd_sc_hd__nor4_1 _29847_ (.A(_01420_),
    .B(_01416_),
    .C(_01417_),
    .D(_01418_),
    .Y(_01421_));
 sky130_fd_sc_hd__clkbuf_2 _29848_ (.A(_23583_),
    .X(_01422_));
 sky130_fd_sc_hd__a21oi_2 _29849_ (.A1(_19795_),
    .A2(_23561_),
    .B1(_23560_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_1 _29850_ (.A(_01423_),
    .B(_23569_),
    .Y(_01425_));
 sky130_fd_sc_hd__and2_1 _29851_ (.A(_23566_),
    .B(_01423_),
    .X(_01426_));
 sky130_fd_sc_hd__nor3_1 _29852_ (.A(_01422_),
    .B(_01425_),
    .C(_01426_),
    .Y(_01427_));
 sky130_fd_sc_hd__o21a_1 _29853_ (.A1(_01425_),
    .A2(_01426_),
    .B1(_01422_),
    .X(_01428_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29854_ (.A(_20928_),
    .X(_01429_));
 sky130_fd_sc_hd__o21a_1 _29855_ (.A1(_01429_),
    .A2(_25260_),
    .B1(_25263_),
    .X(_01430_));
 sky130_fd_sc_hd__o21ai_1 _29856_ (.A1(_01427_),
    .A2(_01428_),
    .B1(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__or3_1 _29857_ (.A(_01430_),
    .B(_01427_),
    .C(_01428_),
    .X(_01432_));
 sky130_fd_sc_hd__nand2_1 _29858_ (.A(_01431_),
    .B(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__or3_1 _29859_ (.A(_01419_),
    .B(net204),
    .C(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__o21ai_1 _29860_ (.A1(_01419_),
    .A2(net205),
    .B1(_01433_),
    .Y(_01436_));
 sky130_fd_sc_hd__nand2_1 _29861_ (.A(_01434_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__xnor2_1 _29862_ (.A(_01414_),
    .B(_01437_),
    .Y(_01438_));
 sky130_fd_sc_hd__or3b_1 _29863_ (.A(_01411_),
    .B(_01412_),
    .C_N(_01438_),
    .X(_01439_));
 sky130_fd_sc_hd__o21bai_2 _29864_ (.A1(_01411_),
    .A2(_01412_),
    .B1_N(_01438_),
    .Y(_01440_));
 sky130_fd_sc_hd__nand2_2 _29865_ (.A(_01439_),
    .B(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__a21boi_2 _29866_ (.A1(_23694_),
    .A2(_25231_),
    .B1_N(_25230_),
    .Y(_01442_));
 sky130_fd_sc_hd__buf_1 _29867_ (.A(_25217_),
    .X(_01443_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _29868_ (.A(\delay_line[20][12] ),
    .X(_01444_));
 sky130_fd_sc_hd__nor2_1 _29869_ (.A(_25217_),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__and2_2 _29870_ (.A(\delay_line[20][11] ),
    .B(\delay_line[20][12] ),
    .X(_01447_));
 sky130_fd_sc_hd__nor2_2 _29871_ (.A(_01445_),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__and3_1 _29872_ (.A(_25216_),
    .B(_01443_),
    .C(_01448_),
    .X(_01449_));
 sky130_fd_sc_hd__o2bb2a_1 _29873_ (.A1_N(_25216_),
    .A2_N(_01443_),
    .B1(_01445_),
    .B2(_01447_),
    .X(_01450_));
 sky130_fd_sc_hd__xnor2_1 _29874_ (.A(_23563_),
    .B(_23685_),
    .Y(_01451_));
 sky130_fd_sc_hd__clkbuf_2 _29875_ (.A(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__nor3_2 _29876_ (.A(_01449_),
    .B(_01450_),
    .C(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__o21a_1 _29877_ (.A1(_01449_),
    .A2(_01450_),
    .B1(_01452_),
    .X(_01454_));
 sky130_fd_sc_hd__or4_1 _29878_ (.A(_15427_),
    .B(_24282_),
    .C(_01453_),
    .D(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__a2bb2o_1 _29879_ (.A1_N(_01453_),
    .A2_N(_01454_),
    .B1(_15394_),
    .B2(_24289_),
    .X(_01456_));
 sky130_fd_sc_hd__o211a_1 _29880_ (.A1(_25221_),
    .A2(_25225_),
    .B1(_01455_),
    .C1(_01456_),
    .X(_01458_));
 sky130_fd_sc_hd__a221oi_2 _29881_ (.A1(_23684_),
    .A2(_25220_),
    .B1(_01455_),
    .B2(_01456_),
    .C1(_25225_),
    .Y(_01459_));
 sky130_fd_sc_hd__a211o_1 _29882_ (.A1(_00441_),
    .A2(_00442_),
    .B1(_01458_),
    .C1(_01459_),
    .X(_01460_));
 sky130_fd_sc_hd__o211ai_1 _29883_ (.A1(_01458_),
    .A2(_01459_),
    .B1(_00441_),
    .C1(_00442_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand3_1 _29884_ (.A(_01460_),
    .B(_25228_),
    .C(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__a21o_1 _29885_ (.A1(_01461_),
    .A2(_01460_),
    .B1(_25228_),
    .X(_01463_));
 sky130_fd_sc_hd__nand2_1 _29886_ (.A(_01462_),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__xor2_1 _29887_ (.A(_01442_),
    .B(_01464_),
    .X(_01465_));
 sky130_fd_sc_hd__xor2_1 _29888_ (.A(_01441_),
    .B(_01465_),
    .X(_01466_));
 sky130_fd_sc_hd__o21ai_1 _29889_ (.A1(_25207_),
    .A2(_00461_),
    .B1(_00456_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand3_1 _29890_ (.A(_00453_),
    .B(_01466_),
    .C(_01467_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_1 _29891_ (.A(_01406_),
    .B(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__a21oi_2 _29892_ (.A1(_00452_),
    .A2(_01467_),
    .B1(_01466_),
    .Y(_01471_));
 sky130_fd_sc_hd__inv_2 _29893_ (.A(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__a21o_1 _29894_ (.A1(_01472_),
    .A2(_01469_),
    .B1(_01406_),
    .X(_01473_));
 sky130_fd_sc_hd__o21ai_2 _29895_ (.A1(_00448_),
    .A2(_00449_),
    .B1(_00430_),
    .Y(_01474_));
 sky130_fd_sc_hd__nand2_1 _29896_ (.A(_00450_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__inv_2 _29897_ (.A(_01324_),
    .Y(_01476_));
 sky130_fd_sc_hd__inv_2 _29898_ (.A(_01328_),
    .Y(_01477_));
 sky130_fd_sc_hd__a21oi_2 _29899_ (.A1(_00424_),
    .A2(_00428_),
    .B1(_00420_),
    .Y(_01478_));
 sky130_fd_sc_hd__o211a_1 _29900_ (.A1(_00305_),
    .A2(_00306_),
    .B1(_00307_),
    .C1(_00308_),
    .X(_01480_));
 sky130_fd_sc_hd__xnor2_1 _29901_ (.A(_00358_),
    .B(_00356_),
    .Y(_01481_));
 sky130_fd_sc_hd__a31oi_4 _29902_ (.A1(_00296_),
    .A2(_00301_),
    .A3(_00295_),
    .B1(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _29903_ (.A(_00345_),
    .B(_00351_),
    .Y(_01483_));
 sky130_fd_sc_hd__o21ba_1 _29904_ (.A1(_00312_),
    .A2(_00339_),
    .B1_N(_00340_),
    .X(_01484_));
 sky130_fd_sc_hd__o21bai_2 _29905_ (.A1(_00228_),
    .A2(_00245_),
    .B1_N(_00229_),
    .Y(_01485_));
 sky130_fd_sc_hd__a21oi_2 _29906_ (.A1(_00316_),
    .A2(_00336_),
    .B1(_00335_),
    .Y(_01486_));
 sky130_fd_sc_hd__or2_1 _29907_ (.A(_00241_),
    .B(_00240_),
    .X(_01487_));
 sky130_fd_sc_hd__inv_2 _29908_ (.A(_00322_),
    .Y(_01488_));
 sky130_fd_sc_hd__or2b_1 _29909_ (.A(_22023_),
    .B_N(_22235_),
    .X(_01489_));
 sky130_fd_sc_hd__xnor2_1 _29910_ (.A(_00317_),
    .B(_01489_),
    .Y(_01491_));
 sky130_fd_sc_hd__inv_2 _29911_ (.A(\delay_line[1][12] ),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_2 _29912_ (.A(net448),
    .B(_01492_),
    .Y(_01493_));
 sky130_fd_sc_hd__clkbuf_2 _29913_ (.A(\delay_line[1][12] ),
    .X(_01494_));
 sky130_fd_sc_hd__and2b_1 _29914_ (.A_N(_01494_),
    .B(net448),
    .X(_01495_));
 sky130_fd_sc_hd__nor3_1 _29915_ (.A(net441),
    .B(_01493_),
    .C(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__o21a_1 _29916_ (.A1(_01493_),
    .A2(_01495_),
    .B1(net441),
    .X(_01497_));
 sky130_fd_sc_hd__nor3b_1 _29917_ (.A(_01496_),
    .B(_01497_),
    .C_N(_00321_),
    .Y(_01498_));
 sky130_fd_sc_hd__o21ba_1 _29918_ (.A1(_01496_),
    .A2(_01497_),
    .B1_N(_00321_),
    .X(_01499_));
 sky130_fd_sc_hd__or3_1 _29919_ (.A(_01491_),
    .B(_01498_),
    .C(_01499_),
    .X(_01500_));
 sky130_fd_sc_hd__o21ai_1 _29920_ (.A1(_01498_),
    .A2(_01499_),
    .B1(_01491_),
    .Y(_01502_));
 sky130_fd_sc_hd__and4_1 _29921_ (.A(_01488_),
    .B(_00331_),
    .C(_01500_),
    .D(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__a22oi_1 _29922_ (.A1(_01488_),
    .A2(_00331_),
    .B1(_01500_),
    .B2(_01502_),
    .Y(_01504_));
 sky130_fd_sc_hd__nor2_1 _29923_ (.A(_00327_),
    .B(_00330_),
    .Y(_01505_));
 sky130_fd_sc_hd__o21ai_1 _29924_ (.A1(_01503_),
    .A2(_01504_),
    .B1(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__or3_1 _29925_ (.A(_01505_),
    .B(_01503_),
    .C(_01504_),
    .X(_01507_));
 sky130_fd_sc_hd__nand2_1 _29926_ (.A(_01506_),
    .B(_01507_),
    .Y(_01508_));
 sky130_fd_sc_hd__o211ai_1 _29927_ (.A1(_00230_),
    .A2(_00242_),
    .B1(_01487_),
    .C1(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__a21o_1 _29928_ (.A1(_01487_),
    .A2(_00243_),
    .B1(_01508_),
    .X(_01510_));
 sky130_fd_sc_hd__nand2_1 _29929_ (.A(_01509_),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__xor2_2 _29930_ (.A(_01486_),
    .B(_01511_),
    .X(_01513_));
 sky130_fd_sc_hd__xnor2_2 _29931_ (.A(_01485_),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__xor2_1 _29932_ (.A(_01484_),
    .B(_01514_),
    .X(_01515_));
 sky130_fd_sc_hd__xnor2_2 _29933_ (.A(_01483_),
    .B(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__a32o_2 _29934_ (.A1(_00288_),
    .A2(_24003_),
    .A3(_00195_),
    .B1(_00192_),
    .B2(_24112_),
    .X(_01517_));
 sky130_fd_sc_hd__nand3_2 _29935_ (.A(_00289_),
    .B(_01516_),
    .C(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__a21oi_1 _29936_ (.A1(_00289_),
    .A2(_01517_),
    .B1(_01516_),
    .Y(_01519_));
 sky130_fd_sc_hd__nor2_1 _29937_ (.A(_00354_),
    .B(_01519_),
    .Y(_01520_));
 sky130_fd_sc_hd__a21o_1 _29938_ (.A1(_00289_),
    .A2(_01517_),
    .B1(_01516_),
    .X(_01521_));
 sky130_fd_sc_hd__a32oi_4 _29939_ (.A1(_00352_),
    .A2(_00350_),
    .A3(_00351_),
    .B1(_01521_),
    .B2(_01518_),
    .Y(_01522_));
 sky130_fd_sc_hd__a21o_1 _29940_ (.A1(_01518_),
    .A2(_01520_),
    .B1(_01522_),
    .X(_01524_));
 sky130_fd_sc_hd__o21ai_1 _29941_ (.A1(_02491_),
    .A2(_17982_),
    .B1(_00130_),
    .Y(_01525_));
 sky130_fd_sc_hd__buf_1 _29942_ (.A(_00120_),
    .X(_01526_));
 sky130_fd_sc_hd__clkbuf_2 _29943_ (.A(\delay_line[12][12] ),
    .X(_01527_));
 sky130_fd_sc_hd__a21o_1 _29944_ (.A1(_00123_),
    .A2(_01526_),
    .B1(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__clkbuf_2 _29945_ (.A(_00123_),
    .X(_01529_));
 sky130_fd_sc_hd__nand3_1 _29946_ (.A(_01529_),
    .B(_01526_),
    .C(_01527_),
    .Y(_01530_));
 sky130_fd_sc_hd__a21o_1 _29947_ (.A1(_01528_),
    .A2(_01530_),
    .B1(_21805_),
    .X(_01531_));
 sky130_fd_sc_hd__nand3_1 _29948_ (.A(_01528_),
    .B(_01530_),
    .C(_21805_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _29949_ (.A(_01531_),
    .B(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__xnor2_1 _29950_ (.A(_01525_),
    .B(_01533_),
    .Y(_01535_));
 sky130_fd_sc_hd__a21boi_1 _29951_ (.A1(_23886_),
    .A2(_00109_),
    .B1_N(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__buf_2 _29952_ (.A(_00092_),
    .X(_01537_));
 sky130_fd_sc_hd__and4b_1 _29953_ (.A_N(_01535_),
    .B(_00109_),
    .C(_23880_),
    .D(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__nor2_1 _29954_ (.A(_01536_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__and2_1 _29955_ (.A(_01539_),
    .B(_00132_),
    .X(_01540_));
 sky130_fd_sc_hd__nor2_1 _29956_ (.A(_00132_),
    .B(_01539_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _29957_ (.A(_00079_),
    .B(_00080_),
    .Y(_01542_));
 sky130_fd_sc_hd__a21oi_1 _29958_ (.A1(_00070_),
    .A2(_00072_),
    .B1(_00068_),
    .Y(_01543_));
 sky130_fd_sc_hd__o21ai_2 _29959_ (.A1(_01542_),
    .A2(_01543_),
    .B1(_00074_),
    .Y(_01544_));
 sky130_fd_sc_hd__or2_1 _29960_ (.A(\delay_line[0][8] ),
    .B(\delay_line[13][12] ),
    .X(_01546_));
 sky130_fd_sc_hd__buf_1 _29961_ (.A(\delay_line[13][12] ),
    .X(_01547_));
 sky130_fd_sc_hd__nand2_2 _29962_ (.A(_21736_),
    .B(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__clkbuf_2 _29963_ (.A(\delay_line[13][11] ),
    .X(_01549_));
 sky130_fd_sc_hd__and4_1 _29964_ (.A(_01546_),
    .B(_01548_),
    .C(_21746_),
    .D(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__a22o_1 _29965_ (.A1(_21746_),
    .A2(_01549_),
    .B1(_01546_),
    .B2(_01548_),
    .X(_01551_));
 sky130_fd_sc_hd__inv_2 _29966_ (.A(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__a211o_1 _29967_ (.A1(_22313_),
    .A2(_23838_),
    .B1(_25430_),
    .C1(_00049_),
    .X(_01553_));
 sky130_fd_sc_hd__and2_2 _29968_ (.A(_21718_),
    .B(\delay_line[11][10] ),
    .X(_01554_));
 sky130_fd_sc_hd__clkbuf_2 _29969_ (.A(\delay_line[11][10] ),
    .X(_01555_));
 sky130_fd_sc_hd__nor2_1 _29970_ (.A(_01555_),
    .B(_21728_),
    .Y(_01557_));
 sky130_fd_sc_hd__nor2b_1 _29971_ (.A(_20003_),
    .B_N(_25433_),
    .Y(_01558_));
 sky130_fd_sc_hd__a21o_1 _29972_ (.A1(_25436_),
    .A2(_00049_),
    .B1(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__o21bai_2 _29973_ (.A1(_01554_),
    .A2(_01557_),
    .B1_N(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__or2_1 _29974_ (.A(_01555_),
    .B(_21728_),
    .X(_01561_));
 sky130_fd_sc_hd__nand3b_1 _29975_ (.A_N(_01554_),
    .B(_01561_),
    .C(_01559_),
    .Y(_01562_));
 sky130_fd_sc_hd__clkbuf_2 _29976_ (.A(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__nand2_2 _29977_ (.A(_01560_),
    .B(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__a211oi_2 _29978_ (.A1(_25438_),
    .A2(_25440_),
    .B1(_23844_),
    .C1(_23845_),
    .Y(_01565_));
 sky130_fd_sc_hd__nand2_1 _29979_ (.A(_01565_),
    .B(_23849_),
    .Y(_01566_));
 sky130_fd_sc_hd__o211a_1 _29980_ (.A1(_01553_),
    .A2(_25437_),
    .B1(_01564_),
    .C1(_01566_),
    .X(_01568_));
 sky130_fd_sc_hd__a22oi_4 _29981_ (.A1(_23844_),
    .A2(_25439_),
    .B1(_01565_),
    .B2(_23848_),
    .Y(_01569_));
 sky130_fd_sc_hd__buf_6 _29982_ (.A(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__nor2_1 _29983_ (.A(_01564_),
    .B(_01570_),
    .Y(_01571_));
 sky130_fd_sc_hd__a21oi_4 _29984_ (.A1(_25409_),
    .A2(_25410_),
    .B1(_25426_),
    .Y(_01572_));
 sky130_fd_sc_hd__and2b_2 _29985_ (.A_N(\delay_line[4][6] ),
    .B(\delay_line[4][8] ),
    .X(_01573_));
 sky130_fd_sc_hd__a21oi_4 _29986_ (.A1(_25418_),
    .A2(_25419_),
    .B1(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2b_1 _29987_ (.A_N(\delay_line[4][7] ),
    .B(\delay_line[4][9] ),
    .Y(_01575_));
 sky130_fd_sc_hd__nand2b_1 _29988_ (.A_N(\delay_line[4][9] ),
    .B(\delay_line[4][7] ),
    .Y(_01576_));
 sky130_fd_sc_hd__and2_1 _29989_ (.A(_01575_),
    .B(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__buf_2 _29990_ (.A(_01577_),
    .X(_01579_));
 sky130_fd_sc_hd__xnor2_2 _29991_ (.A(_01574_),
    .B(_01579_),
    .Y(_01580_));
 sky130_fd_sc_hd__clkbuf_2 _29992_ (.A(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__and4_2 _29993_ (.A(_25416_),
    .B(_25412_),
    .C(_23828_),
    .D(_23829_),
    .X(_01582_));
 sky130_fd_sc_hd__nor2_1 _29994_ (.A(_01581_),
    .B(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__o21ai_4 _29995_ (.A1(_25423_),
    .A2(_01572_),
    .B1(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_1 _29996_ (.A(_25411_),
    .B(_25415_),
    .Y(_01585_));
 sky130_fd_sc_hd__o21ai_4 _29997_ (.A1(_25421_),
    .A2(_25422_),
    .B1(_01580_),
    .Y(_01586_));
 sky130_fd_sc_hd__inv_2 _29998_ (.A(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__a22oi_1 _29999_ (.A1(_01581_),
    .A2(_01582_),
    .B1(_01585_),
    .B2(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__a2bb2oi_2 _30000_ (.A1_N(_01568_),
    .A2_N(_01571_),
    .B1(_01584_),
    .B2(_01588_),
    .Y(_01590_));
 sky130_fd_sc_hd__xor2_4 _30001_ (.A(_01574_),
    .B(_01579_),
    .X(_01591_));
 sky130_fd_sc_hd__nand4_2 _30002_ (.A(_25416_),
    .B(_25412_),
    .C(_23828_),
    .D(_23829_),
    .Y(_01592_));
 sky130_fd_sc_hd__o22ai_4 _30003_ (.A1(_01591_),
    .A2(_01592_),
    .B1(_01586_),
    .B2(_01572_),
    .Y(_01593_));
 sky130_fd_sc_hd__nand2_1 _30004_ (.A(_01570_),
    .B(_01564_),
    .Y(_01594_));
 sky130_fd_sc_hd__a221o_1 _30005_ (.A1(_22310_),
    .A2(_23837_),
    .B1(_25431_),
    .B2(_23840_),
    .C1(_22304_),
    .X(_01595_));
 sky130_fd_sc_hd__nand3_1 _30006_ (.A(_01553_),
    .B(_01595_),
    .C(_25441_),
    .Y(_01596_));
 sky130_fd_sc_hd__o22ai_2 _30007_ (.A1(_01553_),
    .A2(_25437_),
    .B1(_01596_),
    .B2(_23859_),
    .Y(_01597_));
 sky130_fd_sc_hd__and2_1 _30008_ (.A(_01560_),
    .B(_01563_),
    .X(_01598_));
 sky130_fd_sc_hd__nand2_1 _30009_ (.A(_01597_),
    .B(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__nand2_1 _30010_ (.A(_01594_),
    .B(_01599_),
    .Y(_01601_));
 sky130_fd_sc_hd__nor3b_4 _30011_ (.A(_01593_),
    .B(_01601_),
    .C_N(_01584_),
    .Y(_01602_));
 sky130_fd_sc_hd__o21bai_2 _30012_ (.A1(_01590_),
    .A2(_01602_),
    .B1_N(net454),
    .Y(_01603_));
 sky130_fd_sc_hd__o21bai_4 _30013_ (.A1(_25426_),
    .A2(_25428_),
    .B1_N(_01586_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _30014_ (.A(_01581_),
    .B(_01582_),
    .Y(_01605_));
 sky130_fd_sc_hd__nand3_1 _30015_ (.A(_01584_),
    .B(_01604_),
    .C(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__o21ai_2 _30016_ (.A1(_01568_),
    .A2(_01571_),
    .B1(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__nor2_1 _30017_ (.A(_01568_),
    .B(_01571_),
    .Y(_01608_));
 sky130_fd_sc_hd__o2111ai_4 _30018_ (.A1(_00042_),
    .A2(_01591_),
    .B1(_01584_),
    .C1(_01605_),
    .D1(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand3_1 _30019_ (.A(_01607_),
    .B(_01609_),
    .C(net454),
    .Y(_01610_));
 sky130_fd_sc_hd__a22oi_2 _30020_ (.A1(_00055_),
    .A2(_00043_),
    .B1(_01603_),
    .B2(_01610_),
    .Y(_01612_));
 sky130_fd_sc_hd__a21oi_1 _30021_ (.A1(_00042_),
    .A2(_01583_),
    .B1(_01593_),
    .Y(_01613_));
 sky130_fd_sc_hd__o21ai_1 _30022_ (.A1(_01608_),
    .A2(_01613_),
    .B1(net454),
    .Y(_01614_));
 sky130_fd_sc_hd__o21a_1 _30023_ (.A1(_00046_),
    .A2(_00045_),
    .B1(_00055_),
    .X(_01615_));
 sky130_fd_sc_hd__o211a_2 _30024_ (.A1(_01614_),
    .A2(_01602_),
    .B1(_01615_),
    .C1(_01603_),
    .X(_01616_));
 sky130_fd_sc_hd__clkbuf_2 _30025_ (.A(_00046_),
    .X(_01617_));
 sky130_fd_sc_hd__o21bai_4 _30026_ (.A1(_01612_),
    .A2(_01616_),
    .B1_N(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__o21ai_1 _30027_ (.A1(_01602_),
    .A2(_01614_),
    .B1(_01603_),
    .Y(_01619_));
 sky130_fd_sc_hd__a21o_1 _30028_ (.A1(_01603_),
    .A2(_01610_),
    .B1(_01615_),
    .X(_01620_));
 sky130_fd_sc_hd__o211ai_2 _30029_ (.A1(_00041_),
    .A2(_01619_),
    .B1(_01617_),
    .C1(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__o211a_1 _30030_ (.A1(_00056_),
    .A2(_00045_),
    .B1(_23865_),
    .C1(_00057_),
    .X(_01623_));
 sky130_fd_sc_hd__a21o_1 _30031_ (.A1(_00077_),
    .A2(_00048_),
    .B1(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__a21oi_2 _30032_ (.A1(_01618_),
    .A2(_01621_),
    .B1(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__inv_2 _30033_ (.A(net454),
    .Y(_01626_));
 sky130_fd_sc_hd__a21oi_1 _30034_ (.A1(_01601_),
    .A2(_01606_),
    .B1(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__nand2_1 _30035_ (.A(_01607_),
    .B(_01609_),
    .Y(_01628_));
 sky130_fd_sc_hd__a22oi_1 _30036_ (.A1(_01627_),
    .A2(_01609_),
    .B1(_01626_),
    .B2(_01628_),
    .Y(_01629_));
 sky130_fd_sc_hd__clkbuf_2 _30037_ (.A(_01617_),
    .X(_01630_));
 sky130_fd_sc_hd__o21ai_2 _30038_ (.A1(_01615_),
    .A2(_01629_),
    .B1(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__o221a_1 _30039_ (.A1(_01623_),
    .A2(_00071_),
    .B1(_01616_),
    .B2(_01631_),
    .C1(_01618_),
    .X(_01632_));
 sky130_fd_sc_hd__o22ai_2 _30040_ (.A1(_01550_),
    .A2(_01552_),
    .B1(_01625_),
    .B2(_01632_),
    .Y(_01634_));
 sky130_fd_sc_hd__nand4_4 _30041_ (.A(_01546_),
    .B(_01548_),
    .C(_19986_),
    .D(\delay_line[13][11] ),
    .Y(_01635_));
 sky130_fd_sc_hd__nand2_1 _30042_ (.A(_01635_),
    .B(_01551_),
    .Y(_01636_));
 sky130_fd_sc_hd__a21o_1 _30043_ (.A1(_01618_),
    .A2(_01621_),
    .B1(_01624_),
    .X(_01637_));
 sky130_fd_sc_hd__o221ai_4 _30044_ (.A1(_01623_),
    .A2(_00071_),
    .B1(_01616_),
    .B2(_01631_),
    .C1(_01618_),
    .Y(_01638_));
 sky130_fd_sc_hd__nand3b_2 _30045_ (.A_N(_01636_),
    .B(_01637_),
    .C(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__nand3_2 _30046_ (.A(_01544_),
    .B(_01634_),
    .C(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__o21bai_1 _30047_ (.A1(_01625_),
    .A2(_01632_),
    .B1_N(_01636_),
    .Y(_01641_));
 sky130_fd_sc_hd__o32a_1 _30048_ (.A1(_00067_),
    .A2(_00061_),
    .A3(_00066_),
    .B1(_01542_),
    .B2(_01543_),
    .X(_01642_));
 sky130_fd_sc_hd__o211ai_1 _30049_ (.A1(_01550_),
    .A2(_01552_),
    .B1(_01637_),
    .C1(_01638_),
    .Y(_01643_));
 sky130_fd_sc_hd__nand3_1 _30050_ (.A(_01641_),
    .B(_01642_),
    .C(_01643_),
    .Y(_01645_));
 sky130_fd_sc_hd__and3_1 _30051_ (.A(_22362_),
    .B(_23879_),
    .C(_00093_),
    .X(_01646_));
 sky130_fd_sc_hd__nand2_1 _30052_ (.A(_18918_),
    .B(_00093_),
    .Y(_01647_));
 sky130_fd_sc_hd__or2_1 _30053_ (.A(_18918_),
    .B(\delay_line[13][10] ),
    .X(_01648_));
 sky130_fd_sc_hd__and3_1 _30054_ (.A(_00082_),
    .B(_01647_),
    .C(_01648_),
    .X(_01649_));
 sky130_fd_sc_hd__a21oi_2 _30055_ (.A1(_01647_),
    .A2(_01648_),
    .B1(_00082_),
    .Y(_01650_));
 sky130_fd_sc_hd__a2111oi_1 _30056_ (.A1(_00094_),
    .A2(_00099_),
    .B1(_01646_),
    .C1(_01649_),
    .D1(_01650_),
    .Y(_01651_));
 sky130_fd_sc_hd__o22a_1 _30057_ (.A1(_01646_),
    .A2(_00098_),
    .B1(_01649_),
    .B2(_01650_),
    .X(_01652_));
 sky130_fd_sc_hd__o2bb2ai_1 _30058_ (.A1_N(_01640_),
    .A2_N(_01645_),
    .B1(net257),
    .B2(_01652_),
    .Y(_01653_));
 sky130_fd_sc_hd__a32oi_2 _30059_ (.A1(_00086_),
    .A2(_00089_),
    .A3(_00090_),
    .B1(_00115_),
    .B2(_00149_),
    .Y(_01654_));
 sky130_fd_sc_hd__a21oi_1 _30060_ (.A1(_00094_),
    .A2(_18962_),
    .B1(_01646_),
    .Y(_01656_));
 sky130_fd_sc_hd__nor3_1 _30061_ (.A(_01656_),
    .B(_01649_),
    .C(_01650_),
    .Y(_01657_));
 sky130_fd_sc_hd__o21a_1 _30062_ (.A1(_01649_),
    .A2(_01650_),
    .B1(_01656_),
    .X(_01658_));
 sky130_fd_sc_hd__clkbuf_2 _30063_ (.A(_01645_),
    .X(_01659_));
 sky130_fd_sc_hd__o211ai_1 _30064_ (.A1(net256),
    .A2(_01658_),
    .B1(_01640_),
    .C1(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand3_1 _30065_ (.A(_01653_),
    .B(_01654_),
    .C(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__clkbuf_2 _30066_ (.A(_01661_),
    .X(_01662_));
 sky130_fd_sc_hd__o21ai_1 _30067_ (.A1(_01540_),
    .A2(_01541_),
    .B1(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__a32o_1 _30068_ (.A1(_00086_),
    .A2(_00089_),
    .A3(_00090_),
    .B1(_00115_),
    .B2(_00149_),
    .X(_01664_));
 sky130_fd_sc_hd__o2bb2ai_1 _30069_ (.A1_N(_01640_),
    .A2_N(_01659_),
    .B1(net256),
    .B2(_01658_),
    .Y(_01665_));
 sky130_fd_sc_hd__o211ai_2 _30070_ (.A1(net257),
    .A2(_01652_),
    .B1(_01640_),
    .C1(_01659_),
    .Y(_01667_));
 sky130_fd_sc_hd__and3_1 _30071_ (.A(_01664_),
    .B(_01665_),
    .C(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__a2bb2o_1 _30072_ (.A1_N(_00151_),
    .A2_N(_00152_),
    .B1(_00142_),
    .B2(_00114_),
    .X(_01669_));
 sky130_fd_sc_hd__nand3_1 _30073_ (.A(_01664_),
    .B(_01665_),
    .C(_01667_),
    .Y(_01670_));
 sky130_fd_sc_hd__and4_1 _30074_ (.A(_00125_),
    .B(_00127_),
    .C(_00129_),
    .D(_00131_),
    .X(_01671_));
 sky130_fd_sc_hd__and2_1 _30075_ (.A(_01671_),
    .B(_01539_),
    .X(_01672_));
 sky130_fd_sc_hd__nor2_1 _30076_ (.A(_01671_),
    .B(_01539_),
    .Y(_01673_));
 sky130_fd_sc_hd__o2bb2ai_1 _30077_ (.A1_N(_01670_),
    .A2_N(_01662_),
    .B1(_01672_),
    .B2(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__o211ai_2 _30078_ (.A1(_01663_),
    .A2(_01668_),
    .B1(_01669_),
    .C1(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__o2bb2ai_1 _30079_ (.A1_N(_01670_),
    .A2_N(_01661_),
    .B1(_01540_),
    .B2(_01541_),
    .Y(_01676_));
 sky130_fd_sc_hd__o2bb2a_1 _30080_ (.A1_N(_00142_),
    .A2_N(_00113_),
    .B1(_00152_),
    .B2(_00151_),
    .X(_01678_));
 sky130_fd_sc_hd__o211ai_1 _30081_ (.A1(_01672_),
    .A2(_01673_),
    .B1(_01670_),
    .C1(_01662_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand3_1 _30082_ (.A(_01676_),
    .B(_01678_),
    .C(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__inv_2 _30083_ (.A(net417),
    .Y(_01681_));
 sky130_fd_sc_hd__buf_1 _30084_ (.A(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__or2_1 _30085_ (.A(_25396_),
    .B(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__nand2_1 _30086_ (.A(_01682_),
    .B(_25396_),
    .Y(_01684_));
 sky130_fd_sc_hd__a21oi_1 _30087_ (.A1(_01683_),
    .A2(_01684_),
    .B1(_25386_),
    .Y(_01685_));
 sky130_fd_sc_hd__and3_1 _30088_ (.A(_01683_),
    .B(_01684_),
    .C(_25386_),
    .X(_01686_));
 sky130_fd_sc_hd__nor3_2 _30089_ (.A(_01685_),
    .B(_25393_),
    .C(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__o21a_1 _30090_ (.A1(_01686_),
    .A2(_01685_),
    .B1(_25393_),
    .X(_01689_));
 sky130_fd_sc_hd__or2_1 _30091_ (.A(_22447_),
    .B(_19956_),
    .X(_01690_));
 sky130_fd_sc_hd__nand2_1 _30092_ (.A(_19964_),
    .B(_25392_),
    .Y(_01691_));
 sky130_fd_sc_hd__clkbuf_2 _30093_ (.A(_23771_),
    .X(_01692_));
 sky130_fd_sc_hd__nand3_1 _30094_ (.A(_01690_),
    .B(_01691_),
    .C(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__clkbuf_2 _30095_ (.A(_01692_),
    .X(_01694_));
 sky130_fd_sc_hd__a21o_1 _30096_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__and3b_1 _30097_ (.A_N(_25387_),
    .B(_01693_),
    .C(_01695_),
    .X(_01696_));
 sky130_fd_sc_hd__a21boi_1 _30098_ (.A1(_01693_),
    .A2(_01695_),
    .B1_N(_25387_),
    .Y(_01697_));
 sky130_fd_sc_hd__or4_1 _30099_ (.A(_01687_),
    .B(_01689_),
    .C(_01696_),
    .D(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__o22ai_1 _30100_ (.A1(_01687_),
    .A2(_01689_),
    .B1(_01696_),
    .B2(_01697_),
    .Y(_01700_));
 sky130_fd_sc_hd__nand2_1 _30101_ (.A(_01698_),
    .B(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__clkbuf_2 _30102_ (.A(_25376_),
    .X(_01702_));
 sky130_fd_sc_hd__and3b_1 _30103_ (.A_N(_01526_),
    .B(_23800_),
    .C(_23799_),
    .X(_01703_));
 sky130_fd_sc_hd__o211a_1 _30104_ (.A1(_23800_),
    .A2(_01526_),
    .B1(_18985_),
    .C1(_00122_),
    .X(_01704_));
 sky130_fd_sc_hd__and2_1 _30105_ (.A(_18984_),
    .B(\delay_line[10][12] ),
    .X(_01705_));
 sky130_fd_sc_hd__nor2_1 _30106_ (.A(_18984_),
    .B(\delay_line[10][12] ),
    .Y(_01706_));
 sky130_fd_sc_hd__nand4bb_1 _30107_ (.A_N(_01705_),
    .B_N(_01706_),
    .C(_18987_),
    .D(_25375_),
    .Y(_01707_));
 sky130_fd_sc_hd__a2bb2o_1 _30108_ (.A1_N(_01705_),
    .A2_N(_01706_),
    .B1(_18988_),
    .B2(_25376_),
    .X(_01708_));
 sky130_fd_sc_hd__o211a_1 _30109_ (.A1(_01703_),
    .A2(_01704_),
    .B1(_01707_),
    .C1(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__buf_1 _30110_ (.A(_01707_),
    .X(_01711_));
 sky130_fd_sc_hd__a221oi_1 _30111_ (.A1(_18986_),
    .A2(_00126_),
    .B1(_01711_),
    .B2(_01708_),
    .C1(_01703_),
    .Y(_01712_));
 sky130_fd_sc_hd__or4_1 _30112_ (.A(_01702_),
    .B(_17995_),
    .C(_01709_),
    .D(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__o22ai_1 _30113_ (.A1(_01702_),
    .A2(_17995_),
    .B1(_01709_),
    .B2(_01712_),
    .Y(_01714_));
 sky130_fd_sc_hd__a31o_1 _30114_ (.A1(_23769_),
    .A2(_22460_),
    .A3(_25381_),
    .B1(_25378_),
    .X(_01715_));
 sky130_fd_sc_hd__a21oi_1 _30115_ (.A1(_01713_),
    .A2(_01714_),
    .B1(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__and3_1 _30116_ (.A(_01715_),
    .B(_01713_),
    .C(_01714_),
    .X(_01717_));
 sky130_fd_sc_hd__nor2_1 _30117_ (.A(_01716_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__xor2_2 _30118_ (.A(_01701_),
    .B(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__a21oi_2 _30119_ (.A1(_00135_),
    .A2(_00137_),
    .B1(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__or3b_1 _30120_ (.A(_00136_),
    .B(_00138_),
    .C_N(_01719_),
    .X(_01722_));
 sky130_fd_sc_hd__a32o_1 _30121_ (.A1(_25384_),
    .A2(_25400_),
    .A3(_25401_),
    .B1(_25382_),
    .B2(_25383_),
    .X(_01723_));
 sky130_fd_sc_hd__inv_2 _30122_ (.A(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__and3b_1 _30123_ (.A_N(_01720_),
    .B(_01722_),
    .C(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__and2b_1 _30124_ (.A_N(_01720_),
    .B(_01722_),
    .X(_01726_));
 sky130_fd_sc_hd__nor2_1 _30125_ (.A(_01724_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__o2bb2ai_1 _30126_ (.A1_N(_01675_),
    .A2_N(_01680_),
    .B1(_01725_),
    .B2(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__nor2_1 _30127_ (.A(_00162_),
    .B(_00163_),
    .Y(_01729_));
 sky130_fd_sc_hd__a21oi_1 _30128_ (.A1(_00173_),
    .A2(_01729_),
    .B1(_00148_),
    .Y(_01730_));
 sky130_fd_sc_hd__and2_2 _30129_ (.A(_01726_),
    .B(_01723_),
    .X(_01731_));
 sky130_fd_sc_hd__nor2_1 _30130_ (.A(_01723_),
    .B(_01726_),
    .Y(_01733_));
 sky130_fd_sc_hd__clkbuf_2 _30131_ (.A(_01680_),
    .X(_01734_));
 sky130_fd_sc_hd__o211ai_1 _30132_ (.A1(_01731_),
    .A2(_01733_),
    .B1(_01675_),
    .C1(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__nand3_1 _30133_ (.A(_01728_),
    .B(_01730_),
    .C(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__clkbuf_2 _30134_ (.A(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__a21oi_1 _30135_ (.A1(_25368_),
    .A2(_25405_),
    .B1(_00160_),
    .Y(_01738_));
 sky130_fd_sc_hd__buf_1 _30136_ (.A(_21869_),
    .X(_01739_));
 sky130_fd_sc_hd__buf_1 _30137_ (.A(_25313_),
    .X(_01740_));
 sky130_fd_sc_hd__clkbuf_2 _30138_ (.A(_23943_),
    .X(_01741_));
 sky130_fd_sc_hd__and3_1 _30139_ (.A(_01739_),
    .B(_01740_),
    .C(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__buf_1 _30140_ (.A(\delay_line[7][12] ),
    .X(_01744_));
 sky130_fd_sc_hd__clkbuf_2 _30141_ (.A(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__or2_1 _30142_ (.A(_01745_),
    .B(_11833_),
    .X(_01746_));
 sky130_fd_sc_hd__buf_2 _30143_ (.A(_25297_),
    .X(_01747_));
 sky130_fd_sc_hd__nand2_2 _30144_ (.A(_11866_),
    .B(_01745_),
    .Y(_01748_));
 sky130_fd_sc_hd__nand4_4 _30145_ (.A(_18844_),
    .B(_01746_),
    .C(_01747_),
    .D(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__a22o_1 _30146_ (.A1(_25297_),
    .A2(_18844_),
    .B1(_01746_),
    .B2(_01748_),
    .X(_01750_));
 sky130_fd_sc_hd__o211a_1 _30147_ (.A1(_01742_),
    .A2(_25319_),
    .B1(_01749_),
    .C1(_01750_),
    .X(_01751_));
 sky130_fd_sc_hd__a221oi_2 _30148_ (.A1(_25318_),
    .A2(_18044_),
    .B1(_01750_),
    .B2(_01749_),
    .C1(_01742_),
    .Y(_01752_));
 sky130_fd_sc_hd__nor3_1 _30149_ (.A(_25300_),
    .B(_01751_),
    .C(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__o21a_1 _30150_ (.A1(_01751_),
    .A2(_01752_),
    .B1(_25300_),
    .X(_01755_));
 sky130_fd_sc_hd__nor2_2 _30151_ (.A(_01753_),
    .B(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__clkbuf_2 _30152_ (.A(_25308_),
    .X(_01757_));
 sky130_fd_sc_hd__o21ai_2 _30153_ (.A1(_23943_),
    .A2(_25311_),
    .B1(_25313_),
    .Y(_01758_));
 sky130_fd_sc_hd__a21o_1 _30154_ (.A1(_01741_),
    .A2(_01757_),
    .B1(_01758_),
    .X(_01759_));
 sky130_fd_sc_hd__clkbuf_2 _30155_ (.A(\delay_line[8][10] ),
    .X(_01760_));
 sky130_fd_sc_hd__and2_1 _30156_ (.A(_01760_),
    .B(_25311_),
    .X(_01761_));
 sky130_fd_sc_hd__nor2_1 _30157_ (.A(_01760_),
    .B(_01757_),
    .Y(_01762_));
 sky130_fd_sc_hd__o21bai_2 _30158_ (.A1(_01761_),
    .A2(_01762_),
    .B1_N(_25313_),
    .Y(_01763_));
 sky130_fd_sc_hd__a21o_1 _30159_ (.A1(_01759_),
    .A2(_01763_),
    .B1(_23947_),
    .X(_01764_));
 sky130_fd_sc_hd__o211ai_4 _30160_ (.A1(_01758_),
    .A2(_01761_),
    .B1(_23947_),
    .C1(_01763_),
    .Y(_01766_));
 sky130_fd_sc_hd__clkbuf_2 _30161_ (.A(_20099_),
    .X(_01767_));
 sky130_fd_sc_hd__a21o_1 _30162_ (.A1(_01764_),
    .A2(_01766_),
    .B1(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__nand3_2 _30163_ (.A(_01764_),
    .B(_01766_),
    .C(_01767_),
    .Y(_01769_));
 sky130_fd_sc_hd__buf_1 _30164_ (.A(\delay_line[8][12] ),
    .X(_01770_));
 sky130_fd_sc_hd__clkbuf_2 _30165_ (.A(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__xnor2_2 _30166_ (.A(_12987_),
    .B(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__nor2_1 _30167_ (.A(_25309_),
    .B(_25312_),
    .Y(_01773_));
 sky130_fd_sc_hd__a21oi_1 _30168_ (.A1(_18054_),
    .A2(_01773_),
    .B1(_25310_),
    .Y(_01774_));
 sky130_fd_sc_hd__xnor2_1 _30169_ (.A(_01772_),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__a21oi_1 _30170_ (.A1(_01768_),
    .A2(_01769_),
    .B1(_01775_),
    .Y(_01777_));
 sky130_fd_sc_hd__and3_1 _30171_ (.A(_01775_),
    .B(_01768_),
    .C(_01769_),
    .X(_01778_));
 sky130_fd_sc_hd__nor2_1 _30172_ (.A(_01777_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__a31o_1 _30173_ (.A1(_18058_),
    .A2(_22502_),
    .A3(_01773_),
    .B1(_25323_),
    .X(_01780_));
 sky130_fd_sc_hd__nand2_1 _30174_ (.A(_01779_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__a311o_1 _30175_ (.A1(_18058_),
    .A2(_22502_),
    .A3(_01773_),
    .B1(_25323_),
    .C1(_01779_),
    .X(_01782_));
 sky130_fd_sc_hd__nand2_2 _30176_ (.A(_01781_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__xor2_4 _30177_ (.A(_01756_),
    .B(_01783_),
    .X(_01784_));
 sky130_fd_sc_hd__o2bb2a_1 _30178_ (.A1_N(_23752_),
    .A2_N(_23754_),
    .B1(_25340_),
    .B2(_25343_),
    .X(_01785_));
 sky130_fd_sc_hd__nor2_1 _30179_ (.A(_23978_),
    .B(_23975_),
    .Y(_01786_));
 sky130_fd_sc_hd__clkbuf_2 _30180_ (.A(_23969_),
    .X(_01788_));
 sky130_fd_sc_hd__clkbuf_2 _30181_ (.A(_25337_),
    .X(_01789_));
 sky130_fd_sc_hd__and4bb_1 _30182_ (.A_N(_01786_),
    .B_N(_25346_),
    .C(_01788_),
    .D(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__nand2_1 _30183_ (.A(_25389_),
    .B(_25401_),
    .Y(_01791_));
 sky130_fd_sc_hd__a21oi_1 _30184_ (.A1(_25339_),
    .A2(_25337_),
    .B1(_17916_),
    .Y(_01792_));
 sky130_fd_sc_hd__xnor2_4 _30185_ (.A(_23971_),
    .B(net418),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _30186_ (.A(_25339_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__or3b_1 _30187_ (.A(_22436_),
    .B(net418),
    .C_N(_23971_),
    .X(_01795_));
 sky130_fd_sc_hd__a21oi_2 _30188_ (.A1(_01794_),
    .A2(_01795_),
    .B1(_20123_),
    .Y(_01796_));
 sky130_fd_sc_hd__and3_2 _30189_ (.A(_01795_),
    .B(_20123_),
    .C(_01794_),
    .X(_01797_));
 sky130_fd_sc_hd__a211oi_4 _30190_ (.A1(_25397_),
    .A2(_25398_),
    .B1(_01796_),
    .C1(_01797_),
    .Y(_01799_));
 sky130_fd_sc_hd__o211a_1 _30191_ (.A1(_01796_),
    .A2(_01797_),
    .B1(_25397_),
    .C1(_25398_),
    .X(_01800_));
 sky130_fd_sc_hd__nor4_1 _30192_ (.A(_23978_),
    .B(_01792_),
    .C(_01799_),
    .D(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__o22a_1 _30193_ (.A1(_23978_),
    .A2(_01792_),
    .B1(_01799_),
    .B2(_01800_),
    .X(_01802_));
 sky130_fd_sc_hd__nor2_1 _30194_ (.A(_01801_),
    .B(_01802_),
    .Y(_01803_));
 sky130_fd_sc_hd__or2_1 _30195_ (.A(_01791_),
    .B(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__a211oi_2 _30196_ (.A1(_25389_),
    .A2(_25401_),
    .B1(_01801_),
    .C1(_01802_),
    .Y(_01805_));
 sky130_fd_sc_hd__inv_2 _30197_ (.A(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__o211a_1 _30198_ (.A1(_01785_),
    .A2(_01790_),
    .B1(_01804_),
    .C1(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__a221oi_1 _30199_ (.A1(_25344_),
    .A2(_25345_),
    .B1(_01804_),
    .B2(_01806_),
    .C1(_01790_),
    .Y(_01808_));
 sky130_fd_sc_hd__nor2_1 _30200_ (.A(_01807_),
    .B(_01808_),
    .Y(_01810_));
 sky130_fd_sc_hd__a21bo_1 _30201_ (.A1(_25334_),
    .A2(_25349_),
    .B1_N(_25350_),
    .X(_01811_));
 sky130_fd_sc_hd__nand2_1 _30202_ (.A(_01810_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__or2_1 _30203_ (.A(_01811_),
    .B(_01810_),
    .X(_01813_));
 sky130_fd_sc_hd__nand2_1 _30204_ (.A(_01812_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__xnor2_2 _30205_ (.A(_01784_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__a22o_1 _30206_ (.A1(_25354_),
    .A2(_25356_),
    .B1(_01738_),
    .B2(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__o21ba_1 _30207_ (.A1(_01738_),
    .A2(_01815_),
    .B1_N(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__or2b_1 _30208_ (.A(_01738_),
    .B_N(_01815_),
    .X(_01818_));
 sky130_fd_sc_hd__a211o_1 _30209_ (.A1(_25368_),
    .A2(_25405_),
    .B1(_00162_),
    .C1(_01815_),
    .X(_01819_));
 sky130_fd_sc_hd__and4_1 _30210_ (.A(_25354_),
    .B(_25356_),
    .C(_01818_),
    .D(_01819_),
    .X(_01821_));
 sky130_fd_sc_hd__nor2_2 _30211_ (.A(_01817_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__nand2_1 _30212_ (.A(_01737_),
    .B(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__nor2_1 _30213_ (.A(_01731_),
    .B(_01733_),
    .Y(_01824_));
 sky130_fd_sc_hd__nand2_1 _30214_ (.A(_01734_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__o211a_2 _30215_ (.A1(_01663_),
    .A2(_01668_),
    .B1(_01669_),
    .C1(_01674_),
    .X(_01826_));
 sky130_fd_sc_hd__a22o_1 _30216_ (.A1(_00154_),
    .A2(_00170_),
    .B1(_00173_),
    .B2(_01729_),
    .X(_01827_));
 sky130_fd_sc_hd__o2bb2ai_2 _30217_ (.A1_N(_01675_),
    .A2_N(_01734_),
    .B1(_01731_),
    .B2(_01733_),
    .Y(_01828_));
 sky130_fd_sc_hd__o211a_2 _30218_ (.A1(_01825_),
    .A2(_01826_),
    .B1(_01827_),
    .C1(_01828_),
    .X(_01829_));
 sky130_fd_sc_hd__a22o_1 _30219_ (.A1(_00175_),
    .A2(_00174_),
    .B1(_00169_),
    .B2(_00184_),
    .X(_01830_));
 sky130_fd_sc_hd__o211ai_4 _30220_ (.A1(_01825_),
    .A2(_01826_),
    .B1(_01827_),
    .C1(_01828_),
    .Y(_01832_));
 sky130_fd_sc_hd__o2bb2ai_2 _30221_ (.A1_N(_01832_),
    .A2_N(_01737_),
    .B1(_01817_),
    .B2(_01821_),
    .Y(_01833_));
 sky130_fd_sc_hd__o211ai_4 _30222_ (.A1(_01823_),
    .A2(_01829_),
    .B1(_01830_),
    .C1(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__a21bo_1 _30223_ (.A1(_01832_),
    .A2(_01736_),
    .B1_N(_01822_),
    .X(_01835_));
 sky130_fd_sc_hd__o211ai_2 _30224_ (.A1(_01817_),
    .A2(_01821_),
    .B1(_01832_),
    .C1(_01737_),
    .Y(_01836_));
 sky130_fd_sc_hd__o2bb2a_1 _30225_ (.A1_N(_00184_),
    .A2_N(_00169_),
    .B1(_00182_),
    .B2(_00180_),
    .X(_01837_));
 sky130_fd_sc_hd__nand3_4 _30226_ (.A(_01835_),
    .B(_01836_),
    .C(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__a21oi_1 _30227_ (.A1(_22648_),
    .A2(_22651_),
    .B1(_24047_),
    .Y(_01839_));
 sky130_fd_sc_hd__a32o_1 _30228_ (.A1(_01839_),
    .A2(_00200_),
    .A3(_00202_),
    .B1(_00206_),
    .B2(_00209_),
    .X(_01840_));
 sky130_fd_sc_hd__clkbuf_2 _30229_ (.A(\delay_line[2][11] ),
    .X(_01841_));
 sky130_fd_sc_hd__or2b_1 _30230_ (.A(\delay_line[3][10] ),
    .B_N(\delay_line[2][12] ),
    .X(_01843_));
 sky130_fd_sc_hd__or2b_1 _30231_ (.A(\delay_line[2][12] ),
    .B_N(\delay_line[3][10] ),
    .X(_01844_));
 sky130_fd_sc_hd__a22o_1 _30232_ (.A1(_19044_),
    .A2(_00207_),
    .B1(_01843_),
    .B2(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__nand4_2 _30233_ (.A(_19044_),
    .B(_01843_),
    .C(_01844_),
    .D(_00207_),
    .Y(_01846_));
 sky130_fd_sc_hd__a22o_1 _30234_ (.A1(_01841_),
    .A2(_22640_),
    .B1(_01845_),
    .B2(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__o21a_1 _30235_ (.A1(_21958_),
    .A2(_00208_),
    .B1(_24040_),
    .X(_01848_));
 sky130_fd_sc_hd__nand4_2 _30236_ (.A(_22640_),
    .B(_01845_),
    .C(_01841_),
    .D(_01846_),
    .Y(_01849_));
 sky130_fd_sc_hd__and3_1 _30237_ (.A(_01847_),
    .B(_01848_),
    .C(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__a21oi_1 _30238_ (.A1(_01849_),
    .A2(_01847_),
    .B1(_01848_),
    .Y(_01851_));
 sky130_fd_sc_hd__o21ai_1 _30239_ (.A1(_01850_),
    .A2(_01851_),
    .B1(_00234_),
    .Y(_01852_));
 sky130_fd_sc_hd__or3_1 _30240_ (.A(_01851_),
    .B(_00234_),
    .C(_01850_),
    .X(_01854_));
 sky130_fd_sc_hd__and3_1 _30241_ (.A(_01840_),
    .B(_01852_),
    .C(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__a21oi_1 _30242_ (.A1(_01852_),
    .A2(_01854_),
    .B1(_01840_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _30243_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__or2b_1 _30244_ (.A(_00235_),
    .B_N(_00239_),
    .X(_01858_));
 sky130_fd_sc_hd__xnor2_1 _30245_ (.A(_01857_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__or2b_1 _30246_ (.A(_19882_),
    .B_N(\delay_line[3][12] ),
    .X(_01860_));
 sky130_fd_sc_hd__buf_1 _30247_ (.A(\delay_line[3][12] ),
    .X(_01861_));
 sky130_fd_sc_hd__or2b_1 _30248_ (.A(_01861_),
    .B_N(_19883_),
    .X(_01862_));
 sky130_fd_sc_hd__buf_1 _30249_ (.A(\delay_line[5][10] ),
    .X(_01863_));
 sky130_fd_sc_hd__buf_2 _30250_ (.A(_01863_),
    .X(_01865_));
 sky130_fd_sc_hd__a21o_1 _30251_ (.A1(_01860_),
    .A2(_01862_),
    .B1(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__nand3_2 _30252_ (.A(_01860_),
    .B(_01862_),
    .C(_01865_),
    .Y(_01867_));
 sky130_fd_sc_hd__a32o_1 _30253_ (.A1(_00199_),
    .A2(_22627_),
    .A3(_00201_),
    .B1(_01865_),
    .B2(_09228_),
    .X(_01868_));
 sky130_fd_sc_hd__clkbuf_2 _30254_ (.A(\delay_line[5][12] ),
    .X(_01869_));
 sky130_fd_sc_hd__or2b_1 _30255_ (.A(_01869_),
    .B_N(_18082_),
    .X(_01870_));
 sky130_fd_sc_hd__or2b_2 _30256_ (.A(_18080_),
    .B_N(\delay_line[5][12] ),
    .X(_01871_));
 sky130_fd_sc_hd__clkbuf_2 _30257_ (.A(\delay_line[5][11] ),
    .X(_01872_));
 sky130_fd_sc_hd__nand3_2 _30258_ (.A(_01870_),
    .B(_01871_),
    .C(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__a21o_1 _30259_ (.A1(_01870_),
    .A2(_01871_),
    .B1(_01872_),
    .X(_01874_));
 sky130_fd_sc_hd__nand2_2 _30260_ (.A(_01873_),
    .B(_01874_),
    .Y(_01876_));
 sky130_fd_sc_hd__nand3_1 _30261_ (.A(_00196_),
    .B(_00201_),
    .C(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__a21o_1 _30262_ (.A1(_00196_),
    .A2(_00201_),
    .B1(_01876_),
    .X(_01878_));
 sky130_fd_sc_hd__a22o_1 _30263_ (.A1(_00200_),
    .A2(_01868_),
    .B1(_01877_),
    .B2(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__nand4_2 _30264_ (.A(_00200_),
    .B(_01868_),
    .C(_01877_),
    .D(_01878_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand4_2 _30265_ (.A(_01866_),
    .B(_01867_),
    .C(_01879_),
    .D(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__a22o_1 _30266_ (.A1(_01866_),
    .A2(_01867_),
    .B1(_01879_),
    .B2(_01880_),
    .X(_01882_));
 sky130_fd_sc_hd__a21oi_2 _30267_ (.A1(_24088_),
    .A2(_24096_),
    .B1(_00217_),
    .Y(_01883_));
 sky130_fd_sc_hd__clkbuf_2 _30268_ (.A(_24084_),
    .X(_01884_));
 sky130_fd_sc_hd__clkbuf_2 _30269_ (.A(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__o211ai_2 _30270_ (.A1(_00211_),
    .A2(_01885_),
    .B1(_24059_),
    .C1(_00213_),
    .Y(_01887_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30271_ (.A(_24062_),
    .X(_01888_));
 sky130_fd_sc_hd__nor3_1 _30272_ (.A(_00211_),
    .B(_01885_),
    .C(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__o21a_1 _30273_ (.A1(_00211_),
    .A2(_01884_),
    .B1(_01888_),
    .X(_01890_));
 sky130_fd_sc_hd__nand4_1 _30274_ (.A(_03238_),
    .B(_00256_),
    .C(_11976_),
    .D(_00257_),
    .Y(_01891_));
 sky130_fd_sc_hd__o211a_1 _30275_ (.A1(_01889_),
    .A2(_01890_),
    .B1(_00257_),
    .C1(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__a211oi_2 _30276_ (.A1(_00257_),
    .A2(_01891_),
    .B1(_01889_),
    .C1(_01890_),
    .Y(_01893_));
 sky130_fd_sc_hd__a211o_1 _30277_ (.A1(_00212_),
    .A2(_01887_),
    .B1(_01892_),
    .C1(_01893_),
    .X(_01894_));
 sky130_fd_sc_hd__o211ai_2 _30278_ (.A1(_01892_),
    .A2(_01893_),
    .B1(_00212_),
    .C1(_01887_),
    .Y(_01895_));
 sky130_fd_sc_hd__o211ai_4 _30279_ (.A1(_01883_),
    .A2(_00220_),
    .B1(_01894_),
    .C1(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__a221o_1 _30280_ (.A1(_24066_),
    .A2(_00219_),
    .B1(_01894_),
    .B2(_01895_),
    .C1(_01883_),
    .X(_01898_));
 sky130_fd_sc_hd__nand4_2 _30281_ (.A(_01881_),
    .B(_01882_),
    .C(_01896_),
    .D(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__a22o_1 _30282_ (.A1(_01881_),
    .A2(_01882_),
    .B1(_01896_),
    .B2(_01898_),
    .X(_01900_));
 sky130_fd_sc_hd__o21bai_1 _30283_ (.A1(_00210_),
    .A2(_00223_),
    .B1_N(_00222_),
    .Y(_01901_));
 sky130_fd_sc_hd__a21o_1 _30284_ (.A1(_01899_),
    .A2(_01900_),
    .B1(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__nand3_1 _30285_ (.A(_01901_),
    .B(_01899_),
    .C(_01900_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_1 _30286_ (.A(_01902_),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__xnor2_1 _30287_ (.A(_01859_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__nor2_1 _30288_ (.A(_00279_),
    .B(_00284_),
    .Y(_01906_));
 sky130_fd_sc_hd__inv_2 _30289_ (.A(_00278_),
    .Y(_01907_));
 sky130_fd_sc_hd__clkbuf_2 _30290_ (.A(_00268_),
    .X(_01909_));
 sky130_fd_sc_hd__nand4_1 _30291_ (.A(_00264_),
    .B(_00267_),
    .C(_01909_),
    .D(_24093_),
    .Y(_01910_));
 sky130_fd_sc_hd__nand2_1 _30292_ (.A(_01910_),
    .B(_00272_),
    .Y(_01911_));
 sky130_fd_sc_hd__buf_1 _30293_ (.A(_00261_),
    .X(_01912_));
 sky130_fd_sc_hd__or2_1 _30294_ (.A(_01912_),
    .B(_22527_),
    .X(_01913_));
 sky130_fd_sc_hd__nand2_1 _30295_ (.A(_00265_),
    .B(_21862_),
    .Y(_01914_));
 sky130_fd_sc_hd__buf_1 _30296_ (.A(_00253_),
    .X(_01915_));
 sky130_fd_sc_hd__a21o_1 _30297_ (.A1(_01913_),
    .A2(_01914_),
    .B1(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__nand3_1 _30298_ (.A(_01913_),
    .B(_01914_),
    .C(_01915_),
    .Y(_01917_));
 sky130_fd_sc_hd__o21ai_1 _30299_ (.A1(_24092_),
    .A2(_00265_),
    .B1(_00252_),
    .Y(_01918_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30300_ (.A(\delay_line[6][12] ),
    .X(_01920_));
 sky130_fd_sc_hd__nand2_1 _30301_ (.A(_11976_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__or2_1 _30302_ (.A(_11965_),
    .B(\delay_line[6][12] ),
    .X(_01922_));
 sky130_fd_sc_hd__a22o_1 _30303_ (.A1(_00266_),
    .A2(_01918_),
    .B1(_01921_),
    .B2(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30304_ (.A(net427),
    .X(_01924_));
 sky130_fd_sc_hd__nand4_1 _30305_ (.A(_00266_),
    .B(_01918_),
    .C(_01921_),
    .D(_01922_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand4_2 _30306_ (.A(_22591_),
    .B(_01923_),
    .C(_01924_),
    .D(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__a22o_1 _30307_ (.A1(net427),
    .A2(_22591_),
    .B1(_01923_),
    .B2(_01925_),
    .X(_01927_));
 sky130_fd_sc_hd__and4_1 _30308_ (.A(_01916_),
    .B(_01917_),
    .C(_01926_),
    .D(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__inv_2 _30309_ (.A(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__a22o_1 _30310_ (.A1(_01916_),
    .A2(_01917_),
    .B1(_01926_),
    .B2(_01927_),
    .X(_01931_));
 sky130_fd_sc_hd__nand2_1 _30311_ (.A(_01929_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__a21oi_1 _30312_ (.A1(_23933_),
    .A2(_25306_),
    .B1(_25304_),
    .Y(_01933_));
 sky130_fd_sc_hd__xnor2_1 _30313_ (.A(_01932_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__xnor2_1 _30314_ (.A(_01911_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__o21ai_1 _30315_ (.A1(_25327_),
    .A2(_25330_),
    .B1(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__or3_1 _30316_ (.A(_25327_),
    .B(_25330_),
    .C(_01935_),
    .X(_01937_));
 sky130_fd_sc_hd__o211a_2 _30317_ (.A1(_00275_),
    .A2(_01907_),
    .B1(_01936_),
    .C1(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__a211oi_2 _30318_ (.A1(_01936_),
    .A2(_01937_),
    .B1(_00275_),
    .C1(_01907_),
    .Y(_01939_));
 sky130_fd_sc_hd__or3_2 _30319_ (.A(_01906_),
    .B(_01938_),
    .C(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__o21ai_1 _30320_ (.A1(_01938_),
    .A2(_01939_),
    .B1(_01906_),
    .Y(_01942_));
 sky130_fd_sc_hd__nand3b_1 _30321_ (.A_N(_01905_),
    .B(_01940_),
    .C(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__a21bo_1 _30322_ (.A1(_01940_),
    .A2(_01942_),
    .B1_N(_01905_),
    .X(_01944_));
 sky130_fd_sc_hd__o21ai_4 _30323_ (.A1(_25364_),
    .A2(_25360_),
    .B1(_25361_),
    .Y(_01945_));
 sky130_fd_sc_hd__a21o_1 _30324_ (.A1(_01943_),
    .A2(_01944_),
    .B1(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__nand3_2 _30325_ (.A(_01945_),
    .B(_01943_),
    .C(_01944_),
    .Y(_01947_));
 sky130_fd_sc_hd__and2b_1 _30326_ (.A_N(_00248_),
    .B(_00286_),
    .X(_01948_));
 sky130_fd_sc_hd__or2_1 _30327_ (.A(net136),
    .B(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__a21oi_2 _30328_ (.A1(_01946_),
    .A2(_01947_),
    .B1(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__and3_1 _30329_ (.A(_01949_),
    .B(_01946_),
    .C(_01947_),
    .X(_01951_));
 sky130_fd_sc_hd__o2bb2ai_4 _30330_ (.A1_N(_01834_),
    .A2_N(_01838_),
    .B1(_01950_),
    .B2(_01951_),
    .Y(_01953_));
 sky130_fd_sc_hd__nor2_1 _30331_ (.A(_01950_),
    .B(_01951_),
    .Y(_01954_));
 sky130_fd_sc_hd__nand3_4 _30332_ (.A(_01834_),
    .B(_01838_),
    .C(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__o22a_1 _30333_ (.A1(_00297_),
    .A2(_00298_),
    .B1(_00177_),
    .B2(_00186_),
    .X(_01956_));
 sky130_fd_sc_hd__o2bb2ai_1 _30334_ (.A1_N(_01953_),
    .A2_N(_01955_),
    .B1(_01956_),
    .B2(_00306_),
    .Y(_01957_));
 sky130_fd_sc_hd__o2111ai_4 _30335_ (.A1(_00294_),
    .A2(_00187_),
    .B1(_00300_),
    .C1(_01953_),
    .D1(_01955_),
    .Y(_01958_));
 sky130_fd_sc_hd__nand2_1 _30336_ (.A(_01957_),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__a2bb2oi_1 _30337_ (.A1_N(_01480_),
    .A2_N(_01482_),
    .B1(_01524_),
    .B2(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__nand3b_2 _30338_ (.A_N(_01524_),
    .B(_01957_),
    .C(_01958_),
    .Y(_01961_));
 sky130_fd_sc_hd__clkbuf_2 _30339_ (.A(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__nor2_1 _30340_ (.A(_00310_),
    .B(_00355_),
    .Y(_01964_));
 sky130_fd_sc_hd__or2_1 _30341_ (.A(_01964_),
    .B(_00360_),
    .X(_01965_));
 sky130_fd_sc_hd__nand2_1 _30342_ (.A(_01521_),
    .B(_01518_),
    .Y(_01966_));
 sky130_fd_sc_hd__and4b_2 _30343_ (.A_N(_01966_),
    .B(_00351_),
    .C(_00350_),
    .D(_00352_),
    .X(_01967_));
 sky130_fd_sc_hd__a21oi_2 _30344_ (.A1(_00292_),
    .A2(_00363_),
    .B1(_00191_),
    .Y(_01968_));
 sky130_fd_sc_hd__a21oi_4 _30345_ (.A1(_01953_),
    .A2(_01955_),
    .B1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__o211a_2 _30346_ (.A1(_01823_),
    .A2(_01829_),
    .B1(_01830_),
    .C1(_01833_),
    .X(_01970_));
 sky130_fd_sc_hd__nand2_1 _30347_ (.A(_01838_),
    .B(_01954_),
    .Y(_01971_));
 sky130_fd_sc_hd__o211a_2 _30348_ (.A1(_01970_),
    .A2(_01971_),
    .B1(_01968_),
    .C1(_01953_),
    .X(_01972_));
 sky130_fd_sc_hd__o22ai_4 _30349_ (.A1(_01522_),
    .A2(_01967_),
    .B1(_01969_),
    .B2(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__a2bb2o_1 _30350_ (.A1_N(_00364_),
    .A2_N(_00365_),
    .B1(_00361_),
    .B2(_00303_),
    .X(_01975_));
 sky130_fd_sc_hd__a21oi_2 _30351_ (.A1(_01973_),
    .A2(_01961_),
    .B1(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__a211o_1 _30352_ (.A1(_01960_),
    .A2(_01962_),
    .B1(_01965_),
    .C1(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__o211a_1 _30353_ (.A1(_01480_),
    .A2(_01482_),
    .B1(_01973_),
    .C1(_01961_),
    .X(_01978_));
 sky130_fd_sc_hd__o22ai_1 _30354_ (.A1(_01964_),
    .A2(_00360_),
    .B1(_01976_),
    .B2(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__o22a_1 _30355_ (.A1(_00368_),
    .A2(_00362_),
    .B1(_00377_),
    .B2(_00373_),
    .X(_01980_));
 sky130_fd_sc_hd__nand3_1 _30356_ (.A(_01977_),
    .B(_01979_),
    .C(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__o22a_2 _30357_ (.A1(_01522_),
    .A2(_01967_),
    .B1(_01969_),
    .B2(_01972_),
    .X(_01982_));
 sky130_fd_sc_hd__o21ai_2 _30358_ (.A1(_01480_),
    .A2(_01482_),
    .B1(_01962_),
    .Y(_01983_));
 sky130_fd_sc_hd__a21o_1 _30359_ (.A1(_01973_),
    .A2(_01962_),
    .B1(_01975_),
    .X(_01984_));
 sky130_fd_sc_hd__o221ai_4 _30360_ (.A1(_01964_),
    .A2(_00360_),
    .B1(_01982_),
    .B2(_01983_),
    .C1(_01984_),
    .Y(_01986_));
 sky130_fd_sc_hd__inv_2 _30361_ (.A(_01965_),
    .Y(_01987_));
 sky130_fd_sc_hd__o21ai_2 _30362_ (.A1(_01976_),
    .A2(_01978_),
    .B1(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hd__nand3b_4 _30363_ (.A_N(_01980_),
    .B(_01986_),
    .C(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_2 _30364_ (.A(_01981_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__o21ai_1 _30365_ (.A1(_22729_),
    .A2(_23745_),
    .B1(_23746_),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _30366_ (.A(_00406_),
    .B(_00407_),
    .Y(_01992_));
 sky130_fd_sc_hd__nand4b_1 _30367_ (.A_N(_24214_),
    .B(_01991_),
    .C(_00387_),
    .D(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__o2bb2ai_1 _30368_ (.A1_N(_00406_),
    .A2_N(_00407_),
    .B1(_24217_),
    .B2(_24207_),
    .Y(_01994_));
 sky130_fd_sc_hd__o21ai_1 _30369_ (.A1(_00402_),
    .A2(_00404_),
    .B1(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__nand3_2 _30370_ (.A(_01990_),
    .B(_01993_),
    .C(_01995_),
    .Y(_01997_));
 sky130_fd_sc_hd__o21ai_1 _30371_ (.A1(_24231_),
    .A2(_24232_),
    .B1(_00408_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand4_2 _30372_ (.A(_00387_),
    .B(_01998_),
    .C(_01981_),
    .D(_01989_),
    .Y(_01999_));
 sky130_fd_sc_hd__buf_2 _30373_ (.A(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__nand2_1 _30374_ (.A(_01997_),
    .B(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__clkbuf_2 _30375_ (.A(\delay_line[23][11] ),
    .X(_02002_));
 sky130_fd_sc_hd__nor2_1 _30376_ (.A(_02002_),
    .B(net347),
    .Y(_02003_));
 sky130_fd_sc_hd__and2_2 _30377_ (.A(_02002_),
    .B(net347),
    .X(_02004_));
 sky130_fd_sc_hd__nor2_1 _30378_ (.A(_02003_),
    .B(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _30379_ (.A(_02001_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__a32o_2 _30380_ (.A1(_01228_),
    .A2(_01229_),
    .A3(_01251_),
    .B1(_01252_),
    .B2(_01265_),
    .X(_02008_));
 sky130_fd_sc_hd__inv_2 _30381_ (.A(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__o211ai_1 _30382_ (.A1(_02003_),
    .A2(_02004_),
    .B1(_01997_),
    .C1(_02000_),
    .Y(_02010_));
 sky130_fd_sc_hd__and3_2 _30383_ (.A(_02006_),
    .B(_02009_),
    .C(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__o21ai_1 _30384_ (.A1(_02003_),
    .A2(_02004_),
    .B1(_02001_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand3_1 _30385_ (.A(_01997_),
    .B(_02000_),
    .C(_02005_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand3_2 _30386_ (.A(_02008_),
    .B(_02012_),
    .C(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__clkbuf_2 _30387_ (.A(_24225_),
    .X(_02015_));
 sky130_fd_sc_hd__clkbuf_2 _30388_ (.A(_02002_),
    .X(_02016_));
 sky130_fd_sc_hd__clkbuf_2 _30389_ (.A(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__buf_2 _30390_ (.A(_24225_),
    .X(_02019_));
 sky130_fd_sc_hd__o211a_1 _30391_ (.A1(_02019_),
    .A2(_02002_),
    .B1(_00390_),
    .C1(_00393_),
    .X(_02020_));
 sky130_fd_sc_hd__a21oi_1 _30392_ (.A1(_02015_),
    .A2(_02017_),
    .B1(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__nand2_1 _30393_ (.A(_02014_),
    .B(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__o31a_1 _30394_ (.A1(_01266_),
    .A2(_01267_),
    .A3(_01319_),
    .B1(_01320_),
    .X(_02023_));
 sky130_fd_sc_hd__nand3_1 _30395_ (.A(_02006_),
    .B(_02009_),
    .C(_02010_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _30396_ (.A(_02024_),
    .B(_02014_),
    .Y(_02025_));
 sky130_fd_sc_hd__o21ai_1 _30397_ (.A1(_00399_),
    .A2(_02020_),
    .B1(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__o211ai_4 _30398_ (.A1(_02011_),
    .A2(_02022_),
    .B1(_02023_),
    .C1(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__o21ai_1 _30399_ (.A1(_00399_),
    .A2(_02020_),
    .B1(_02014_),
    .Y(_02028_));
 sky130_fd_sc_hd__o21ai_2 _30400_ (.A1(_01319_),
    .A2(_01268_),
    .B1(_01320_),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2_1 _30401_ (.A(_02025_),
    .B(_02021_),
    .Y(_02031_));
 sky130_fd_sc_hd__o211ai_4 _30402_ (.A1(_02028_),
    .A2(_02011_),
    .B1(_02030_),
    .C1(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__nand2_1 _30403_ (.A(_00411_),
    .B(_00422_),
    .Y(_02033_));
 sky130_fd_sc_hd__a21oi_2 _30404_ (.A1(_02027_),
    .A2(_02032_),
    .B1(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__o211a_1 _30405_ (.A1(_25293_),
    .A2(_25061_),
    .B1(_00398_),
    .C1(_00410_),
    .X(_02035_));
 sky130_fd_sc_hd__o211a_1 _30406_ (.A1(_02035_),
    .A2(_00419_),
    .B1(_02027_),
    .C1(_02032_),
    .X(_02036_));
 sky130_fd_sc_hd__nor3_4 _30407_ (.A(_01478_),
    .B(_02034_),
    .C(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30408_ (.A(_04601_),
    .X(_02038_));
 sky130_fd_sc_hd__nor2_1 _30409_ (.A(_22781_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__a21oi_1 _30410_ (.A1(_02038_),
    .A2(_10372_),
    .B1(_02039_),
    .Y(_02041_));
 sky130_fd_sc_hd__and2_1 _30411_ (.A(_22111_),
    .B(net348),
    .X(_02042_));
 sky130_fd_sc_hd__nor2_1 _30412_ (.A(_22111_),
    .B(net348),
    .Y(_02043_));
 sky130_fd_sc_hd__and4bb_1 _30413_ (.A_N(_02042_),
    .B_N(_02043_),
    .C(_22109_),
    .D(_22749_),
    .X(_02044_));
 sky130_fd_sc_hd__o2bb2a_1 _30414_ (.A1_N(_22109_),
    .A2_N(_22749_),
    .B1(_02042_),
    .B2(_02043_),
    .X(_02045_));
 sky130_fd_sc_hd__or2_1 _30415_ (.A(_02044_),
    .B(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__nor2_1 _30416_ (.A(_02041_),
    .B(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__o21a_1 _30417_ (.A1(_02044_),
    .A2(_02045_),
    .B1(_02041_),
    .X(_02048_));
 sky130_fd_sc_hd__o21ai_2 _30418_ (.A1(_02034_),
    .A2(_02036_),
    .B1(_01478_),
    .Y(_02049_));
 sky130_fd_sc_hd__o21ai_2 _30419_ (.A1(_02047_),
    .A2(_02048_),
    .B1(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__a21o_1 _30420_ (.A1(_02027_),
    .A2(_02032_),
    .B1(_02033_),
    .X(_02052_));
 sky130_fd_sc_hd__o211ai_2 _30421_ (.A1(_02035_),
    .A2(_00419_),
    .B1(_02027_),
    .C1(_02032_),
    .Y(_02053_));
 sky130_fd_sc_hd__a21o_1 _30422_ (.A1(_00424_),
    .A2(_00428_),
    .B1(_00420_),
    .X(_02054_));
 sky130_fd_sc_hd__a21oi_1 _30423_ (.A1(_02052_),
    .A2(_02053_),
    .B1(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__nor2_1 _30424_ (.A(_02047_),
    .B(_02048_),
    .Y(_02056_));
 sky130_fd_sc_hd__o21ai_2 _30425_ (.A1(_02055_),
    .A2(_02037_),
    .B1(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__o221ai_2 _30426_ (.A1(_01476_),
    .A2(_01477_),
    .B1(_02037_),
    .B2(_02050_),
    .C1(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__nand3_1 _30427_ (.A(_02054_),
    .B(_02052_),
    .C(_02053_),
    .Y(_02059_));
 sky130_fd_sc_hd__a21o_1 _30428_ (.A1(_02049_),
    .A2(_02059_),
    .B1(_02056_),
    .X(_02060_));
 sky130_fd_sc_hd__nand3_1 _30429_ (.A(_02049_),
    .B(_02059_),
    .C(_02056_),
    .Y(_02061_));
 sky130_fd_sc_hd__o21ai_2 _30430_ (.A1(_01066_),
    .A2(_01327_),
    .B1(_01324_),
    .Y(_02063_));
 sky130_fd_sc_hd__inv_2 _30431_ (.A(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__nand3_1 _30432_ (.A(_02060_),
    .B(_02061_),
    .C(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__and3_2 _30433_ (.A(_01475_),
    .B(_02058_),
    .C(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__a21o_1 _30434_ (.A1(_02058_),
    .A2(_02065_),
    .B1(_01475_),
    .X(_02067_));
 sky130_fd_sc_hd__inv_2 _30435_ (.A(_01064_),
    .Y(_02068_));
 sky130_fd_sc_hd__or2b_1 _30436_ (.A(_01065_),
    .B_N(_01330_),
    .X(_02069_));
 sky130_fd_sc_hd__o21ai_2 _30437_ (.A1(_00463_),
    .A2(_02068_),
    .B1(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__a21bo_1 _30438_ (.A1(_00879_),
    .A2(_01063_),
    .B1_N(_00880_),
    .X(_02071_));
 sky130_fd_sc_hd__and2b_2 _30439_ (.A_N(_00964_),
    .B(_01056_),
    .X(_02072_));
 sky130_fd_sc_hd__or2b_1 _30440_ (.A(_20332_),
    .B_N(net321),
    .X(_02074_));
 sky130_fd_sc_hd__or4b_2 _30441_ (.A(_19323_),
    .B(_00917_),
    .C(_00918_),
    .D_N(net322),
    .X(_02075_));
 sky130_fd_sc_hd__and2b_1 _30442_ (.A_N(_21300_),
    .B(\delay_line[29][10] ),
    .X(_02076_));
 sky130_fd_sc_hd__and2b_1 _30443_ (.A_N(\delay_line[29][10] ),
    .B(_21300_),
    .X(_02077_));
 sky130_fd_sc_hd__nor2_1 _30444_ (.A(_02076_),
    .B(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__a21oi_1 _30445_ (.A1(_02074_),
    .A2(_02075_),
    .B1(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__and3_1 _30446_ (.A(_02074_),
    .B(_02075_),
    .C(_02078_),
    .X(_02080_));
 sky130_fd_sc_hd__a41o_1 _30447_ (.A1(_18451_),
    .A2(_00915_),
    .A3(_24433_),
    .A4(_00920_),
    .B1(_00925_),
    .X(_02081_));
 sky130_fd_sc_hd__or3_1 _30448_ (.A(_02079_),
    .B(_02080_),
    .C(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__o21ai_2 _30449_ (.A1(_02079_),
    .A2(_02080_),
    .B1(_02081_),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _30450_ (.A(_02082_),
    .B(_02083_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand2_2 _30451_ (.A(_00953_),
    .B(_00927_),
    .Y(_02086_));
 sky130_fd_sc_hd__a221oi_2 _30452_ (.A1(_24399_),
    .A2(_24398_),
    .B1(_00946_),
    .B2(_00948_),
    .C1(_00931_),
    .Y(_02087_));
 sky130_fd_sc_hd__o21ai_4 _30453_ (.A1(_00928_),
    .A2(_02087_),
    .B1(_00949_),
    .Y(_02088_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30454_ (.A(_00940_),
    .X(_02089_));
 sky130_fd_sc_hd__and3_1 _30455_ (.A(_06337_),
    .B(_18453_),
    .C(_02089_),
    .X(_02090_));
 sky130_fd_sc_hd__a31oi_4 _30456_ (.A1(_00943_),
    .A2(_00942_),
    .A3(_20346_),
    .B1(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__clkbuf_2 _30457_ (.A(_00934_),
    .X(_02092_));
 sky130_fd_sc_hd__o211a_1 _30458_ (.A1(_20350_),
    .A2(_23246_),
    .B1(_23251_),
    .C1(_23252_),
    .X(_02093_));
 sky130_fd_sc_hd__a2111oi_4 _30459_ (.A1(_15569_),
    .A2(_02092_),
    .B1(_23268_),
    .C1(_06315_),
    .D1(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__and3_1 _30460_ (.A(_15569_),
    .B(_19336_),
    .C(_23269_),
    .X(_02096_));
 sky130_fd_sc_hd__o22a_1 _30461_ (.A1(_23268_),
    .A2(_06326_),
    .B1(_02096_),
    .B2(_02093_),
    .X(_02097_));
 sky130_fd_sc_hd__nor2_1 _30462_ (.A(_02094_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__clkbuf_2 _30463_ (.A(\delay_line[30][11] ),
    .X(_02099_));
 sky130_fd_sc_hd__nor2_1 _30464_ (.A(_00933_),
    .B(_02092_),
    .Y(_02100_));
 sky130_fd_sc_hd__inv_2 _30465_ (.A(\delay_line[30][12] ),
    .Y(_02101_));
 sky130_fd_sc_hd__clkbuf_2 _30466_ (.A(_23248_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_1 _30467_ (.A(_00940_),
    .B(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__and2_1 _30468_ (.A(_20348_),
    .B(_23248_),
    .X(_02104_));
 sky130_fd_sc_hd__or3_2 _30469_ (.A(_02101_),
    .B(_02103_),
    .C(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__clkbuf_2 _30470_ (.A(_02104_),
    .X(_02107_));
 sky130_fd_sc_hd__o21ai_2 _30471_ (.A1(_02103_),
    .A2(_02107_),
    .B1(_02101_),
    .Y(_02108_));
 sky130_fd_sc_hd__a22o_1 _30472_ (.A1(_02099_),
    .A2(_02100_),
    .B1(_02105_),
    .B2(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__clkbuf_2 _30473_ (.A(_02099_),
    .X(_02110_));
 sky130_fd_sc_hd__nand4_4 _30474_ (.A(_02105_),
    .B(_02108_),
    .C(_02110_),
    .D(_02100_),
    .Y(_02111_));
 sky130_fd_sc_hd__nand3_2 _30475_ (.A(_02098_),
    .B(_02109_),
    .C(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__o2bb2ai_1 _30476_ (.A1_N(_02111_),
    .A2_N(_02109_),
    .B1(_02094_),
    .B2(_02097_),
    .Y(_02113_));
 sky130_fd_sc_hd__nor3_1 _30477_ (.A(_00937_),
    .B(_00938_),
    .C(_00947_),
    .Y(_02114_));
 sky130_fd_sc_hd__a211oi_1 _30478_ (.A1(_02112_),
    .A2(_02113_),
    .B1(_00937_),
    .C1(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__o211a_1 _30479_ (.A1(_00937_),
    .A2(_02114_),
    .B1(_02112_),
    .C1(_02113_),
    .X(_02116_));
 sky130_fd_sc_hd__nor2_2 _30480_ (.A(_02115_),
    .B(_02116_),
    .Y(_02118_));
 sky130_fd_sc_hd__xnor2_4 _30481_ (.A(_02091_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__xor2_4 _30482_ (.A(_02088_),
    .B(_02119_),
    .X(_02120_));
 sky130_fd_sc_hd__xnor2_4 _30483_ (.A(_02086_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__a31oi_2 _30484_ (.A1(_23280_),
    .A2(_24393_),
    .A3(_24426_),
    .B1(_24423_),
    .Y(_02122_));
 sky130_fd_sc_hd__o2bb2ai_4 _30485_ (.A1_N(_00926_),
    .A2_N(_00955_),
    .B1(_00954_),
    .B2(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__xor2_2 _30486_ (.A(_02121_),
    .B(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__xor2_1 _30487_ (.A(_02085_),
    .B(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__or2_2 _30488_ (.A(_24472_),
    .B(_00911_),
    .X(_02126_));
 sky130_fd_sc_hd__buf_1 _30489_ (.A(\delay_line[31][12] ),
    .X(_02127_));
 sky130_fd_sc_hd__nor2_1 _30490_ (.A(net316),
    .B(_02127_),
    .Y(_02129_));
 sky130_fd_sc_hd__nand2_1 _30491_ (.A(_00885_),
    .B(_02127_),
    .Y(_02130_));
 sky130_fd_sc_hd__nand3b_1 _30492_ (.A_N(_02129_),
    .B(_02130_),
    .C(_00884_),
    .Y(_02131_));
 sky130_fd_sc_hd__and2_1 _30493_ (.A(\delay_line[31][11] ),
    .B(_02127_),
    .X(_02132_));
 sky130_fd_sc_hd__o21bai_2 _30494_ (.A1(_02129_),
    .A2(_02132_),
    .B1_N(_00884_),
    .Y(_02133_));
 sky130_fd_sc_hd__o21ai_1 _30495_ (.A1(_23207_),
    .A2(_00883_),
    .B1(_00886_),
    .Y(_02134_));
 sky130_fd_sc_hd__and3_1 _30496_ (.A(_02131_),
    .B(_02133_),
    .C(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30497_ (.A(_02131_),
    .X(_02136_));
 sky130_fd_sc_hd__a21o_1 _30498_ (.A1(_02136_),
    .A2(_02133_),
    .B1(_02134_),
    .X(_02137_));
 sky130_fd_sc_hd__nand3b_1 _30499_ (.A_N(_02135_),
    .B(_02137_),
    .C(_00896_),
    .Y(_02138_));
 sky130_fd_sc_hd__a21oi_1 _30500_ (.A1(_02136_),
    .A2(_02133_),
    .B1(_02134_),
    .Y(_02140_));
 sky130_fd_sc_hd__o21ai_1 _30501_ (.A1(_02135_),
    .A2(_02140_),
    .B1(_00894_),
    .Y(_02141_));
 sky130_fd_sc_hd__or2_1 _30502_ (.A(_21270_),
    .B(_24447_),
    .X(_02142_));
 sky130_fd_sc_hd__buf_1 _30503_ (.A(_20307_),
    .X(_02143_));
 sky130_fd_sc_hd__buf_1 _30504_ (.A(_21270_),
    .X(_02144_));
 sky130_fd_sc_hd__nand2_1 _30505_ (.A(_24447_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__nand4_1 _30506_ (.A(_06271_),
    .B(_02142_),
    .C(_02143_),
    .D(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__a22o_1 _30507_ (.A1(_02143_),
    .A2(_06271_),
    .B1(_02142_),
    .B2(_02145_),
    .X(_02147_));
 sky130_fd_sc_hd__a22o_1 _30508_ (.A1(_02138_),
    .A2(_02141_),
    .B1(_02146_),
    .B2(_02147_),
    .X(_02148_));
 sky130_fd_sc_hd__nand4_1 _30509_ (.A(_02138_),
    .B(_02141_),
    .C(_02146_),
    .D(_02147_),
    .Y(_02149_));
 sky130_fd_sc_hd__nand2_1 _30510_ (.A(_00895_),
    .B(_00905_),
    .Y(_02151_));
 sky130_fd_sc_hd__nand3_1 _30511_ (.A(_02148_),
    .B(_02149_),
    .C(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__a21o_1 _30512_ (.A1(_02148_),
    .A2(_02149_),
    .B1(_02151_),
    .X(_02153_));
 sky130_fd_sc_hd__nand2_1 _30513_ (.A(_02152_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__xor2_1 _30514_ (.A(_00901_),
    .B(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__o211ai_1 _30515_ (.A1(_24449_),
    .A2(_00908_),
    .B1(_02155_),
    .C1(_00906_),
    .Y(_02156_));
 sky130_fd_sc_hd__a21o_1 _30516_ (.A1(_00906_),
    .A2(_00909_),
    .B1(_02155_),
    .X(_02157_));
 sky130_fd_sc_hd__nand2_2 _30517_ (.A(_02156_),
    .B(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__xnor2_4 _30518_ (.A(_02126_),
    .B(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _30519_ (.A(_23221_),
    .B(_24473_),
    .Y(_02160_));
 sky130_fd_sc_hd__inv_2 _30520_ (.A(_00911_),
    .Y(_02162_));
 sky130_fd_sc_hd__a22oi_4 _30521_ (.A1(_02160_),
    .A2(_02162_),
    .B1(_00913_),
    .B2(_00912_),
    .Y(_02163_));
 sky130_fd_sc_hd__xnor2_2 _30522_ (.A(_02159_),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_2 _30523_ (.A(_02125_),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__and2_1 _30524_ (.A(_02125_),
    .B(_02164_),
    .X(_02166_));
 sky130_fd_sc_hd__nor2_2 _30525_ (.A(_02165_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__o21bai_1 _30526_ (.A1(_01047_),
    .A2(_01048_),
    .B1_N(_01045_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _30527_ (.A(_01036_),
    .B(_19304_),
    .Y(_02169_));
 sky130_fd_sc_hd__a21oi_1 _30528_ (.A1(_01028_),
    .A2(_01032_),
    .B1(net325),
    .Y(_02170_));
 sky130_fd_sc_hd__and3_1 _30529_ (.A(_24311_),
    .B(net326),
    .C(net325),
    .X(_02171_));
 sky130_fd_sc_hd__buf_1 _30530_ (.A(_20407_),
    .X(_02173_));
 sky130_fd_sc_hd__o21ba_1 _30531_ (.A1(_02170_),
    .A2(_02171_),
    .B1_N(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__nor3b_1 _30532_ (.A(_02170_),
    .B(_02171_),
    .C_N(_02173_),
    .Y(_02175_));
 sky130_fd_sc_hd__a211oi_2 _30533_ (.A1(_01034_),
    .A2(_02169_),
    .B1(_02174_),
    .C1(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__o211a_1 _30534_ (.A1(_02174_),
    .A2(_02175_),
    .B1(_01034_),
    .C1(_02169_),
    .X(_02177_));
 sky130_fd_sc_hd__nor3_1 _30535_ (.A(_02176_),
    .B(_19301_),
    .C(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__o21a_1 _30536_ (.A1(_02177_),
    .A2(_02176_),
    .B1(_19301_),
    .X(_02179_));
 sky130_fd_sc_hd__nor2_1 _30537_ (.A(_02178_),
    .B(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__or3_1 _30538_ (.A(_01038_),
    .B(_01041_),
    .C(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__o21ai_1 _30539_ (.A1(_01038_),
    .A2(_01041_),
    .B1(_02180_),
    .Y(_02182_));
 sky130_fd_sc_hd__a21oi_1 _30540_ (.A1(_02181_),
    .A2(_02182_),
    .B1(_01043_),
    .Y(_02184_));
 sky130_fd_sc_hd__and3_1 _30541_ (.A(_02181_),
    .B(_02182_),
    .C(_01043_),
    .X(_02185_));
 sky130_fd_sc_hd__nor2_1 _30542_ (.A(_02184_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__xnor2_1 _30543_ (.A(_02168_),
    .B(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__nor2_1 _30544_ (.A(_01004_),
    .B(_01006_),
    .Y(_02188_));
 sky130_fd_sc_hd__or4b_1 _30545_ (.A(_23132_),
    .B(_24350_),
    .C(_24351_),
    .D_N(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__o211ai_2 _30546_ (.A1(_24340_),
    .A2(_00997_),
    .B1(_01001_),
    .C1(_01003_),
    .Y(_02190_));
 sky130_fd_sc_hd__buf_1 _30547_ (.A(\delay_line[26][7] ),
    .X(_02191_));
 sky130_fd_sc_hd__nor2_1 _30548_ (.A(_00998_),
    .B(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__nand2_1 _30549_ (.A(_20397_),
    .B(_21228_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand3b_1 _30550_ (.A_N(_02192_),
    .B(_02193_),
    .C(_16020_),
    .Y(_02195_));
 sky130_fd_sc_hd__and2_1 _30551_ (.A(_00998_),
    .B(_02191_),
    .X(_02196_));
 sky130_fd_sc_hd__o21ai_1 _30552_ (.A1(_02192_),
    .A2(_02196_),
    .B1(_21223_),
    .Y(_02197_));
 sky130_fd_sc_hd__o21ai_1 _30553_ (.A1(_06480_),
    .A2(_00999_),
    .B1(_01000_),
    .Y(_02198_));
 sky130_fd_sc_hd__and3_1 _30554_ (.A(_02195_),
    .B(_02197_),
    .C(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__a21oi_1 _30555_ (.A1(_02195_),
    .A2(_02197_),
    .B1(_02198_),
    .Y(_02200_));
 sky130_fd_sc_hd__nor2_1 _30556_ (.A(_02199_),
    .B(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__o211a_1 _30557_ (.A1(_24344_),
    .A2(_01006_),
    .B1(_02190_),
    .C1(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__buf_1 _30558_ (.A(_02199_),
    .X(_02203_));
 sky130_fd_sc_hd__a32o_1 _30559_ (.A1(_01001_),
    .A2(_01003_),
    .A3(_01005_),
    .B1(_02188_),
    .B2(_24350_),
    .X(_02204_));
 sky130_fd_sc_hd__o21a_1 _30560_ (.A1(_02203_),
    .A2(_02200_),
    .B1(_02204_),
    .X(_02206_));
 sky130_fd_sc_hd__buf_1 _30561_ (.A(\delay_line[26][11] ),
    .X(_02207_));
 sky130_fd_sc_hd__o21a_1 _30562_ (.A1(_02202_),
    .A2(_02206_),
    .B1(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__nor3_1 _30563_ (.A(_02207_),
    .B(_02202_),
    .C(_02206_),
    .Y(_02209_));
 sky130_fd_sc_hd__a211oi_1 _30564_ (.A1(_01012_),
    .A2(_02189_),
    .B1(_02208_),
    .C1(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__o211a_1 _30565_ (.A1(_02208_),
    .A2(_02209_),
    .B1(_01012_),
    .C1(_02189_),
    .X(_02211_));
 sky130_fd_sc_hd__o211a_1 _30566_ (.A1(_02210_),
    .A2(_02211_),
    .B1(_01015_),
    .C1(_01020_),
    .X(_02212_));
 sky130_fd_sc_hd__a211oi_1 _30567_ (.A1(_01015_),
    .A2(_01020_),
    .B1(_02210_),
    .C1(_02211_),
    .Y(_02213_));
 sky130_fd_sc_hd__buf_1 _30568_ (.A(_00967_),
    .X(_02214_));
 sky130_fd_sc_hd__nor2_1 _30569_ (.A(_24360_),
    .B(\delay_line[27][12] ),
    .Y(_02215_));
 sky130_fd_sc_hd__buf_1 _30570_ (.A(\delay_line[27][12] ),
    .X(_02217_));
 sky130_fd_sc_hd__nand2_1 _30571_ (.A(_24366_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nand3b_1 _30572_ (.A_N(_02215_),
    .B(_02218_),
    .C(_00968_),
    .Y(_02219_));
 sky130_fd_sc_hd__and2_2 _30573_ (.A(_24360_),
    .B(\delay_line[27][12] ),
    .X(_02220_));
 sky130_fd_sc_hd__o21ai_2 _30574_ (.A1(_02215_),
    .A2(_02220_),
    .B1(_00966_),
    .Y(_02221_));
 sky130_fd_sc_hd__nand2_1 _30575_ (.A(_02219_),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__clkbuf_2 _30576_ (.A(\delay_line[27][12] ),
    .X(_02223_));
 sky130_fd_sc_hd__nor2_1 _30577_ (.A(_02223_),
    .B(_00967_),
    .Y(_02224_));
 sky130_fd_sc_hd__nand2_1 _30578_ (.A(_19277_),
    .B(_19280_),
    .Y(_02225_));
 sky130_fd_sc_hd__a211oi_1 _30579_ (.A1(_02214_),
    .A2(_02222_),
    .B1(_02224_),
    .C1(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__nor3_1 _30580_ (.A(_00965_),
    .B(_24361_),
    .C(_00968_),
    .Y(_02228_));
 sky130_fd_sc_hd__a21oi_1 _30581_ (.A1(_02219_),
    .A2(_02221_),
    .B1(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__o22a_1 _30582_ (.A1(net274),
    .A2(_19286_),
    .B1(_02229_),
    .B2(_02224_),
    .X(_02230_));
 sky130_fd_sc_hd__a22oi_1 _30583_ (.A1(_23155_),
    .A2(_00972_),
    .B1(_00967_),
    .B2(_00969_),
    .Y(_02231_));
 sky130_fd_sc_hd__o22ai_2 _30584_ (.A1(_00971_),
    .A2(_24362_),
    .B1(_18499_),
    .B2(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__o21bai_1 _30585_ (.A1(_02226_),
    .A2(_02230_),
    .B1_N(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__a211o_1 _30586_ (.A1(_02214_),
    .A2(_02222_),
    .B1(_02224_),
    .C1(_02225_),
    .X(_02234_));
 sky130_fd_sc_hd__o21ai_1 _30587_ (.A1(_02229_),
    .A2(_02224_),
    .B1(_02225_),
    .Y(_02235_));
 sky130_fd_sc_hd__nand3_2 _30588_ (.A(_02232_),
    .B(_02234_),
    .C(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand3b_1 _30589_ (.A_N(_18494_),
    .B(_02233_),
    .C(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__a2bb2o_1 _30590_ (.A1_N(_18496_),
    .A2_N(_19274_),
    .B1(_02233_),
    .B2(_02236_),
    .X(_02239_));
 sky130_fd_sc_hd__nand2_1 _30591_ (.A(_02237_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand2_1 _30592_ (.A(_00980_),
    .B(_00981_),
    .Y(_02241_));
 sky130_fd_sc_hd__xor2_1 _30593_ (.A(_02240_),
    .B(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__xnor2_1 _30594_ (.A(_00986_),
    .B(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__inv_2 _30595_ (.A(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__or3_1 _30596_ (.A(net135),
    .B(_00992_),
    .C(_02244_),
    .X(_02245_));
 sky130_fd_sc_hd__o21ai_1 _30597_ (.A1(net135),
    .A2(_00992_),
    .B1(_02244_),
    .Y(_02246_));
 sky130_fd_sc_hd__nand2_1 _30598_ (.A(_02245_),
    .B(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__or3_1 _30599_ (.A(_02212_),
    .B(_02213_),
    .C(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__a2bb2o_1 _30600_ (.A1_N(_02212_),
    .A2_N(_02213_),
    .B1(_02245_),
    .B2(_02246_),
    .X(_02250_));
 sky130_fd_sc_hd__nand2_1 _30601_ (.A(_02248_),
    .B(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__or2_1 _30602_ (.A(_02187_),
    .B(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__nand2_1 _30603_ (.A(_02251_),
    .B(_02187_),
    .Y(_02253_));
 sky130_fd_sc_hd__nand2_1 _30604_ (.A(_02252_),
    .B(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__o311a_1 _30605_ (.A1(_01022_),
    .A2(net107),
    .A3(_00993_),
    .B1(_01052_),
    .C1(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__a21oi_2 _30606_ (.A1(_01024_),
    .A2(_01052_),
    .B1(_02254_),
    .Y(_02256_));
 sky130_fd_sc_hd__nor2_2 _30607_ (.A(_02255_),
    .B(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__xor2_4 _30608_ (.A(_02167_),
    .B(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__or3_1 _30609_ (.A(_00594_),
    .B(net92),
    .C(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__o21ai_2 _30610_ (.A1(_00594_),
    .A2(net92),
    .B1(_02258_),
    .Y(_02261_));
 sky130_fd_sc_hd__nand2_1 _30611_ (.A(_02259_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__o21bai_4 _30612_ (.A1(_01055_),
    .A2(_02072_),
    .B1_N(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__or3b_1 _30613_ (.A(_01055_),
    .B(_02072_),
    .C_N(_02262_),
    .X(_02264_));
 sky130_fd_sc_hd__nand2_1 _30614_ (.A(_02263_),
    .B(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__o21bai_2 _30615_ (.A1(_00599_),
    .A2(_00873_),
    .B1_N(_00875_),
    .Y(_02266_));
 sky130_fd_sc_hd__o21a_1 _30616_ (.A1(_00509_),
    .A2(_00589_),
    .B1(_00587_),
    .X(_02267_));
 sky130_fd_sc_hd__a32o_1 _30617_ (.A1(_24529_),
    .A2(_24531_),
    .A3(_24532_),
    .B1(_00501_),
    .B2(_00503_),
    .X(_02268_));
 sky130_fd_sc_hd__a21oi_2 _30618_ (.A1(_00464_),
    .A2(_02268_),
    .B1(_00507_),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_1 _30619_ (.A(_00500_),
    .B(_00503_),
    .Y(_02270_));
 sky130_fd_sc_hd__or3b_1 _30620_ (.A(_06821_),
    .B(_00465_),
    .C_N(_24499_),
    .X(_02272_));
 sky130_fd_sc_hd__and2b_1 _30621_ (.A_N(_22822_),
    .B(_18324_),
    .X(_02273_));
 sky130_fd_sc_hd__o21a_1 _30622_ (.A1(_18325_),
    .A2(_18326_),
    .B1(_22822_),
    .X(_02274_));
 sky130_fd_sc_hd__buf_1 _30623_ (.A(\delay_line[25][12] ),
    .X(_02275_));
 sky130_fd_sc_hd__nor2_1 _30624_ (.A(_24511_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__and2_1 _30625_ (.A(_24505_),
    .B(\delay_line[25][12] ),
    .X(_02277_));
 sky130_fd_sc_hd__o21bai_1 _30626_ (.A1(_02276_),
    .A2(_02277_),
    .B1_N(_00473_),
    .Y(_02278_));
 sky130_fd_sc_hd__nand2_1 _30627_ (.A(_24511_),
    .B(_02275_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand3b_1 _30628_ (.A_N(_02276_),
    .B(_02279_),
    .C(_00473_),
    .Y(_02280_));
 sky130_fd_sc_hd__nand3_1 _30629_ (.A(_02278_),
    .B(_21565_),
    .C(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__a21o_1 _30630_ (.A1(_02280_),
    .A2(_02278_),
    .B1(_21565_),
    .X(_02283_));
 sky130_fd_sc_hd__a2bb2o_1 _30631_ (.A1_N(_00473_),
    .A2_N(_00475_),
    .B1(_21569_),
    .B2(_00477_),
    .X(_02284_));
 sky130_fd_sc_hd__nand3_1 _30632_ (.A(_02281_),
    .B(_02283_),
    .C(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__a21o_1 _30633_ (.A1(_02281_),
    .A2(_02283_),
    .B1(_02284_),
    .X(_02286_));
 sky130_fd_sc_hd__o211a_1 _30634_ (.A1(_02273_),
    .A2(_02274_),
    .B1(_02285_),
    .C1(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__or2_1 _30635_ (.A(_02273_),
    .B(_02274_),
    .X(_02288_));
 sky130_fd_sc_hd__a21oi_1 _30636_ (.A1(_02285_),
    .A2(_02286_),
    .B1(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__a21boi_1 _30637_ (.A1(_00488_),
    .A2(_00486_),
    .B1_N(_00483_),
    .Y(_02290_));
 sky130_fd_sc_hd__o21ai_2 _30638_ (.A1(_02287_),
    .A2(_02289_),
    .B1(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__o211ai_1 _30639_ (.A1(_02273_),
    .A2(_02274_),
    .B1(_02285_),
    .C1(_02286_),
    .Y(_02292_));
 sky130_fd_sc_hd__a21o_1 _30640_ (.A1(_02285_),
    .A2(_02286_),
    .B1(_02288_),
    .X(_02294_));
 sky130_fd_sc_hd__nand3b_1 _30641_ (.A_N(_02290_),
    .B(_02292_),
    .C(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__clkbuf_2 _30642_ (.A(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__nand2_1 _30643_ (.A(_00470_),
    .B(_06799_),
    .Y(_02297_));
 sky130_fd_sc_hd__a21o_1 _30644_ (.A1(_02291_),
    .A2(_02296_),
    .B1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__nand3_1 _30645_ (.A(_02297_),
    .B(_02291_),
    .C(_02296_),
    .Y(_02299_));
 sky130_fd_sc_hd__nand4_1 _30646_ (.A(_00490_),
    .B(_00495_),
    .C(_02298_),
    .D(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__a21boi_1 _30647_ (.A1(_00494_),
    .A2(_00496_),
    .B1_N(_00490_),
    .Y(_02301_));
 sky130_fd_sc_hd__nand4_2 _30648_ (.A(_02291_),
    .B(_00465_),
    .C(_17237_),
    .D(_02296_),
    .Y(_02302_));
 sky130_fd_sc_hd__a22o_1 _30649_ (.A1(_00465_),
    .A2(_17237_),
    .B1(_02291_),
    .B2(_02295_),
    .X(_02303_));
 sky130_fd_sc_hd__nand3b_2 _30650_ (.A_N(_02301_),
    .B(_02302_),
    .C(_02303_),
    .Y(_02305_));
 sky130_fd_sc_hd__nand3_1 _30651_ (.A(_02272_),
    .B(_02300_),
    .C(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__a21o_1 _30652_ (.A1(_02300_),
    .A2(_02305_),
    .B1(_02272_),
    .X(_02307_));
 sky130_fd_sc_hd__nand2_1 _30653_ (.A(_02306_),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__xnor2_2 _30654_ (.A(_02270_),
    .B(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__xor2_2 _30655_ (.A(_02269_),
    .B(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__a21boi_1 _30656_ (.A1(_00578_),
    .A2(_24596_),
    .B1_N(_00580_),
    .Y(_02311_));
 sky130_fd_sc_hd__a21boi_1 _30657_ (.A1(_00572_),
    .A2(_00573_),
    .B1_N(_00574_),
    .Y(_02312_));
 sky130_fd_sc_hd__o21a_1 _30658_ (.A1(_19519_),
    .A2(_00549_),
    .B1(_00550_),
    .X(_02313_));
 sky130_fd_sc_hd__and2_1 _30659_ (.A(_00548_),
    .B(net342),
    .X(_02314_));
 sky130_fd_sc_hd__o21ai_2 _30660_ (.A1(_00548_),
    .A2(_22883_),
    .B1(_20463_),
    .Y(_02316_));
 sky130_fd_sc_hd__clkbuf_2 _30661_ (.A(\delay_line[24][11] ),
    .X(_02317_));
 sky130_fd_sc_hd__nor2_1 _30662_ (.A(_00548_),
    .B(net342),
    .Y(_02318_));
 sky130_fd_sc_hd__o21ai_2 _30663_ (.A1(_02314_),
    .A2(_02318_),
    .B1(_20467_),
    .Y(_02319_));
 sky130_fd_sc_hd__o211a_1 _30664_ (.A1(_02314_),
    .A2(_02316_),
    .B1(_02317_),
    .C1(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__a21o_1 _30665_ (.A1(_21619_),
    .A2(_22883_),
    .B1(_02316_),
    .X(_02321_));
 sky130_fd_sc_hd__clkbuf_2 _30666_ (.A(_02317_),
    .X(_02322_));
 sky130_fd_sc_hd__a21oi_1 _30667_ (.A1(_02321_),
    .A2(_02319_),
    .B1(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__o21ai_1 _30668_ (.A1(_02320_),
    .A2(_02323_),
    .B1(_00554_),
    .Y(_02324_));
 sky130_fd_sc_hd__o211ai_1 _30669_ (.A1(_02314_),
    .A2(_02316_),
    .B1(_02322_),
    .C1(_02319_),
    .Y(_02325_));
 sky130_fd_sc_hd__a21o_1 _30670_ (.A1(_02321_),
    .A2(_02319_),
    .B1(_02317_),
    .X(_02327_));
 sky130_fd_sc_hd__nand3_1 _30671_ (.A(_00561_),
    .B(_02325_),
    .C(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__nand3b_1 _30672_ (.A_N(_02313_),
    .B(_02324_),
    .C(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand3_1 _30673_ (.A(_02327_),
    .B(_00554_),
    .C(_02325_),
    .Y(_02330_));
 sky130_fd_sc_hd__o21ai_1 _30674_ (.A1(_02320_),
    .A2(_02323_),
    .B1(_00561_),
    .Y(_02331_));
 sky130_fd_sc_hd__o2111ai_2 _30675_ (.A1(_19519_),
    .A2(_00549_),
    .B1(_00550_),
    .C1(_02330_),
    .D1(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__o21a_1 _30676_ (.A1(_00554_),
    .A2(_00556_),
    .B1(_24581_),
    .X(_02333_));
 sky130_fd_sc_hd__o21ai_1 _30677_ (.A1(_00547_),
    .A2(_02333_),
    .B1(_00567_),
    .Y(_02334_));
 sky130_fd_sc_hd__a21o_1 _30678_ (.A1(_02329_),
    .A2(_02332_),
    .B1(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30679_ (.A(_22877_),
    .X(_02336_));
 sky130_fd_sc_hd__nand2_1 _30680_ (.A(_02336_),
    .B(_22871_),
    .Y(_02338_));
 sky130_fd_sc_hd__and3_1 _30681_ (.A(_02338_),
    .B(_18310_),
    .C(_06909_),
    .X(_02339_));
 sky130_fd_sc_hd__a21oi_1 _30682_ (.A1(_02338_),
    .A2(_18310_),
    .B1(_06920_),
    .Y(_02340_));
 sky130_fd_sc_hd__nor2_1 _30683_ (.A(_02339_),
    .B(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__nand3_1 _30684_ (.A(_02334_),
    .B(_02329_),
    .C(_02332_),
    .Y(_02342_));
 sky130_fd_sc_hd__nand3_1 _30685_ (.A(_02335_),
    .B(_02341_),
    .C(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__nand2_1 _30686_ (.A(_02342_),
    .B(_02335_),
    .Y(_02344_));
 sky130_fd_sc_hd__o21ai_1 _30687_ (.A1(_02339_),
    .A2(_02340_),
    .B1(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand3b_2 _30688_ (.A_N(_02312_),
    .B(_02343_),
    .C(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__nand2_1 _30689_ (.A(_02344_),
    .B(_02341_),
    .Y(_02347_));
 sky130_fd_sc_hd__o211ai_1 _30690_ (.A1(_02339_),
    .A2(_02340_),
    .B1(_02342_),
    .C1(_02335_),
    .Y(_02349_));
 sky130_fd_sc_hd__nand3_1 _30691_ (.A(_02347_),
    .B(_02349_),
    .C(_02312_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand4_1 _30692_ (.A(_02346_),
    .B(_01457_),
    .C(_02350_),
    .D(_22878_),
    .Y(_02351_));
 sky130_fd_sc_hd__nand2_1 _30693_ (.A(_02350_),
    .B(_02346_),
    .Y(_02352_));
 sky130_fd_sc_hd__o21ai_1 _30694_ (.A1(_19508_),
    .A2(_24572_),
    .B1(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__nand2_1 _30695_ (.A(_02351_),
    .B(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _30696_ (.A(_02311_),
    .B(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__nand2_1 _30697_ (.A(_02354_),
    .B(_02311_),
    .Y(_02356_));
 sky130_fd_sc_hd__or2b_1 _30698_ (.A(_02355_),
    .B_N(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__xnor2_2 _30699_ (.A(_00586_),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__clkbuf_2 _30700_ (.A(\delay_line[22][3] ),
    .X(_02360_));
 sky130_fd_sc_hd__nand2_1 _30701_ (.A(_01413_),
    .B(_06865_),
    .Y(_02361_));
 sky130_fd_sc_hd__o21ai_1 _30702_ (.A1(_00527_),
    .A2(_00523_),
    .B1(_00529_),
    .Y(_02362_));
 sky130_fd_sc_hd__buf_1 _30703_ (.A(\delay_line[22][7] ),
    .X(_02363_));
 sky130_fd_sc_hd__nor2_1 _30704_ (.A(_02363_),
    .B(\delay_line[22][11] ),
    .Y(_02364_));
 sky130_fd_sc_hd__nand2_1 _30705_ (.A(_02363_),
    .B(\delay_line[22][11] ),
    .Y(_02365_));
 sky130_fd_sc_hd__nand3b_1 _30706_ (.A_N(_02364_),
    .B(_00521_),
    .C(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__inv_2 _30707_ (.A(\delay_line[22][10] ),
    .Y(_02367_));
 sky130_fd_sc_hd__and2_1 _30708_ (.A(net352),
    .B(\delay_line[22][11] ),
    .X(_02368_));
 sky130_fd_sc_hd__o22ai_2 _30709_ (.A1(_21599_),
    .A2(_02367_),
    .B1(_02368_),
    .B2(_02364_),
    .Y(_02369_));
 sky130_fd_sc_hd__inv_2 _30710_ (.A(\delay_line[22][4] ),
    .Y(_02371_));
 sky130_fd_sc_hd__or3_1 _30711_ (.A(_21600_),
    .B(_02371_),
    .C(_17073_),
    .X(_02372_));
 sky130_fd_sc_hd__o21ai_1 _30712_ (.A1(_21600_),
    .A2(_17084_),
    .B1(_02371_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand4_2 _30713_ (.A(_02366_),
    .B(_02369_),
    .C(_02372_),
    .D(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__a22o_1 _30714_ (.A1(_02366_),
    .A2(_02369_),
    .B1(_02372_),
    .B2(_02373_),
    .X(_02375_));
 sky130_fd_sc_hd__nand3_2 _30715_ (.A(_02362_),
    .B(_02374_),
    .C(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21o_1 _30716_ (.A1(_02374_),
    .A2(_02375_),
    .B1(_02362_),
    .X(_02377_));
 sky130_fd_sc_hd__o2111ai_4 _30717_ (.A1(_02360_),
    .A2(_02361_),
    .B1(_02376_),
    .C1(_06876_),
    .D1(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__a22o_1 _30718_ (.A1(_00525_),
    .A2(_06876_),
    .B1(_02377_),
    .B2(_02376_),
    .X(_02379_));
 sky130_fd_sc_hd__and3_1 _30719_ (.A(_00528_),
    .B(_00531_),
    .C(_00533_),
    .X(_02380_));
 sky130_fd_sc_hd__a31oi_1 _30720_ (.A1(_00534_),
    .A2(_01413_),
    .A3(_24554_),
    .B1(_02380_),
    .Y(_02382_));
 sky130_fd_sc_hd__a21bo_1 _30721_ (.A1(_02378_),
    .A2(_02379_),
    .B1_N(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__nand3b_2 _30722_ (.A_N(_02382_),
    .B(_02378_),
    .C(_02379_),
    .Y(_02384_));
 sky130_fd_sc_hd__nand3b_2 _30723_ (.A_N(_24554_),
    .B(_02383_),
    .C(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__a2bb2o_1 _30724_ (.A1_N(_22852_),
    .A2_N(_06887_),
    .B1(_02384_),
    .B2(_02383_),
    .X(_02386_));
 sky130_fd_sc_hd__a21oi_1 _30725_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_00540_),
    .Y(_02387_));
 sky130_fd_sc_hd__nor4_1 _30726_ (.A(_24541_),
    .B(_24566_),
    .C(_00539_),
    .D(_00540_),
    .Y(_02388_));
 sky130_fd_sc_hd__a21oi_1 _30727_ (.A1(_00511_),
    .A2(_00542_),
    .B1(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__and3_1 _30728_ (.A(_02386_),
    .B(_00540_),
    .C(_02385_),
    .X(_02390_));
 sky130_fd_sc_hd__o21ai_1 _30729_ (.A1(_02390_),
    .A2(_02387_),
    .B1(_02389_),
    .Y(_02391_));
 sky130_fd_sc_hd__o21ai_2 _30730_ (.A1(_02387_),
    .A2(_02389_),
    .B1(_02391_),
    .Y(_02393_));
 sky130_fd_sc_hd__xor2_1 _30731_ (.A(_02358_),
    .B(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__nand2_1 _30732_ (.A(_02310_),
    .B(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__or2_1 _30733_ (.A(_02310_),
    .B(_02394_),
    .X(_02396_));
 sky130_fd_sc_hd__a21bo_2 _30734_ (.A1(_00649_),
    .A2(_00738_),
    .B1_N(_00737_),
    .X(_02397_));
 sky130_fd_sc_hd__a21oi_1 _30735_ (.A1(_02395_),
    .A2(_02396_),
    .B1(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__nand3_1 _30736_ (.A(_02397_),
    .B(_02395_),
    .C(_02396_),
    .Y(_02399_));
 sky130_fd_sc_hd__or3b_2 _30737_ (.A(_02267_),
    .B(_02398_),
    .C_N(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__or2b_1 _30738_ (.A(_02398_),
    .B_N(_02399_),
    .X(_02401_));
 sky130_fd_sc_hd__nand2_1 _30739_ (.A(_02401_),
    .B(_02267_),
    .Y(_02402_));
 sky130_fd_sc_hd__nand2_4 _30740_ (.A(_02400_),
    .B(_02402_),
    .Y(_02404_));
 sky130_fd_sc_hd__clkbuf_2 _30741_ (.A(_00749_),
    .X(_02405_));
 sky130_fd_sc_hd__nor2_1 _30742_ (.A(_00743_),
    .B(_00745_),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _30743_ (.A(\delay_line[14][6] ),
    .B(_21492_),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_1 _30744_ (.A(_20587_),
    .B(_21492_),
    .Y(_02408_));
 sky130_fd_sc_hd__nand3b_2 _30745_ (.A_N(_02407_),
    .B(_02408_),
    .C(\delay_line[14][11] ),
    .Y(_02409_));
 sky130_fd_sc_hd__and2_1 _30746_ (.A(_20587_),
    .B(_21497_),
    .X(_02410_));
 sky130_fd_sc_hd__o21bai_1 _30747_ (.A1(_02407_),
    .A2(_02410_),
    .B1_N(\delay_line[14][11] ),
    .Y(_02411_));
 sky130_fd_sc_hd__a22oi_2 _30748_ (.A1(_02405_),
    .A2(_02406_),
    .B1(_02409_),
    .B2(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__a21oi_1 _30749_ (.A1(_19452_),
    .A2(_20589_),
    .B1(_16832_),
    .Y(_02413_));
 sky130_fd_sc_hd__and3_1 _30750_ (.A(_16832_),
    .B(_19452_),
    .C(_20589_),
    .X(_02415_));
 sky130_fd_sc_hd__nor2_1 _30751_ (.A(_02413_),
    .B(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__nand4_1 _30752_ (.A(_02411_),
    .B(_02405_),
    .C(_02409_),
    .D(_02406_),
    .Y(_02417_));
 sky130_fd_sc_hd__nand3b_1 _30753_ (.A_N(_02412_),
    .B(_02416_),
    .C(_02417_),
    .Y(_02418_));
 sky130_fd_sc_hd__and4_1 _30754_ (.A(_02411_),
    .B(_00749_),
    .C(_02409_),
    .D(_02406_),
    .X(_02419_));
 sky130_fd_sc_hd__o22ai_1 _30755_ (.A1(_02413_),
    .A2(_02415_),
    .B1(_02419_),
    .B2(_02412_),
    .Y(_02420_));
 sky130_fd_sc_hd__a211o_1 _30756_ (.A1(_02418_),
    .A2(_02420_),
    .B1(_00751_),
    .C1(_00753_),
    .X(_02421_));
 sky130_fd_sc_hd__o211ai_1 _30757_ (.A1(_00751_),
    .A2(_00753_),
    .B1(_02418_),
    .C1(_02420_),
    .Y(_02422_));
 sky130_fd_sc_hd__nand2_1 _30758_ (.A(_02421_),
    .B(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__xnor2_2 _30759_ (.A(_00742_),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand2_1 _30760_ (.A(_00756_),
    .B(_00758_),
    .Y(_02426_));
 sky130_fd_sc_hd__xor2_2 _30761_ (.A(_02424_),
    .B(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__a311o_2 _30762_ (.A1(_00760_),
    .A2(_00758_),
    .A3(_00759_),
    .B1(_00764_),
    .C1(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__o21ai_2 _30763_ (.A1(_00762_),
    .A2(_00764_),
    .B1(_02427_),
    .Y(_02429_));
 sky130_fd_sc_hd__and2_1 _30764_ (.A(_24736_),
    .B(\delay_line[15][12] ),
    .X(_02430_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30765_ (.A(\delay_line[15][12] ),
    .X(_02431_));
 sky130_fd_sc_hd__o211ai_2 _30766_ (.A1(_24736_),
    .A2(_02431_),
    .B1(_00774_),
    .C1(_23078_),
    .Y(_02432_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30767_ (.A(_20599_),
    .X(_02433_));
 sky130_fd_sc_hd__inv_2 _30768_ (.A(\delay_line[15][11] ),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_1 _30769_ (.A(_24736_),
    .B(_02431_),
    .Y(_02435_));
 sky130_fd_sc_hd__o22ai_2 _30770_ (.A1(_24739_),
    .A2(_02434_),
    .B1(_02430_),
    .B2(_02435_),
    .Y(_02437_));
 sky130_fd_sc_hd__o211a_1 _30771_ (.A1(_02430_),
    .A2(_02432_),
    .B1(_02433_),
    .C1(_02437_),
    .X(_02438_));
 sky130_fd_sc_hd__a21o_1 _30772_ (.A1(_24737_),
    .A2(_02431_),
    .B1(_02432_),
    .X(_02439_));
 sky130_fd_sc_hd__a21o_1 _30773_ (.A1(_02439_),
    .A2(_02437_),
    .B1(_02433_),
    .X(_02440_));
 sky130_fd_sc_hd__o2bb2ai_1 _30774_ (.A1_N(_21458_),
    .A2_N(_00779_),
    .B1(_00776_),
    .B2(_00775_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand3b_2 _30775_ (.A_N(_02438_),
    .B(_02440_),
    .C(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__buf_1 _30776_ (.A(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__a21oi_1 _30777_ (.A1(_02439_),
    .A2(_02437_),
    .B1(_02433_),
    .Y(_02444_));
 sky130_fd_sc_hd__o21bai_4 _30778_ (.A1(_02438_),
    .A2(_02444_),
    .B1_N(_02441_),
    .Y(_02445_));
 sky130_fd_sc_hd__nor2_1 _30779_ (.A(_18412_),
    .B(_21454_),
    .Y(_02446_));
 sky130_fd_sc_hd__o21a_1 _30780_ (.A1(_18415_),
    .A2(_18418_),
    .B1(_18412_),
    .X(_02448_));
 sky130_fd_sc_hd__o2bb2ai_1 _30781_ (.A1_N(_02443_),
    .A2_N(_02445_),
    .B1(_02446_),
    .B2(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__o21a_1 _30782_ (.A1(_16788_),
    .A2(_18429_),
    .B1(_21454_),
    .X(_02450_));
 sky130_fd_sc_hd__and3b_1 _30783_ (.A_N(_16788_),
    .B(_18423_),
    .C(_18412_),
    .X(_02451_));
 sky130_fd_sc_hd__o211ai_1 _30784_ (.A1(_02450_),
    .A2(_02451_),
    .B1(_02443_),
    .C1(_02445_),
    .Y(_02452_));
 sky130_fd_sc_hd__nand4_2 _30785_ (.A(_00785_),
    .B(_00790_),
    .C(_02449_),
    .D(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__a211oi_1 _30786_ (.A1(_24746_),
    .A2(_24744_),
    .B1(_00780_),
    .C1(_00786_),
    .Y(_02454_));
 sky130_fd_sc_hd__a21o_1 _30787_ (.A1(_00791_),
    .A2(_00789_),
    .B1(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__o211ai_2 _30788_ (.A1(_02446_),
    .A2(_02448_),
    .B1(_02442_),
    .C1(_02445_),
    .Y(_02456_));
 sky130_fd_sc_hd__o2bb2ai_1 _30789_ (.A1_N(_02443_),
    .A2_N(_02445_),
    .B1(_02450_),
    .B2(_02451_),
    .Y(_02457_));
 sky130_fd_sc_hd__nand3_2 _30790_ (.A(_02455_),
    .B(_02456_),
    .C(_02457_),
    .Y(_02459_));
 sky130_fd_sc_hd__o21ai_1 _30791_ (.A1(_18413_),
    .A2(_00798_),
    .B1(_00769_),
    .Y(_02460_));
 sky130_fd_sc_hd__a21o_1 _30792_ (.A1(_02453_),
    .A2(_02459_),
    .B1(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__nand3_1 _30793_ (.A(_02460_),
    .B(_02453_),
    .C(_02459_),
    .Y(_02462_));
 sky130_fd_sc_hd__and4_1 _30794_ (.A(_00803_),
    .B(_00797_),
    .C(_02461_),
    .D(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__nand2_1 _30795_ (.A(_00803_),
    .B(_00797_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _30796_ (.A(_02453_),
    .B(_02459_),
    .Y(_02465_));
 sky130_fd_sc_hd__or2_1 _30797_ (.A(_02460_),
    .B(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__or3b_2 _30798_ (.A(_00798_),
    .B(_18412_),
    .C_N(_07107_),
    .X(_02467_));
 sky130_fd_sc_hd__a22o_1 _30799_ (.A1(_00769_),
    .A2(_02467_),
    .B1(_02453_),
    .B2(_02459_),
    .X(_02468_));
 sky130_fd_sc_hd__and3_1 _30800_ (.A(_02464_),
    .B(_02466_),
    .C(_02468_),
    .X(_02470_));
 sky130_fd_sc_hd__o32a_2 _30801_ (.A1(_24763_),
    .A2(_00798_),
    .A3(_00769_),
    .B1(_02463_),
    .B2(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__a22o_1 _30802_ (.A1(_00803_),
    .A2(_00797_),
    .B1(_02461_),
    .B2(_02462_),
    .X(_02472_));
 sky130_fd_sc_hd__and4b_1 _30803_ (.A_N(_02463_),
    .B(_02472_),
    .C(_01820_),
    .D(_07129_),
    .X(_02473_));
 sky130_fd_sc_hd__a21o_1 _30804_ (.A1(_00802_),
    .A2(_00809_),
    .B1(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__o211a_2 _30805_ (.A1(_02471_),
    .A2(_02473_),
    .B1(_00802_),
    .C1(_00809_),
    .X(_02475_));
 sky130_fd_sc_hd__o21ba_1 _30806_ (.A1(_02471_),
    .A2(_02474_),
    .B1_N(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__a311o_1 _30807_ (.A1(_24767_),
    .A2(_00811_),
    .A3(_00809_),
    .B1(_00815_),
    .C1(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__o21ai_1 _30808_ (.A1(_24775_),
    .A2(_24779_),
    .B1(_24771_),
    .Y(_02478_));
 sky130_fd_sc_hd__a22oi_4 _30809_ (.A1(_00812_),
    .A2(_00809_),
    .B1(_02478_),
    .B2(_00813_),
    .Y(_02479_));
 sky130_fd_sc_hd__or2_1 _30810_ (.A(_02479_),
    .B(_02475_),
    .X(_02481_));
 sky130_fd_sc_hd__a22o_1 _30811_ (.A1(_02428_),
    .A2(_02429_),
    .B1(_02477_),
    .B2(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__a21boi_1 _30812_ (.A1(_24836_),
    .A2(_00856_),
    .B1_N(_00860_),
    .Y(_02483_));
 sky130_fd_sc_hd__a21boi_1 _30813_ (.A1(_00848_),
    .A2(_00852_),
    .B1_N(_00846_),
    .Y(_02484_));
 sky130_fd_sc_hd__o21ai_1 _30814_ (.A1(_19435_),
    .A2(_00826_),
    .B1(_00837_),
    .Y(_02485_));
 sky130_fd_sc_hd__nor2_1 _30815_ (.A(net384),
    .B(\delay_line[16][8] ),
    .Y(_02486_));
 sky130_fd_sc_hd__and2_1 _30816_ (.A(net384),
    .B(net383),
    .X(_02487_));
 sky130_fd_sc_hd__o21bai_1 _30817_ (.A1(_02486_),
    .A2(_02487_),
    .B1_N(_24816_),
    .Y(_02488_));
 sky130_fd_sc_hd__clkbuf_2 _30818_ (.A(net381),
    .X(_02489_));
 sky130_fd_sc_hd__nand2_1 _30819_ (.A(net384),
    .B(net383),
    .Y(_02490_));
 sky130_fd_sc_hd__nand3b_1 _30820_ (.A_N(_02486_),
    .B(_02490_),
    .C(_24816_),
    .Y(_02492_));
 sky130_fd_sc_hd__nand3_1 _30821_ (.A(_02488_),
    .B(_02489_),
    .C(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__clkbuf_2 _30822_ (.A(net381),
    .X(_02494_));
 sky130_fd_sc_hd__a21o_1 _30823_ (.A1(_02492_),
    .A2(_02488_),
    .B1(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__a21o_1 _30824_ (.A1(_02493_),
    .A2(_02495_),
    .B1(_00838_),
    .X(_02496_));
 sky130_fd_sc_hd__inv_2 _30825_ (.A(\delay_line[16][10] ),
    .Y(_02497_));
 sky130_fd_sc_hd__buf_2 _30826_ (.A(_02497_),
    .X(_02498_));
 sky130_fd_sc_hd__o21ai_1 _30827_ (.A1(_00826_),
    .A2(_00837_),
    .B1(_00830_),
    .Y(_02499_));
 sky130_fd_sc_hd__buf_1 _30828_ (.A(_02493_),
    .X(_02500_));
 sky130_fd_sc_hd__o211ai_1 _30829_ (.A1(_02498_),
    .A2(_02499_),
    .B1(_02500_),
    .C1(_02495_),
    .Y(_02501_));
 sky130_fd_sc_hd__nand3_1 _30830_ (.A(_02485_),
    .B(_02496_),
    .C(_02501_),
    .Y(_02503_));
 sky130_fd_sc_hd__nand3_1 _30831_ (.A(_02495_),
    .B(_00831_),
    .C(_02493_),
    .Y(_02504_));
 sky130_fd_sc_hd__o2bb2ai_1 _30832_ (.A1_N(_02493_),
    .A2_N(_02495_),
    .B1(_02498_),
    .B2(_02499_),
    .Y(_02505_));
 sky130_fd_sc_hd__o2111ai_2 _30833_ (.A1(_19441_),
    .A2(_00826_),
    .B1(_00837_),
    .C1(_02504_),
    .D1(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__nand2_1 _30834_ (.A(_02503_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__a21boi_1 _30835_ (.A1(_00842_),
    .A2(_00824_),
    .B1_N(_00844_),
    .Y(_02508_));
 sky130_fd_sc_hd__nand2_1 _30836_ (.A(_02507_),
    .B(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__and3_1 _30837_ (.A(_24814_),
    .B(_24835_),
    .C(_21509_),
    .X(_02510_));
 sky130_fd_sc_hd__a21oi_1 _30838_ (.A1(_24814_),
    .A2(_24835_),
    .B1(_21536_),
    .Y(_02511_));
 sky130_fd_sc_hd__nor2_1 _30839_ (.A(_02510_),
    .B(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__nand2_1 _30840_ (.A(_00844_),
    .B(_00845_),
    .Y(_02514_));
 sky130_fd_sc_hd__nand3_1 _30841_ (.A(_02514_),
    .B(_02503_),
    .C(_02506_),
    .Y(_02515_));
 sky130_fd_sc_hd__nand3_1 _30842_ (.A(_02509_),
    .B(_02512_),
    .C(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__a2bb2o_1 _30843_ (.A1_N(_02510_),
    .A2_N(_02511_),
    .B1(_02515_),
    .B2(_02509_),
    .X(_02517_));
 sky130_fd_sc_hd__nand3b_1 _30844_ (.A_N(_02484_),
    .B(_02516_),
    .C(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__nand2_1 _30845_ (.A(_02515_),
    .B(_02509_),
    .Y(_02519_));
 sky130_fd_sc_hd__nand2_1 _30846_ (.A(_02519_),
    .B(_02512_),
    .Y(_02520_));
 sky130_fd_sc_hd__o211ai_1 _30847_ (.A1(_02510_),
    .A2(_02511_),
    .B1(_02515_),
    .C1(_02509_),
    .Y(_02521_));
 sky130_fd_sc_hd__nand4_1 _30848_ (.A(_00847_),
    .B(_00858_),
    .C(_02520_),
    .D(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__nand4_1 _30849_ (.A(_02518_),
    .B(_01886_),
    .C(_02522_),
    .D(_00850_),
    .Y(_02523_));
 sky130_fd_sc_hd__a22o_1 _30850_ (.A1(_01886_),
    .A2(_00850_),
    .B1(_02522_),
    .B2(_02518_),
    .X(_02525_));
 sky130_fd_sc_hd__nand2_1 _30851_ (.A(_02523_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__nor2_1 _30852_ (.A(_02483_),
    .B(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__buf_1 _30853_ (.A(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__nand2_1 _30854_ (.A(_02526_),
    .B(_02483_),
    .Y(_02529_));
 sky130_fd_sc_hd__or2b_1 _30855_ (.A(_02528_),
    .B_N(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__xor2_1 _30856_ (.A(_00864_),
    .B(_02530_),
    .X(_02531_));
 sky130_fd_sc_hd__o2111ai_4 _30857_ (.A1(_02479_),
    .A2(_02475_),
    .B1(_02477_),
    .C1(_02429_),
    .D1(_02428_),
    .Y(_02532_));
 sky130_fd_sc_hd__and3_1 _30858_ (.A(_02482_),
    .B(_02531_),
    .C(_02532_),
    .X(_02533_));
 sky130_fd_sc_hd__a21oi_1 _30859_ (.A1(_02532_),
    .A2(_02482_),
    .B1(_02531_),
    .Y(_02534_));
 sky130_fd_sc_hd__nor2_1 _30860_ (.A(_02533_),
    .B(_02534_),
    .Y(_02536_));
 sky130_fd_sc_hd__nor3_1 _30861_ (.A(net101),
    .B(_00867_),
    .C(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__o21a_4 _30862_ (.A1(net101),
    .A2(_00867_),
    .B1(_02536_),
    .X(_02538_));
 sky130_fd_sc_hd__nor2_2 _30863_ (.A(_02537_),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__nor2_1 _30864_ (.A(net358),
    .B(\delay_line[21][11] ),
    .Y(_02540_));
 sky130_fd_sc_hd__and2_1 _30865_ (.A(net358),
    .B(\delay_line[21][11] ),
    .X(_02541_));
 sky130_fd_sc_hd__nand2_1 _30866_ (.A(\delay_line[21][9] ),
    .B(net358),
    .Y(_02542_));
 sky130_fd_sc_hd__o21ai_1 _30867_ (.A1(_02540_),
    .A2(_02541_),
    .B1(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__or2_1 _30868_ (.A(\delay_line[21][11] ),
    .B(_02542_),
    .X(_02544_));
 sky130_fd_sc_hd__and3_1 _30869_ (.A(_02543_),
    .B(_02544_),
    .C(_20521_),
    .X(_02545_));
 sky130_fd_sc_hd__a21oi_2 _30870_ (.A1(_02543_),
    .A2(_02544_),
    .B1(_21423_),
    .Y(_02547_));
 sky130_fd_sc_hd__a211o_1 _30871_ (.A1(_00618_),
    .A2(_00620_),
    .B1(_02545_),
    .C1(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _30872_ (.A(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__clkbuf_2 _30873_ (.A(_00613_),
    .X(_02550_));
 sky130_fd_sc_hd__o221ai_4 _30874_ (.A1(_00616_),
    .A2(_02550_),
    .B1(_02547_),
    .B2(_02545_),
    .C1(_00621_),
    .Y(_02551_));
 sky130_fd_sc_hd__a21oi_1 _30875_ (.A1(_07305_),
    .A2(_18347_),
    .B1(_18346_),
    .Y(_02552_));
 sky130_fd_sc_hd__a21oi_1 _30876_ (.A1(_19420_),
    .A2(_19421_),
    .B1(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__and3_1 _30877_ (.A(_19420_),
    .B(_02552_),
    .C(_19421_),
    .X(_02554_));
 sky130_fd_sc_hd__or2_1 _30878_ (.A(_02553_),
    .B(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__a21oi_1 _30879_ (.A1(_02549_),
    .A2(_02551_),
    .B1(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__and3_1 _30880_ (.A(_02555_),
    .B(_02548_),
    .C(_02551_),
    .X(_02558_));
 sky130_fd_sc_hd__a32o_1 _30881_ (.A1(_00611_),
    .A2(_00619_),
    .A3(_00621_),
    .B1(_00624_),
    .B2(_00628_),
    .X(_02559_));
 sky130_fd_sc_hd__o21bai_2 _30882_ (.A1(_02556_),
    .A2(_02558_),
    .B1_N(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__nor2_1 _30883_ (.A(_02556_),
    .B(_02558_),
    .Y(_02561_));
 sky130_fd_sc_hd__nand2_1 _30884_ (.A(_02561_),
    .B(_02559_),
    .Y(_02562_));
 sky130_fd_sc_hd__a21o_1 _30885_ (.A1(_07569_),
    .A2(_18353_),
    .B1(_07591_),
    .X(_02563_));
 sky130_fd_sc_hd__o21a_1 _30886_ (.A1(_18359_),
    .A2(_00607_),
    .B1(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__a21oi_1 _30887_ (.A1(_02560_),
    .A2(_02562_),
    .B1(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__and3_1 _30888_ (.A(_02562_),
    .B(_02564_),
    .C(_02560_),
    .X(_02566_));
 sky130_fd_sc_hd__nand2_1 _30889_ (.A(_00631_),
    .B(_00635_),
    .Y(_02567_));
 sky130_fd_sc_hd__o21bai_1 _30890_ (.A1(_02565_),
    .A2(_02566_),
    .B1_N(_02567_),
    .Y(_02569_));
 sky130_fd_sc_hd__o2111ai_2 _30891_ (.A1(_18359_),
    .A2(_00607_),
    .B1(_02563_),
    .C1(_02560_),
    .D1(_02562_),
    .Y(_02570_));
 sky130_fd_sc_hd__nand3b_2 _30892_ (.A_N(_02565_),
    .B(_02570_),
    .C(_02567_),
    .Y(_02571_));
 sky130_fd_sc_hd__nand2_1 _30893_ (.A(_02569_),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__or2_1 _30894_ (.A(_16536_),
    .B(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__a32o_1 _30895_ (.A1(_16547_),
    .A2(_16525_),
    .A3(_16514_),
    .B1(_02569_),
    .B2(_02571_),
    .X(_02574_));
 sky130_fd_sc_hd__nand2_1 _30896_ (.A(_00638_),
    .B(_00640_),
    .Y(_02575_));
 sky130_fd_sc_hd__nand3_1 _30897_ (.A(_02573_),
    .B(_02574_),
    .C(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__a21o_1 _30898_ (.A1(_02573_),
    .A2(_02574_),
    .B1(_02575_),
    .X(_02577_));
 sky130_fd_sc_hd__nand2_1 _30899_ (.A(_00643_),
    .B(_00639_),
    .Y(_02578_));
 sky130_fd_sc_hd__o21ai_2 _30900_ (.A1(_00644_),
    .A2(_00648_),
    .B1(_02578_),
    .Y(_02580_));
 sky130_fd_sc_hd__a21oi_2 _30901_ (.A1(_02576_),
    .A2(_02577_),
    .B1(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__and3_1 _30902_ (.A(_02580_),
    .B(_02576_),
    .C(_02577_),
    .X(_02582_));
 sky130_fd_sc_hd__a22oi_2 _30903_ (.A1(_00693_),
    .A2(_00697_),
    .B1(_00703_),
    .B2(_00699_),
    .Y(_02583_));
 sky130_fd_sc_hd__o2bb2ai_1 _30904_ (.A1_N(_00660_),
    .A2_N(_00663_),
    .B1(_00655_),
    .B2(_00662_),
    .Y(_02584_));
 sky130_fd_sc_hd__clkbuf_2 _30905_ (.A(\delay_line[19][11] ),
    .X(_02585_));
 sky130_fd_sc_hd__buf_2 _30906_ (.A(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__nand2_2 _30907_ (.A(_24654_),
    .B(\delay_line[19][10] ),
    .Y(_02587_));
 sky130_fd_sc_hd__nor2_1 _30908_ (.A(_00658_),
    .B(_02585_),
    .Y(_02588_));
 sky130_fd_sc_hd__and2_1 _30909_ (.A(_00658_),
    .B(\delay_line[19][11] ),
    .X(_02589_));
 sky130_fd_sc_hd__o21ai_2 _30910_ (.A1(_02588_),
    .A2(_02589_),
    .B1(_02587_),
    .Y(_02591_));
 sky130_fd_sc_hd__o211ai_4 _30911_ (.A1(_02586_),
    .A2(_02587_),
    .B1(_20560_),
    .C1(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__or2_1 _30912_ (.A(_02585_),
    .B(_02587_),
    .X(_02593_));
 sky130_fd_sc_hd__a21o_1 _30913_ (.A1(_02591_),
    .A2(_02593_),
    .B1(_20560_),
    .X(_02594_));
 sky130_fd_sc_hd__nand3_2 _30914_ (.A(_02584_),
    .B(_02592_),
    .C(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__buf_1 _30915_ (.A(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__and3_2 _30916_ (.A(_02591_),
    .B(_02593_),
    .C(_20561_),
    .X(_02597_));
 sky130_fd_sc_hd__a21oi_1 _30917_ (.A1(_02591_),
    .A2(_02593_),
    .B1(_20561_),
    .Y(_02598_));
 sky130_fd_sc_hd__o21bai_4 _30918_ (.A1(_02597_),
    .A2(_02598_),
    .B1_N(_02584_),
    .Y(_02599_));
 sky130_fd_sc_hd__a21oi_1 _30919_ (.A1(_07382_),
    .A2(_18375_),
    .B1(_16404_),
    .Y(_02600_));
 sky130_fd_sc_hd__a21oi_2 _30920_ (.A1(_19404_),
    .A2(_19406_),
    .B1(_02600_),
    .Y(_02602_));
 sky130_fd_sc_hd__and3_1 _30921_ (.A(_19404_),
    .B(_19406_),
    .C(_02600_),
    .X(_02603_));
 sky130_fd_sc_hd__nor2_1 _30922_ (.A(_02602_),
    .B(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__a21boi_1 _30923_ (.A1(_02596_),
    .A2(_02599_),
    .B1_N(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__o211a_1 _30924_ (.A1(_02602_),
    .A2(_02603_),
    .B1(_02596_),
    .C1(_02599_),
    .X(_02606_));
 sky130_fd_sc_hd__a21boi_1 _30925_ (.A1(_00679_),
    .A2(_00671_),
    .B1_N(_00666_),
    .Y(_02607_));
 sky130_fd_sc_hd__o21ai_1 _30926_ (.A1(_02605_),
    .A2(_02606_),
    .B1(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__a21bo_1 _30927_ (.A1(_02595_),
    .A2(_02599_),
    .B1_N(_02604_),
    .X(_02609_));
 sky130_fd_sc_hd__o211ai_4 _30928_ (.A1(_02602_),
    .A2(_02603_),
    .B1(_02595_),
    .C1(_02599_),
    .Y(_02610_));
 sky130_fd_sc_hd__nand2_1 _30929_ (.A(_00666_),
    .B(_00685_),
    .Y(_02611_));
 sky130_fd_sc_hd__nand3_1 _30930_ (.A(_02609_),
    .B(_02610_),
    .C(_02611_),
    .Y(_02613_));
 sky130_fd_sc_hd__a21oi_1 _30931_ (.A1(_16426_),
    .A2(_07415_),
    .B1(_18377_),
    .Y(_02614_));
 sky130_fd_sc_hd__o22a_1 _30932_ (.A1(_07459_),
    .A2(_00672_),
    .B1(_18373_),
    .B2(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__a21o_1 _30933_ (.A1(_02608_),
    .A2(_02613_),
    .B1(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__a21oi_1 _30934_ (.A1(_02609_),
    .A2(_02610_),
    .B1(_02611_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand3b_1 _30935_ (.A_N(_02617_),
    .B(_02613_),
    .C(_02615_),
    .Y(_02618_));
 sky130_fd_sc_hd__a21bo_1 _30936_ (.A1(_00651_),
    .A2(_00683_),
    .B1_N(_00686_),
    .X(_02619_));
 sky130_fd_sc_hd__a21oi_1 _30937_ (.A1(_02616_),
    .A2(_02618_),
    .B1(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__and3_1 _30938_ (.A(_02619_),
    .B(_02616_),
    .C(_02618_),
    .X(_02621_));
 sky130_fd_sc_hd__nor3_1 _30939_ (.A(_16437_),
    .B(_02620_),
    .C(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__o21a_1 _30940_ (.A1(_02620_),
    .A2(_02621_),
    .B1(_16437_),
    .X(_02624_));
 sky130_fd_sc_hd__a211o_1 _30941_ (.A1(_00695_),
    .A2(_00692_),
    .B1(net140),
    .C1(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__a21oi_1 _30942_ (.A1(_00691_),
    .A2(_07492_),
    .B1(_00690_),
    .Y(_02626_));
 sky130_fd_sc_hd__o21ai_1 _30943_ (.A1(net140),
    .A2(_02624_),
    .B1(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__nand2_1 _30944_ (.A(_02625_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__nand2_1 _30945_ (.A(_02583_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__or2_1 _30946_ (.A(_02628_),
    .B(_02583_),
    .X(_02630_));
 sky130_fd_sc_hd__nand2_1 _30947_ (.A(_02629_),
    .B(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__o21ai_2 _30948_ (.A1(_00706_),
    .A2(_00734_),
    .B1(_00731_),
    .Y(_02632_));
 sky130_fd_sc_hd__nor2_1 _30949_ (.A(_21358_),
    .B(\delay_line[18][11] ),
    .Y(_02633_));
 sky130_fd_sc_hd__buf_1 _30950_ (.A(\delay_line[18][11] ),
    .X(_02635_));
 sky130_fd_sc_hd__nand2_1 _30951_ (.A(_21363_),
    .B(_02635_),
    .Y(_02636_));
 sky130_fd_sc_hd__nand3b_1 _30952_ (.A_N(_02633_),
    .B(_00715_),
    .C(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__inv_2 _30953_ (.A(\delay_line[18][10] ),
    .Y(_02638_));
 sky130_fd_sc_hd__and2_1 _30954_ (.A(_21358_),
    .B(\delay_line[18][11] ),
    .X(_02639_));
 sky130_fd_sc_hd__o22ai_2 _30955_ (.A1(_21356_),
    .A2(_02638_),
    .B1(_02639_),
    .B2(_02633_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand3_1 _30956_ (.A(_21355_),
    .B(_18384_),
    .C(_24704_),
    .Y(_02641_));
 sky130_fd_sc_hd__o21ai_1 _30957_ (.A1(_07514_),
    .A2(_16327_),
    .B1(_18387_),
    .Y(_02642_));
 sky130_fd_sc_hd__nand4_1 _30958_ (.A(_02637_),
    .B(_02640_),
    .C(_02641_),
    .D(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_1 _30959_ (.A(_02637_),
    .B(_02640_),
    .Y(_02644_));
 sky130_fd_sc_hd__nand2_1 _30960_ (.A(_02641_),
    .B(_02642_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand2_1 _30961_ (.A(_02644_),
    .B(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__o21ai_1 _30962_ (.A1(_00715_),
    .A2(_00713_),
    .B1(_00719_),
    .Y(_02648_));
 sky130_fd_sc_hd__a21o_1 _30963_ (.A1(_02643_),
    .A2(_02647_),
    .B1(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__nand2_1 _30964_ (.A(_16338_),
    .B(_01677_),
    .Y(_02650_));
 sky130_fd_sc_hd__nand3_1 _30965_ (.A(_02648_),
    .B(_02643_),
    .C(_02647_),
    .Y(_02651_));
 sky130_fd_sc_hd__and4_1 _30966_ (.A(_02649_),
    .B(_07525_),
    .C(_02650_),
    .D(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__a22oi_2 _30967_ (.A1(_07536_),
    .A2(_02650_),
    .B1(_02649_),
    .B2(_02651_),
    .Y(_02653_));
 sky130_fd_sc_hd__a211o_1 _30968_ (.A1(_00721_),
    .A2(_00724_),
    .B1(_02652_),
    .C1(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__o211ai_2 _30969_ (.A1(_02652_),
    .A2(_02653_),
    .B1(_00721_),
    .C1(_00724_),
    .Y(_02655_));
 sky130_fd_sc_hd__and3_1 _30970_ (.A(_02654_),
    .B(_00725_),
    .C(_02655_),
    .X(_02657_));
 sky130_fd_sc_hd__a21oi_1 _30971_ (.A1(_02655_),
    .A2(_02654_),
    .B1(_00725_),
    .Y(_02658_));
 sky130_fd_sc_hd__o21bai_2 _30972_ (.A1(_02657_),
    .A2(_02658_),
    .B1_N(_00729_),
    .Y(_02659_));
 sky130_fd_sc_hd__nand2_2 _30973_ (.A(_02632_),
    .B(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__nand3_1 _30974_ (.A(_02654_),
    .B(_00725_),
    .C(_02655_),
    .Y(_02661_));
 sky130_fd_sc_hd__nand3b_2 _30975_ (.A_N(_02658_),
    .B(_00729_),
    .C(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__a21o_1 _30976_ (.A1(_02662_),
    .A2(_02659_),
    .B1(_02632_),
    .X(_02663_));
 sky130_fd_sc_hd__nand3b_4 _30977_ (.A_N(_02631_),
    .B(_02660_),
    .C(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hd__inv_2 _30978_ (.A(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__a21boi_2 _30979_ (.A1(_02663_),
    .A2(_02660_),
    .B1_N(_02631_),
    .Y(_02666_));
 sky130_fd_sc_hd__o22ai_2 _30980_ (.A1(_02581_),
    .A2(_02582_),
    .B1(_02665_),
    .B2(_02666_),
    .Y(_02668_));
 sky130_fd_sc_hd__or4_2 _30981_ (.A(_02581_),
    .B(_02582_),
    .C(_02665_),
    .D(_02666_),
    .X(_02669_));
 sky130_fd_sc_hd__and3_2 _30982_ (.A(_02539_),
    .B(_02668_),
    .C(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__a21oi_1 _30983_ (.A1(_02669_),
    .A2(_02668_),
    .B1(_02539_),
    .Y(_02671_));
 sky130_fd_sc_hd__nor2_2 _30984_ (.A(_02670_),
    .B(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__o21a_1 _30985_ (.A1(_00739_),
    .A2(_00872_),
    .B1(_00871_),
    .X(_02673_));
 sky130_fd_sc_hd__xor2_4 _30986_ (.A(_02672_),
    .B(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__xor2_4 _30987_ (.A(_02404_),
    .B(_02674_),
    .X(_02675_));
 sky130_fd_sc_hd__xor2_1 _30988_ (.A(_02266_),
    .B(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__xnor2_1 _30989_ (.A(_02265_),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__xnor2_1 _30990_ (.A(_02071_),
    .B(_02677_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand3_1 _30991_ (.A(_01212_),
    .B(_01213_),
    .C(_01322_),
    .Y(_02680_));
 sky130_fd_sc_hd__a21oi_2 _30992_ (.A1(_01060_),
    .A2(_01061_),
    .B1(_01059_),
    .Y(_02681_));
 sky130_fd_sc_hd__nor2_1 _30993_ (.A(_01223_),
    .B(net285),
    .Y(_02682_));
 sky130_fd_sc_hd__and2_1 _30994_ (.A(_01223_),
    .B(net285),
    .X(_02683_));
 sky130_fd_sc_hd__buf_1 _30995_ (.A(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__a2111oi_1 _30996_ (.A1(_25032_),
    .A2(_01224_),
    .B1(_02682_),
    .C1(_02684_),
    .D1(_01220_),
    .Y(_02685_));
 sky130_fd_sc_hd__buf_1 _30997_ (.A(\delay_line[38][10] ),
    .X(_02686_));
 sky130_fd_sc_hd__and3_1 _30998_ (.A(_23434_),
    .B(_02686_),
    .C(_01221_),
    .X(_02687_));
 sky130_fd_sc_hd__o22a_1 _30999_ (.A1(_02682_),
    .A2(_02683_),
    .B1(_02687_),
    .B2(_01220_),
    .X(_02688_));
 sky130_fd_sc_hd__a2111oi_1 _31000_ (.A1(_01224_),
    .A2(_01218_),
    .B1(_01226_),
    .C1(net254),
    .D1(_02688_),
    .Y(_02690_));
 sky130_fd_sc_hd__and4_1 _31001_ (.A(_23429_),
    .B(_01223_),
    .C(_25034_),
    .D(_01224_),
    .X(_02691_));
 sky130_fd_sc_hd__o22a_1 _31002_ (.A1(net255),
    .A2(_02688_),
    .B1(_02691_),
    .B2(_01226_),
    .X(_02692_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31003_ (.A(_01231_),
    .X(_02693_));
 sky130_fd_sc_hd__nand2_1 _31004_ (.A(_02693_),
    .B(_01233_),
    .Y(_02694_));
 sky130_fd_sc_hd__nor2_1 _31005_ (.A(_01233_),
    .B(\delay_line[39][12] ),
    .Y(_02695_));
 sky130_fd_sc_hd__and2_1 _31006_ (.A(_01233_),
    .B(\delay_line[39][12] ),
    .X(_02696_));
 sky130_fd_sc_hd__or3b_1 _31007_ (.A(_02695_),
    .B(_02696_),
    .C_N(_01231_),
    .X(_02697_));
 sky130_fd_sc_hd__o21bai_1 _31008_ (.A1(_02695_),
    .A2(_02696_),
    .B1_N(_02693_),
    .Y(_02698_));
 sky130_fd_sc_hd__nand2_1 _31009_ (.A(_02697_),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__a21oi_2 _31010_ (.A1(_02694_),
    .A2(_01236_),
    .B1(_02699_),
    .Y(_02701_));
 sky130_fd_sc_hd__a311oi_2 _31011_ (.A1(_01234_),
    .A2(_02694_),
    .A3(_02699_),
    .B1(_23446_),
    .C1(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__and3_1 _31012_ (.A(_02694_),
    .B(_01236_),
    .C(_02699_),
    .X(_02703_));
 sky130_fd_sc_hd__o21a_1 _31013_ (.A1(_02701_),
    .A2(_02703_),
    .B1(_23446_),
    .X(_02704_));
 sky130_fd_sc_hd__or2_1 _31014_ (.A(_02702_),
    .B(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__or2b_1 _31015_ (.A(_01240_),
    .B_N(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__o21bai_1 _31016_ (.A1(_01240_),
    .A2(_01241_),
    .B1_N(_02705_),
    .Y(_02707_));
 sky130_fd_sc_hd__o221a_2 _31017_ (.A1(_02706_),
    .A2(_01241_),
    .B1(_01246_),
    .B2(_01250_),
    .C1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__o21a_1 _31018_ (.A1(_01241_),
    .A2(_02706_),
    .B1(_02707_),
    .X(_02709_));
 sky130_fd_sc_hd__or3_1 _31019_ (.A(_01246_),
    .B(_01250_),
    .C(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__inv_2 _31020_ (.A(_02710_),
    .Y(_02712_));
 sky130_fd_sc_hd__or4_2 _31021_ (.A(net134),
    .B(_02692_),
    .C(_02708_),
    .D(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__inv_2 _31022_ (.A(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__o22a_1 _31023_ (.A1(net133),
    .A2(_02692_),
    .B1(_02708_),
    .B2(_02712_),
    .X(_02715_));
 sky130_fd_sc_hd__o211ai_1 _31024_ (.A1(_01257_),
    .A2(_01258_),
    .B1(_25047_),
    .C1(_25050_),
    .Y(_02716_));
 sky130_fd_sc_hd__and2_1 _31025_ (.A(_02716_),
    .B(_01262_),
    .X(_02717_));
 sky130_fd_sc_hd__nand2_1 _31026_ (.A(\delay_line[40][11] ),
    .B(\delay_line[40][12] ),
    .Y(_02718_));
 sky130_fd_sc_hd__inv_2 _31027_ (.A(\delay_line[40][11] ),
    .Y(_02719_));
 sky130_fd_sc_hd__o21bai_1 _31028_ (.A1(_01254_),
    .A2(_02719_),
    .B1_N(\delay_line[40][12] ),
    .Y(_02720_));
 sky130_fd_sc_hd__o21a_1 _31029_ (.A1(_01254_),
    .A2(_02718_),
    .B1(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__xor2_1 _31030_ (.A(_23464_),
    .B(_02721_),
    .X(_02723_));
 sky130_fd_sc_hd__a31o_1 _31031_ (.A1(_23465_),
    .A2(_01254_),
    .A3(_02719_),
    .B1(_01257_),
    .X(_02724_));
 sky130_fd_sc_hd__xor2_1 _31032_ (.A(_02723_),
    .B(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__o21a_1 _31033_ (.A1(_01261_),
    .A2(_02717_),
    .B1(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__a211oi_1 _31034_ (.A1(_02716_),
    .A2(_01262_),
    .B1(_02725_),
    .C1(_01261_),
    .Y(_02727_));
 sky130_fd_sc_hd__or2_2 _31035_ (.A(_02726_),
    .B(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__o21ai_1 _31036_ (.A1(_02714_),
    .A2(_02715_),
    .B1(_02728_),
    .Y(_02729_));
 sky130_fd_sc_hd__or3_1 _31037_ (.A(_02715_),
    .B(_02728_),
    .C(_02714_),
    .X(_02730_));
 sky130_fd_sc_hd__and2_2 _31038_ (.A(_02729_),
    .B(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31039_ (.A(\delay_line[37][11] ),
    .X(_02732_));
 sky130_fd_sc_hd__or2b_1 _31040_ (.A(_23521_),
    .B_N(_02732_),
    .X(_02734_));
 sky130_fd_sc_hd__nand3b_1 _31041_ (.A_N(_21036_),
    .B(_01269_),
    .C(_01272_),
    .Y(_02735_));
 sky130_fd_sc_hd__xnor2_1 _31042_ (.A(\delay_line[37][10] ),
    .B(\delay_line[37][12] ),
    .Y(_02736_));
 sky130_fd_sc_hd__a21oi_1 _31043_ (.A1(_02734_),
    .A2(_02735_),
    .B1(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__and3_1 _31044_ (.A(_02734_),
    .B(_02735_),
    .C(_02736_),
    .X(_02738_));
 sky130_fd_sc_hd__nor2_1 _31045_ (.A(_02737_),
    .B(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__a41oi_2 _31046_ (.A1(_02732_),
    .A2(_25068_),
    .A3(_25066_),
    .A4(_25067_),
    .B1(_01275_),
    .Y(_02740_));
 sky130_fd_sc_hd__xnor2_1 _31047_ (.A(_02739_),
    .B(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__nor2_1 _31048_ (.A(_20833_),
    .B(_01302_),
    .Y(_02742_));
 sky130_fd_sc_hd__nor3b_1 _31049_ (.A(_01291_),
    .B(_01292_),
    .C_N(_25098_),
    .Y(_02743_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31050_ (.A(\delay_line[35][11] ),
    .X(_02745_));
 sky130_fd_sc_hd__nor2_1 _31051_ (.A(_02745_),
    .B(\delay_line[35][12] ),
    .Y(_02746_));
 sky130_fd_sc_hd__and2_1 _31052_ (.A(\delay_line[35][11] ),
    .B(net301),
    .X(_02747_));
 sky130_fd_sc_hd__or3b_1 _31053_ (.A(_02746_),
    .B(_02747_),
    .C_N(_25091_),
    .X(_02748_));
 sky130_fd_sc_hd__o21bai_1 _31054_ (.A1(_02746_),
    .A2(_02747_),
    .B1_N(_25091_),
    .Y(_02749_));
 sky130_fd_sc_hd__o211a_1 _31055_ (.A1(_01292_),
    .A2(_02743_),
    .B1(_02748_),
    .C1(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__a221oi_2 _31056_ (.A1(_01290_),
    .A2(_02745_),
    .B1(_02748_),
    .B2(_02749_),
    .C1(_02743_),
    .Y(_02751_));
 sky130_fd_sc_hd__nor3_1 _31057_ (.A(_01298_),
    .B(_02750_),
    .C(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__o21ai_1 _31058_ (.A1(_02750_),
    .A2(_02751_),
    .B1(_01298_),
    .Y(_02753_));
 sky130_fd_sc_hd__inv_2 _31059_ (.A(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__or3_1 _31060_ (.A(_20837_),
    .B(_02752_),
    .C(_02754_),
    .X(_02756_));
 sky130_fd_sc_hd__o21ai_1 _31061_ (.A1(_02752_),
    .A2(_02754_),
    .B1(_20837_),
    .Y(_02757_));
 sky130_fd_sc_hd__o211ai_2 _31062_ (.A1(_01299_),
    .A2(_02742_),
    .B1(_02756_),
    .C1(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__a211o_1 _31063_ (.A1(_02756_),
    .A2(_02757_),
    .B1(_01299_),
    .C1(_02742_),
    .X(_02759_));
 sky130_fd_sc_hd__a221o_1 _31064_ (.A1(_02758_),
    .A2(_02759_),
    .B1(_01309_),
    .B2(_01308_),
    .C1(_01305_),
    .X(_02760_));
 sky130_fd_sc_hd__nand2_1 _31065_ (.A(_02758_),
    .B(_02759_),
    .Y(_02761_));
 sky130_fd_sc_hd__a21oi_1 _31066_ (.A1(_01309_),
    .A2(_01308_),
    .B1(_01305_),
    .Y(_02762_));
 sky130_fd_sc_hd__or2_1 _31067_ (.A(_02761_),
    .B(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__buf_1 _31068_ (.A(\delay_line[36][8] ),
    .X(_02764_));
 sky130_fd_sc_hd__nand2_1 _31069_ (.A(_02764_),
    .B(_01280_),
    .Y(_02765_));
 sky130_fd_sc_hd__and2b_1 _31070_ (.A_N(_25077_),
    .B(_02764_),
    .X(_02767_));
 sky130_fd_sc_hd__and2b_1 _31071_ (.A_N(net297),
    .B(net296),
    .X(_02768_));
 sky130_fd_sc_hd__and2b_1 _31072_ (.A_N(net296),
    .B(\delay_line[36][7] ),
    .X(_02769_));
 sky130_fd_sc_hd__nor2_1 _31073_ (.A(_02768_),
    .B(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__a211oi_2 _31074_ (.A1(_01279_),
    .A2(_01281_),
    .B1(_02767_),
    .C1(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__and3_1 _31075_ (.A(_01278_),
    .B(_01279_),
    .C(_01281_),
    .X(_02772_));
 sky130_fd_sc_hd__o21a_1 _31076_ (.A1(_02767_),
    .A2(_02772_),
    .B1(_02770_),
    .X(_02773_));
 sky130_fd_sc_hd__a211oi_2 _31077_ (.A1(_01288_),
    .A2(_02765_),
    .B1(_02771_),
    .C1(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__o211a_1 _31078_ (.A1(_02773_),
    .A2(_02771_),
    .B1(_02765_),
    .C1(_01288_),
    .X(_02775_));
 sky130_fd_sc_hd__or2_1 _31079_ (.A(_02774_),
    .B(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__a21boi_1 _31080_ (.A1(_02760_),
    .A2(_02763_),
    .B1_N(_02776_),
    .Y(_02778_));
 sky130_fd_sc_hd__nand3b_1 _31081_ (.A_N(_02776_),
    .B(_02760_),
    .C(_02763_),
    .Y(_02779_));
 sky130_fd_sc_hd__or2b_1 _31082_ (.A(_02778_),
    .B_N(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__xnor2_1 _31083_ (.A(_02741_),
    .B(_02780_),
    .Y(_02781_));
 sky130_fd_sc_hd__and3b_1 _31084_ (.A_N(_01312_),
    .B(_01314_),
    .C(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__o21ba_1 _31085_ (.A1(_01277_),
    .A2(_01313_),
    .B1_N(_01312_),
    .X(_02783_));
 sky130_fd_sc_hd__nor2_1 _31086_ (.A(_02783_),
    .B(_02781_),
    .Y(_02784_));
 sky130_fd_sc_hd__nor2_2 _31087_ (.A(_02782_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__xnor2_4 _31088_ (.A(_02731_),
    .B(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__o21ai_4 _31089_ (.A1(_00914_),
    .A2(_00962_),
    .B1(_00960_),
    .Y(_02787_));
 sky130_fd_sc_hd__nor2_1 _31090_ (.A(_01146_),
    .B(_01147_),
    .Y(_02789_));
 sky130_fd_sc_hd__and3_1 _31091_ (.A(_24947_),
    .B(_01151_),
    .C(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__or4_1 _31092_ (.A(_02128_),
    .B(_01133_),
    .C(_19611_),
    .D(_01131_),
    .X(_02791_));
 sky130_fd_sc_hd__nor2_1 _31093_ (.A(_01111_),
    .B(\delay_line[32][12] ),
    .Y(_02792_));
 sky130_fd_sc_hd__buf_1 _31094_ (.A(\delay_line[32][12] ),
    .X(_02793_));
 sky130_fd_sc_hd__nand2_1 _31095_ (.A(_01111_),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__clkbuf_2 _31096_ (.A(\delay_line[32][10] ),
    .X(_02795_));
 sky130_fd_sc_hd__nand3b_2 _31097_ (.A_N(_02792_),
    .B(_02794_),
    .C(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__and2_1 _31098_ (.A(_01111_),
    .B(\delay_line[32][12] ),
    .X(_02797_));
 sky130_fd_sc_hd__o21bai_1 _31099_ (.A1(_02792_),
    .A2(_02797_),
    .B1_N(_24956_),
    .Y(_02798_));
 sky130_fd_sc_hd__o21ai_1 _31100_ (.A1(_01119_),
    .A2(_01112_),
    .B1(_01114_),
    .Y(_02800_));
 sky130_fd_sc_hd__a21oi_1 _31101_ (.A1(_02796_),
    .A2(_02798_),
    .B1(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__and3_1 _31102_ (.A(_02796_),
    .B(_02798_),
    .C(_02800_),
    .X(_02802_));
 sky130_fd_sc_hd__buf_1 _31103_ (.A(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__nor3_1 _31104_ (.A(_02801_),
    .B(_01119_),
    .C(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31105_ (.A(_01119_),
    .X(_02805_));
 sky130_fd_sc_hd__o21a_1 _31106_ (.A1(_02803_),
    .A2(_02801_),
    .B1(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__a21oi_1 _31107_ (.A1(_01116_),
    .A2(_01120_),
    .B1(_01122_),
    .Y(_02807_));
 sky130_fd_sc_hd__o21ai_1 _31108_ (.A1(_01121_),
    .A2(_02807_),
    .B1(_01123_),
    .Y(_02808_));
 sky130_fd_sc_hd__o21bai_1 _31109_ (.A1(_02804_),
    .A2(_02806_),
    .B1_N(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__a21o_1 _31110_ (.A1(_02796_),
    .A2(_02798_),
    .B1(_02800_),
    .X(_02811_));
 sky130_fd_sc_hd__nand3b_1 _31111_ (.A_N(_02802_),
    .B(_02811_),
    .C(_01115_),
    .Y(_02812_));
 sky130_fd_sc_hd__o21ai_1 _31112_ (.A1(_02803_),
    .A2(_02801_),
    .B1(_02805_),
    .Y(_02813_));
 sky130_fd_sc_hd__nand3_2 _31113_ (.A(_02808_),
    .B(_02812_),
    .C(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__nor2_1 _31114_ (.A(_18659_),
    .B(_21112_),
    .Y(_02815_));
 sky130_fd_sc_hd__nor2_1 _31115_ (.A(_20699_),
    .B(_18672_),
    .Y(_02816_));
 sky130_fd_sc_hd__nor2_1 _31116_ (.A(_02815_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__xor2_1 _31117_ (.A(_01131_),
    .B(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__and3_1 _31118_ (.A(_02809_),
    .B(_02814_),
    .C(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__a21oi_1 _31119_ (.A1(_02809_),
    .A2(_02814_),
    .B1(_02818_),
    .Y(_02820_));
 sky130_fd_sc_hd__o211a_1 _31120_ (.A1(_02819_),
    .A2(_02820_),
    .B1(_01130_),
    .C1(_01136_),
    .X(_02822_));
 sky130_fd_sc_hd__a211o_1 _31121_ (.A1(_01130_),
    .A2(_01136_),
    .B1(_02819_),
    .C1(_02820_),
    .X(_02823_));
 sky130_fd_sc_hd__inv_2 _31122_ (.A(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__nor3_1 _31123_ (.A(_02791_),
    .B(_02822_),
    .C(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__buf_1 _31124_ (.A(_01131_),
    .X(_02826_));
 sky130_fd_sc_hd__o32a_1 _31125_ (.A1(_24949_),
    .A2(_02826_),
    .A3(_01133_),
    .B1(_02822_),
    .B2(_02824_),
    .X(_02827_));
 sky130_fd_sc_hd__a211oi_1 _31126_ (.A1(_01141_),
    .A2(_01142_),
    .B1(_02825_),
    .C1(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__o211a_1 _31127_ (.A1(_02825_),
    .A2(_02827_),
    .B1(_01141_),
    .C1(_01142_),
    .X(_02829_));
 sky130_fd_sc_hd__nor2_1 _31128_ (.A(_02828_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__xor2_2 _31129_ (.A(_01146_),
    .B(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__o21ai_2 _31130_ (.A1(_02790_),
    .A2(_01156_),
    .B1(_02831_),
    .Y(_02833_));
 sky130_fd_sc_hd__a311o_1 _31131_ (.A1(_24947_),
    .A2(_01151_),
    .A3(_02789_),
    .B1(_01156_),
    .C1(_02831_),
    .X(_02834_));
 sky130_fd_sc_hd__nor2_1 _31132_ (.A(_01169_),
    .B(_01171_),
    .Y(_02835_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31133_ (.A(_19576_),
    .X(_02836_));
 sky130_fd_sc_hd__and3_1 _31134_ (.A(_05348_),
    .B(_01160_),
    .C(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__inv_2 _31135_ (.A(\delay_line[33][12] ),
    .Y(_02838_));
 sky130_fd_sc_hd__nand2_1 _31136_ (.A(_23356_),
    .B(_20666_),
    .Y(_02839_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31137_ (.A(_21161_),
    .X(_02840_));
 sky130_fd_sc_hd__nand2_1 _31138_ (.A(_20671_),
    .B(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__nand3_1 _31139_ (.A(_02838_),
    .B(_02839_),
    .C(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__a21o_1 _31140_ (.A1(_02839_),
    .A2(_02841_),
    .B1(_02838_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_2 _31141_ (.A(_01163_),
    .X(_02845_));
 sky130_fd_sc_hd__a21oi_1 _31142_ (.A1(_01164_),
    .A2(_01165_),
    .B1(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__a21oi_1 _31143_ (.A1(_02842_),
    .A2(_02844_),
    .B1(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__clkbuf_2 _31144_ (.A(_20671_),
    .X(_02848_));
 sky130_fd_sc_hd__a21oi_1 _31145_ (.A1(_02848_),
    .A2(_19576_),
    .B1(_24914_),
    .Y(_02849_));
 sky130_fd_sc_hd__nand2_1 _31146_ (.A(_23366_),
    .B(_24913_),
    .Y(_02850_));
 sky130_fd_sc_hd__a31o_1 _31147_ (.A1(_24914_),
    .A2(_02836_),
    .A3(_02848_),
    .B1(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__and3_1 _31148_ (.A(_24914_),
    .B(_20671_),
    .C(_19576_),
    .X(_02852_));
 sky130_fd_sc_hd__o21ai_1 _31149_ (.A1(_02852_),
    .A2(_02849_),
    .B1(_02850_),
    .Y(_02853_));
 sky130_fd_sc_hd__o21ai_1 _31150_ (.A1(_02849_),
    .A2(_02851_),
    .B1(_02853_),
    .Y(_02855_));
 sky130_fd_sc_hd__and3_1 _31151_ (.A(_02844_),
    .B(_02846_),
    .C(_02842_),
    .X(_02856_));
 sky130_fd_sc_hd__nor3_1 _31152_ (.A(_02847_),
    .B(_02855_),
    .C(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__o21a_1 _31153_ (.A1(_02856_),
    .A2(_02847_),
    .B1(_02855_),
    .X(_02858_));
 sky130_fd_sc_hd__nor2_1 _31154_ (.A(_02857_),
    .B(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__a311o_1 _31155_ (.A1(_24927_),
    .A2(_01166_),
    .A3(_01167_),
    .B1(_01177_),
    .C1(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__o21ai_2 _31156_ (.A1(_01176_),
    .A2(_01177_),
    .B1(_02859_),
    .Y(_02861_));
 sky130_fd_sc_hd__o211a_1 _31157_ (.A1(_02835_),
    .A2(_02837_),
    .B1(_02860_),
    .C1(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__a211oi_1 _31158_ (.A1(_02860_),
    .A2(_02861_),
    .B1(_02835_),
    .C1(_02837_),
    .Y(_02863_));
 sky130_fd_sc_hd__a211o_1 _31159_ (.A1(_01185_),
    .A2(_01192_),
    .B1(_02862_),
    .C1(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__and3_1 _31160_ (.A(_01192_),
    .B(_01193_),
    .C(_01190_),
    .X(_02866_));
 sky130_fd_sc_hd__o211ai_1 _31161_ (.A1(_02862_),
    .A2(_02863_),
    .B1(_01185_),
    .C1(_01192_),
    .Y(_02867_));
 sky130_fd_sc_hd__and3_1 _31162_ (.A(_02864_),
    .B(_02866_),
    .C(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__a21oi_1 _31163_ (.A1(_02867_),
    .A2(_02864_),
    .B1(_02866_),
    .Y(_02869_));
 sky130_fd_sc_hd__nor2_1 _31164_ (.A(_02868_),
    .B(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__a32oi_4 _31165_ (.A1(_01158_),
    .A2(_01191_),
    .A3(_01195_),
    .B1(_01199_),
    .B2(_01198_),
    .Y(_02871_));
 sky130_fd_sc_hd__xnor2_1 _31166_ (.A(_02870_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__a21o_1 _31167_ (.A1(_02833_),
    .A2(_02834_),
    .B1(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__nand3_2 _31168_ (.A(_02834_),
    .B(_02872_),
    .C(_02833_),
    .Y(_02874_));
 sky130_fd_sc_hd__nand2_1 _31169_ (.A(_02873_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__inv_2 _31170_ (.A(_01096_),
    .Y(_02877_));
 sky130_fd_sc_hd__and2_1 _31171_ (.A(_01076_),
    .B(_24873_),
    .X(_02878_));
 sky130_fd_sc_hd__nor2_1 _31172_ (.A(_24873_),
    .B(_01076_),
    .Y(_02879_));
 sky130_fd_sc_hd__clkbuf_2 _31173_ (.A(_01078_),
    .X(_02880_));
 sky130_fd_sc_hd__or2_1 _31174_ (.A(_01072_),
    .B(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__nand2_2 _31175_ (.A(_01072_),
    .B(_02880_),
    .Y(_02882_));
 sky130_fd_sc_hd__buf_1 _31176_ (.A(net305),
    .X(_02883_));
 sky130_fd_sc_hd__nor2_1 _31177_ (.A(_24880_),
    .B(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__and2_1 _31178_ (.A(_24880_),
    .B(net305),
    .X(_02885_));
 sky130_fd_sc_hd__or3_2 _31179_ (.A(_02884_),
    .B(_01080_),
    .C(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__a2bb2o_1 _31180_ (.A1_N(_02885_),
    .A2_N(_02884_),
    .B1(_01078_),
    .B2(_01079_),
    .X(_02888_));
 sky130_fd_sc_hd__a22o_1 _31181_ (.A1(_02881_),
    .A2(_02882_),
    .B1(_02886_),
    .B2(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__nand4_2 _31182_ (.A(_02881_),
    .B(_02882_),
    .C(_02886_),
    .D(_02888_),
    .Y(_02890_));
 sky130_fd_sc_hd__nand2_1 _31183_ (.A(_01081_),
    .B(_01085_),
    .Y(_02891_));
 sky130_fd_sc_hd__a21o_1 _31184_ (.A1(_02889_),
    .A2(_02890_),
    .B1(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__nand3_1 _31185_ (.A(_02891_),
    .B(_02889_),
    .C(_02890_),
    .Y(_02893_));
 sky130_fd_sc_hd__a2bb2oi_1 _31186_ (.A1_N(_02878_),
    .A2_N(_02879_),
    .B1(_02892_),
    .B2(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__and4bb_2 _31187_ (.A_N(_02878_),
    .B_N(_02879_),
    .C(_02892_),
    .D(_02893_),
    .X(_02895_));
 sky130_fd_sc_hd__a211oi_2 _31188_ (.A1(_01090_),
    .A2(_02877_),
    .B1(_02894_),
    .C1(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__o221ai_2 _31189_ (.A1(_01088_),
    .A2(_01087_),
    .B1(_02894_),
    .B2(_02895_),
    .C1(_02877_),
    .Y(_02897_));
 sky130_fd_sc_hd__or4bb_2 _31190_ (.A(_17812_),
    .B(_02896_),
    .C_N(_24887_),
    .D_N(_02897_),
    .X(_02899_));
 sky130_fd_sc_hd__inv_2 _31191_ (.A(_02896_),
    .Y(_02900_));
 sky130_fd_sc_hd__a21o_1 _31192_ (.A1(_02897_),
    .A2(_02900_),
    .B1(_01092_),
    .X(_02901_));
 sky130_fd_sc_hd__a221o_1 _31193_ (.A1(_24878_),
    .A2(_01099_),
    .B1(_02899_),
    .B2(_02901_),
    .C1(_01098_),
    .X(_02902_));
 sky130_fd_sc_hd__and4b_1 _31194_ (.A_N(_05403_),
    .B(_24873_),
    .C(_24876_),
    .D(_01099_),
    .X(_02903_));
 sky130_fd_sc_hd__o211ai_2 _31195_ (.A1(_01098_),
    .A2(_02903_),
    .B1(_02899_),
    .C1(_02901_),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2_1 _31196_ (.A(_02902_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__a21oi_2 _31197_ (.A1(_01103_),
    .A2(_01108_),
    .B1(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__o211ai_1 _31198_ (.A1(_01101_),
    .A2(_01100_),
    .B1(_02905_),
    .C1(_01108_),
    .Y(_02907_));
 sky130_fd_sc_hd__or2b_1 _31199_ (.A(_02906_),
    .B_N(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__xor2_1 _31200_ (.A(_02875_),
    .B(_02908_),
    .X(_02910_));
 sky130_fd_sc_hd__xnor2_1 _31201_ (.A(_02787_),
    .B(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__a21o_1 _31202_ (.A1(_01109_),
    .A2(_01204_),
    .B1(_01202_),
    .X(_02912_));
 sky130_fd_sc_hd__and2b_1 _31203_ (.A_N(_02911_),
    .B(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__and2b_1 _31204_ (.A_N(_02912_),
    .B(_02911_),
    .X(_02914_));
 sky130_fd_sc_hd__nor2_1 _31205_ (.A(_02913_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__or3_1 _31206_ (.A(_01208_),
    .B(_01211_),
    .C(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__o21ai_1 _31207_ (.A1(_01208_),
    .A2(_01211_),
    .B1(_02915_),
    .Y(_02917_));
 sky130_fd_sc_hd__nand2_1 _31208_ (.A(_02916_),
    .B(_02917_),
    .Y(_02918_));
 sky130_fd_sc_hd__xnor2_2 _31209_ (.A(_02786_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__xnor2_1 _31210_ (.A(_02681_),
    .B(_02919_),
    .Y(_02921_));
 sky130_fd_sc_hd__and3_1 _31211_ (.A(_01212_),
    .B(_02680_),
    .C(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__a21o_1 _31212_ (.A1(_01212_),
    .A2(_02680_),
    .B1(_02921_),
    .X(_02923_));
 sky130_fd_sc_hd__or2b_1 _31213_ (.A(_02922_),
    .B_N(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__xnor2_1 _31214_ (.A(_02679_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__xnor2_2 _31215_ (.A(_02070_),
    .B(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__nand2_1 _31216_ (.A(_02067_),
    .B(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__a21oi_1 _31217_ (.A1(_02058_),
    .A2(_02065_),
    .B1(_01475_),
    .Y(_02928_));
 sky130_fd_sc_hd__o21bai_2 _31218_ (.A1(_02928_),
    .A2(_02066_),
    .B1_N(_02926_),
    .Y(_02929_));
 sky130_fd_sc_hd__a31o_1 _31219_ (.A1(_00460_),
    .A2(_00462_),
    .A3(_01334_),
    .B1(_01332_),
    .X(_02930_));
 sky130_fd_sc_hd__o211ai_4 _31220_ (.A1(_02066_),
    .A2(_02927_),
    .B1(_02929_),
    .C1(_02930_),
    .Y(_02932_));
 sky130_fd_sc_hd__o221a_1 _31221_ (.A1(_01476_),
    .A2(_01477_),
    .B1(_02037_),
    .B2(_02050_),
    .C1(_02057_),
    .X(_02933_));
 sky130_fd_sc_hd__a32o_1 _31222_ (.A1(_02060_),
    .A2(_02061_),
    .A3(_02064_),
    .B1(_01474_),
    .B2(_00450_),
    .X(_02934_));
 sky130_fd_sc_hd__o211ai_2 _31223_ (.A1(_02933_),
    .A2(_02934_),
    .B1(_02067_),
    .C1(_02926_),
    .Y(_02935_));
 sky130_fd_sc_hd__a21o_1 _31224_ (.A1(_02929_),
    .A2(_02935_),
    .B1(_02930_),
    .X(_02936_));
 sky130_fd_sc_hd__o2111ai_1 _31225_ (.A1(_01470_),
    .A2(_01471_),
    .B1(_01473_),
    .C1(_02932_),
    .D1(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__and3_1 _31226_ (.A(_02930_),
    .B(_02929_),
    .C(_02935_),
    .X(_02938_));
 sky130_fd_sc_hd__a21oi_1 _31227_ (.A1(_02929_),
    .A2(_02935_),
    .B1(_02930_),
    .Y(_02939_));
 sky130_fd_sc_hd__o21ai_2 _31228_ (.A1(_01471_),
    .A2(_01470_),
    .B1(_01473_),
    .Y(_02940_));
 sky130_fd_sc_hd__o21ai_1 _31229_ (.A1(_02938_),
    .A2(_02939_),
    .B1(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__nand3_1 _31230_ (.A(_01404_),
    .B(_02937_),
    .C(_02941_),
    .Y(_02943_));
 sky130_fd_sc_hd__a21o_1 _31231_ (.A1(_02932_),
    .A2(_02936_),
    .B1(_02940_),
    .X(_02944_));
 sky130_fd_sc_hd__nand3_1 _31232_ (.A(_02940_),
    .B(_02932_),
    .C(_02936_),
    .Y(_02945_));
 sky130_fd_sc_hd__o21a_1 _31233_ (.A1(_25285_),
    .A2(_01403_),
    .B1(_01341_),
    .X(_02946_));
 sky130_fd_sc_hd__nand3_1 _31234_ (.A(_02944_),
    .B(_02945_),
    .C(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__nand2_1 _31235_ (.A(_02943_),
    .B(_02947_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2_1 _31236_ (.A(_25282_),
    .B(_25280_),
    .Y(_02949_));
 sky130_fd_sc_hd__o21a_1 _31237_ (.A1(_04953_),
    .A2(_10778_),
    .B1(_19827_),
    .X(_02950_));
 sky130_fd_sc_hd__or2_1 _31238_ (.A(_20964_),
    .B(_10844_),
    .X(_02951_));
 sky130_fd_sc_hd__nand2_2 _31239_ (.A(_19809_),
    .B(_10844_),
    .Y(_02952_));
 sky130_fd_sc_hd__o211a_1 _31240_ (.A1(_05172_),
    .A2(_02950_),
    .B1(_02951_),
    .C1(_02952_),
    .X(_02954_));
 sky130_fd_sc_hd__a221oi_1 _31241_ (.A1(_04953_),
    .A2(_20898_),
    .B1(_02951_),
    .B2(_02952_),
    .C1(_02950_),
    .Y(_02955_));
 sky130_fd_sc_hd__nor2_1 _31242_ (.A(_02954_),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__or3_1 _31243_ (.A(_25241_),
    .B(_25245_),
    .C(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__o21ai_2 _31244_ (.A1(_25241_),
    .A2(_25245_),
    .B1(_02956_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand3_1 _31245_ (.A(_02957_),
    .B(_01360_),
    .C(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__a32o_1 _31246_ (.A1(_01357_),
    .A2(_01355_),
    .A3(_01356_),
    .B1(_02958_),
    .B2(_02957_),
    .X(_02960_));
 sky130_fd_sc_hd__nand2_1 _31247_ (.A(_02959_),
    .B(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__o211ai_4 _31248_ (.A1(_25246_),
    .A2(_25272_),
    .B1(_25273_),
    .C1(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__or3_1 _31249_ (.A(_25244_),
    .B(_25245_),
    .C(_25274_),
    .X(_02963_));
 sky130_fd_sc_hd__a21o_2 _31250_ (.A1(_25273_),
    .A2(_02963_),
    .B1(_02961_),
    .X(_02965_));
 sky130_fd_sc_hd__a221o_1 _31251_ (.A1(_01354_),
    .A2(_01361_),
    .B1(_02962_),
    .B2(_02965_),
    .C1(_01364_),
    .X(_02966_));
 sky130_fd_sc_hd__o211ai_4 _31252_ (.A1(_01363_),
    .A2(_01364_),
    .B1(_02962_),
    .C1(_02965_),
    .Y(_02967_));
 sky130_fd_sc_hd__o21ai_2 _31253_ (.A1(_01353_),
    .A2(_01371_),
    .B1(_01369_),
    .Y(_02968_));
 sky130_fd_sc_hd__a21oi_1 _31254_ (.A1(_02966_),
    .A2(_02967_),
    .B1(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__and3_1 _31255_ (.A(_02968_),
    .B(_02966_),
    .C(_02967_),
    .X(_02970_));
 sky130_fd_sc_hd__or2_1 _31256_ (.A(_02969_),
    .B(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__a21oi_1 _31257_ (.A1(_25277_),
    .A2(_02949_),
    .B1(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__nand3_1 _31258_ (.A(_25277_),
    .B(_02949_),
    .C(_02971_),
    .Y(_02973_));
 sky130_fd_sc_hd__and2b_1 _31259_ (.A_N(_02972_),
    .B(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__xor2_1 _31260_ (.A(_01373_),
    .B(_02974_),
    .X(_02976_));
 sky130_fd_sc_hd__nand2_1 _31261_ (.A(_02948_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__a32oi_4 _31262_ (.A1(_01349_),
    .A2(_01350_),
    .A3(_01351_),
    .B1(_01347_),
    .B2(_01386_),
    .Y(_02978_));
 sky130_fd_sc_hd__xnor2_1 _31263_ (.A(_01373_),
    .B(_02974_),
    .Y(_02979_));
 sky130_fd_sc_hd__nand3_1 _31264_ (.A(_02979_),
    .B(_02943_),
    .C(_02947_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand3_1 _31265_ (.A(_02977_),
    .B(_02978_),
    .C(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__a21o_1 _31266_ (.A1(_02980_),
    .A2(_02977_),
    .B1(_02978_),
    .X(_02982_));
 sky130_fd_sc_hd__or4bb_1 _31267_ (.A(_01378_),
    .B(_01384_),
    .C_N(_02981_),
    .D_N(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__a2bb2o_1 _31268_ (.A1_N(_01378_),
    .A2_N(_01384_),
    .B1(_02981_),
    .B2(_02982_),
    .X(_02984_));
 sky130_fd_sc_hd__a21boi_2 _31269_ (.A1(_01390_),
    .A2(_01394_),
    .B1_N(_01391_),
    .Y(_02985_));
 sky130_fd_sc_hd__nand2_1 _31270_ (.A(_02981_),
    .B(_02982_),
    .Y(_02987_));
 sky130_fd_sc_hd__a21oi_2 _31271_ (.A1(_25176_),
    .A2(_01380_),
    .B1(_01378_),
    .Y(_02988_));
 sky130_fd_sc_hd__a21oi_2 _31272_ (.A1(_02987_),
    .A2(_02988_),
    .B1(_02985_),
    .Y(_02989_));
 sky130_fd_sc_hd__or2_1 _31273_ (.A(_02988_),
    .B(_02987_),
    .X(_02990_));
 sky130_fd_sc_hd__a32o_1 _31274_ (.A1(_02983_),
    .A2(_02984_),
    .A3(_02985_),
    .B1(_02989_),
    .B2(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__o22ai_4 _31275_ (.A1(_01395_),
    .A2(_01398_),
    .B1(_01400_),
    .B2(_25205_),
    .Y(_02992_));
 sky130_fd_sc_hd__xnor2_2 _31276_ (.A(_02991_),
    .B(_02992_),
    .Y(_00006_));
 sky130_fd_sc_hd__o21ai_1 _31277_ (.A1(_02939_),
    .A2(_02940_),
    .B1(_02932_),
    .Y(_02993_));
 sky130_fd_sc_hd__a32oi_2 _31278_ (.A1(_02060_),
    .A2(_02061_),
    .A3(_02064_),
    .B1(_01474_),
    .B2(_00450_),
    .Y(_02994_));
 sky130_fd_sc_hd__buf_1 _31279_ (.A(\delay_line[17][12] ),
    .X(_02995_));
 sky130_fd_sc_hd__or2b_1 _31280_ (.A(_02995_),
    .B_N(_01409_),
    .X(_02997_));
 sky130_fd_sc_hd__or3b_1 _31281_ (.A(_01417_),
    .B(_01421_),
    .C_N(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__o21ai_1 _31282_ (.A1(_01418_),
    .A2(_02997_),
    .B1(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__xor2_2 _31283_ (.A(_25251_),
    .B(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__buf_1 _31284_ (.A(\delay_line[17][13] ),
    .X(_03001_));
 sky130_fd_sc_hd__nor2_1 _31285_ (.A(_02995_),
    .B(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__and2_1 _31286_ (.A(_02995_),
    .B(\delay_line[17][13] ),
    .X(_03003_));
 sky130_fd_sc_hd__or2_1 _31287_ (.A(_03002_),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_2 _31288_ (.A(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__nor2_1 _31289_ (.A(_19815_),
    .B(_19800_),
    .Y(_03006_));
 sky130_fd_sc_hd__and2_1 _31290_ (.A(_19800_),
    .B(_19815_),
    .X(_03008_));
 sky130_fd_sc_hd__nor2_1 _31291_ (.A(_03006_),
    .B(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__xor2_2 _31292_ (.A(_03005_),
    .B(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_2 _31293_ (.A(_23707_),
    .X(_03011_));
 sky130_fd_sc_hd__a21oi_1 _31294_ (.A1(_23563_),
    .A2(_23685_),
    .B1(_23684_),
    .Y(_03012_));
 sky130_fd_sc_hd__nor2_1 _31295_ (.A(_03012_),
    .B(_23689_),
    .Y(_03013_));
 sky130_fd_sc_hd__and2_1 _31296_ (.A(_23689_),
    .B(_03012_),
    .X(_03014_));
 sky130_fd_sc_hd__nor3_2 _31297_ (.A(_03011_),
    .B(_03013_),
    .C(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__o21a_1 _31298_ (.A1(_03013_),
    .A2(_03014_),
    .B1(_03011_),
    .X(_03016_));
 sky130_fd_sc_hd__nor2_1 _31299_ (.A(_01425_),
    .B(_01427_),
    .Y(_03017_));
 sky130_fd_sc_hd__o21a_1 _31300_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_03017_),
    .X(_03019_));
 sky130_fd_sc_hd__or3_1 _31301_ (.A(_03017_),
    .B(_03015_),
    .C(_03016_),
    .X(_03020_));
 sky130_fd_sc_hd__and2b_1 _31302_ (.A_N(_03019_),
    .B(_03020_),
    .X(_03021_));
 sky130_fd_sc_hd__xor2_1 _31303_ (.A(_03010_),
    .B(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__o311a_1 _31304_ (.A1(_01419_),
    .A2(net204),
    .A3(_01433_),
    .B1(_01432_),
    .C1(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__a21oi_2 _31305_ (.A1(_01432_),
    .A2(_01434_),
    .B1(_03022_),
    .Y(_03024_));
 sky130_fd_sc_hd__nor2_1 _31306_ (.A(_03023_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__nor2_1 _31307_ (.A(_03000_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__and2_1 _31308_ (.A(_03025_),
    .B(_03000_),
    .X(_03027_));
 sky130_fd_sc_hd__or2_1 _31309_ (.A(_03026_),
    .B(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31310_ (.A(_01444_),
    .X(_03030_));
 sky130_fd_sc_hd__nor2_2 _31311_ (.A(_01444_),
    .B(net364),
    .Y(_03031_));
 sky130_fd_sc_hd__and2_1 _31312_ (.A(_01444_),
    .B(\delay_line[20][13] ),
    .X(_03032_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31313_ (.A(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__o2bb2a_1 _31314_ (.A1_N(_01443_),
    .A2_N(_03030_),
    .B1(_03031_),
    .B2(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__nor2_1 _31315_ (.A(_03031_),
    .B(_03032_),
    .Y(_03035_));
 sky130_fd_sc_hd__and3_1 _31316_ (.A(_01443_),
    .B(_03030_),
    .C(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__xnor2_2 _31317_ (.A(_23558_),
    .B(_25220_),
    .Y(_03037_));
 sky130_fd_sc_hd__nor3_2 _31318_ (.A(_03034_),
    .B(_03036_),
    .C(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__o21a_1 _31319_ (.A1(_03034_),
    .A2(_03036_),
    .B1(_03037_),
    .X(_03039_));
 sky130_fd_sc_hd__or4_1 _31320_ (.A(_17898_),
    .B(_04601_),
    .C(_03038_),
    .D(_03039_),
    .X(_03041_));
 sky130_fd_sc_hd__o22ai_2 _31321_ (.A1(_02038_),
    .A2(_22781_),
    .B1(_03039_),
    .B2(_03038_),
    .Y(_03042_));
 sky130_fd_sc_hd__o211a_1 _31322_ (.A1(_01449_),
    .A2(_01453_),
    .B1(_03041_),
    .C1(_03042_),
    .X(_03043_));
 sky130_fd_sc_hd__a221oi_2 _31323_ (.A1(_25219_),
    .A2(_01448_),
    .B1(_03041_),
    .B2(_03042_),
    .C1(_01453_),
    .Y(_03044_));
 sky130_fd_sc_hd__a211o_1 _31324_ (.A1(_02038_),
    .A2(_10372_),
    .B1(_02039_),
    .C1(_02046_),
    .X(_03045_));
 sky130_fd_sc_hd__o31a_1 _31325_ (.A1(_00438_),
    .A2(_02042_),
    .A3(_02043_),
    .B1(_03045_),
    .X(_03046_));
 sky130_fd_sc_hd__o21a_1 _31326_ (.A1(_03043_),
    .A2(_03044_),
    .B1(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__nor3_2 _31327_ (.A(_03046_),
    .B(_03043_),
    .C(_03044_),
    .Y(_03048_));
 sky130_fd_sc_hd__o21ai_1 _31328_ (.A1(_03047_),
    .A2(_03048_),
    .B1(_01455_),
    .Y(_03049_));
 sky130_fd_sc_hd__nor4_1 _31329_ (.A(_15427_),
    .B(_24282_),
    .C(_01453_),
    .D(_01454_),
    .Y(_03050_));
 sky130_fd_sc_hd__nor2_1 _31330_ (.A(_03047_),
    .B(_03048_),
    .Y(_03052_));
 sky130_fd_sc_hd__o21a_1 _31331_ (.A1(_03050_),
    .A2(_01458_),
    .B1(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__o21bai_1 _31332_ (.A1(_01458_),
    .A2(_03049_),
    .B1_N(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__and3_1 _31333_ (.A(_01460_),
    .B(_01462_),
    .C(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__a21o_1 _31334_ (.A1(_01460_),
    .A2(_01462_),
    .B1(_03054_),
    .X(_03056_));
 sky130_fd_sc_hd__and2b_1 _31335_ (.A_N(_03055_),
    .B(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__xnor2_1 _31336_ (.A(_03028_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__o21ai_1 _31337_ (.A1(_02933_),
    .A2(_02994_),
    .B1(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__a211o_1 _31338_ (.A1(_01475_),
    .A2(_02065_),
    .B1(_03058_),
    .C1(_02933_),
    .X(_03060_));
 sky130_fd_sc_hd__or2b_1 _31339_ (.A(_01441_),
    .B_N(_01465_),
    .X(_03061_));
 sky130_fd_sc_hd__o21ai_2 _31340_ (.A1(_01442_),
    .A2(_01464_),
    .B1(_03061_),
    .Y(_03063_));
 sky130_fd_sc_hd__a21oi_2 _31341_ (.A1(_03059_),
    .A2(_03060_),
    .B1(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__and3_2 _31342_ (.A(_03059_),
    .B(_03060_),
    .C(_03063_),
    .X(_03065_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31343_ (.A(\delay_line[23][13] ),
    .X(_03066_));
 sky130_fd_sc_hd__nor2_2 _31344_ (.A(net347),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__and2_4 _31345_ (.A(net347),
    .B(\delay_line[23][13] ),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_2 _31346_ (.A(_01980_),
    .X(_03069_));
 sky130_fd_sc_hd__nand2_2 _31347_ (.A(_01986_),
    .B(_01988_),
    .Y(_03070_));
 sky130_fd_sc_hd__o2bb2ai_2 _31348_ (.A1_N(_00408_),
    .A2_N(_24224_),
    .B1(_00402_),
    .B2(_00404_),
    .Y(_03071_));
 sky130_fd_sc_hd__o22ai_1 _31349_ (.A1(_03069_),
    .A2(_03070_),
    .B1(_01990_),
    .B2(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__nor2_1 _31350_ (.A(_01524_),
    .B(_01969_),
    .Y(_03074_));
 sky130_fd_sc_hd__and2_2 _31351_ (.A(_01515_),
    .B(_01483_),
    .X(_03075_));
 sky130_fd_sc_hd__nand2_1 _31352_ (.A(_01513_),
    .B(_01485_),
    .Y(_03076_));
 sky130_fd_sc_hd__o21a_1 _31353_ (.A1(_01484_),
    .A2(_01514_),
    .B1(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__o21ba_1 _31354_ (.A1(_01505_),
    .A2(_01503_),
    .B1_N(_01504_),
    .X(_03078_));
 sky130_fd_sc_hd__and2_1 _31355_ (.A(_01857_),
    .B(_01858_),
    .X(_03079_));
 sky130_fd_sc_hd__and2b_2 _31356_ (.A_N(_22235_),
    .B(_00324_),
    .X(_03080_));
 sky130_fd_sc_hd__o21bai_1 _31357_ (.A1(_01496_),
    .A2(_01497_),
    .B1_N(_00321_),
    .Y(_03081_));
 sky130_fd_sc_hd__nor2_1 _31358_ (.A(_01494_),
    .B(net447),
    .Y(_03082_));
 sky130_fd_sc_hd__nand2_1 _31359_ (.A(_01494_),
    .B(net447),
    .Y(_03083_));
 sky130_fd_sc_hd__nand3b_2 _31360_ (.A_N(_03082_),
    .B(_03083_),
    .C(net440),
    .Y(_03085_));
 sky130_fd_sc_hd__and2_1 _31361_ (.A(_01494_),
    .B(net447),
    .X(_03086_));
 sky130_fd_sc_hd__o21bai_1 _31362_ (.A1(_03082_),
    .A2(_03086_),
    .B1_N(net440),
    .Y(_03087_));
 sky130_fd_sc_hd__and3_1 _31363_ (.A(_01497_),
    .B(_03085_),
    .C(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__a21oi_1 _31364_ (.A1(_03085_),
    .A2(_03087_),
    .B1(_01497_),
    .Y(_03089_));
 sky130_fd_sc_hd__buf_1 _31365_ (.A(net448),
    .X(_03090_));
 sky130_fd_sc_hd__buf_1 _31366_ (.A(_01492_),
    .X(_03091_));
 sky130_fd_sc_hd__a21oi_1 _31367_ (.A1(_03090_),
    .A2(_03091_),
    .B1(_03080_),
    .Y(_03092_));
 sky130_fd_sc_hd__and3_1 _31368_ (.A(_03090_),
    .B(_03080_),
    .C(_03091_),
    .X(_03093_));
 sky130_fd_sc_hd__o22ai_2 _31369_ (.A1(_03088_),
    .A2(_03089_),
    .B1(_03092_),
    .B2(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__or4_2 _31370_ (.A(_03088_),
    .B(_03089_),
    .C(_03092_),
    .D(_03093_),
    .X(_03096_));
 sky130_fd_sc_hd__a221o_1 _31371_ (.A1(_01491_),
    .A2(_03081_),
    .B1(_03094_),
    .B2(_03096_),
    .C1(net271),
    .X(_03097_));
 sky130_fd_sc_hd__a21o_1 _31372_ (.A1(_01491_),
    .A2(_03081_),
    .B1(net271),
    .X(_03098_));
 sky130_fd_sc_hd__nand3_2 _31373_ (.A(_03098_),
    .B(_03094_),
    .C(_03096_),
    .Y(_03099_));
 sky130_fd_sc_hd__or2b_1 _31374_ (.A(_03090_),
    .B_N(_00324_),
    .X(_03100_));
 sky130_fd_sc_hd__o2111ai_4 _31375_ (.A1(_22239_),
    .A2(_03080_),
    .B1(_03097_),
    .C1(_03099_),
    .D1(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__a21o_1 _31376_ (.A1(_24156_),
    .A2(_24157_),
    .B1(_03080_),
    .X(_03102_));
 sky130_fd_sc_hd__a22o_1 _31377_ (.A1(_03100_),
    .A2(_03102_),
    .B1(_03097_),
    .B2(_03099_),
    .X(_03103_));
 sky130_fd_sc_hd__o211ai_1 _31378_ (.A1(_01855_),
    .A2(_03079_),
    .B1(_03101_),
    .C1(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__a221o_1 _31379_ (.A1(_01858_),
    .A2(_01857_),
    .B1(_03103_),
    .B2(_03101_),
    .C1(_01855_),
    .X(_03105_));
 sky130_fd_sc_hd__nand2_1 _31380_ (.A(_03104_),
    .B(_03105_),
    .Y(_03107_));
 sky130_fd_sc_hd__xnor2_2 _31381_ (.A(_03078_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__o21a_1 _31382_ (.A1(_01859_),
    .A2(_01904_),
    .B1(_01903_),
    .X(_03109_));
 sky130_fd_sc_hd__xnor2_1 _31383_ (.A(_03108_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__o21ai_1 _31384_ (.A1(_01486_),
    .A2(_01511_),
    .B1(_01510_),
    .Y(_03111_));
 sky130_fd_sc_hd__or2b_1 _31385_ (.A(_03110_),
    .B_N(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__o211ai_1 _31386_ (.A1(_01511_),
    .A2(_01486_),
    .B1(_01510_),
    .C1(_03110_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2_1 _31387_ (.A(_03112_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__nor2_1 _31388_ (.A(_03077_),
    .B(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__o211a_1 _31389_ (.A1(_01514_),
    .A2(_01484_),
    .B1(_03076_),
    .C1(_03114_),
    .X(_03116_));
 sky130_fd_sc_hd__o21ai_1 _31390_ (.A1(net136),
    .A2(_01948_),
    .B1(_01946_),
    .Y(_03118_));
 sky130_fd_sc_hd__o211ai_1 _31391_ (.A1(_03115_),
    .A2(_03116_),
    .B1(_01947_),
    .C1(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__a211o_1 _31392_ (.A1(_01947_),
    .A2(_03118_),
    .B1(_03115_),
    .C1(_03116_),
    .X(_03120_));
 sky130_fd_sc_hd__nand2_1 _31393_ (.A(_03119_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__xnor2_1 _31394_ (.A(_03075_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__o21ai_1 _31395_ (.A1(_02491_),
    .A2(_17982_),
    .B1(_01533_),
    .Y(_03123_));
 sky130_fd_sc_hd__nor2_1 _31396_ (.A(_01649_),
    .B(net256),
    .Y(_03124_));
 sky130_fd_sc_hd__buf_2 _31397_ (.A(net401),
    .X(_03125_));
 sky130_fd_sc_hd__nand2_1 _31398_ (.A(net402),
    .B(net401),
    .Y(_03126_));
 sky130_fd_sc_hd__or2_1 _31399_ (.A(\delay_line[12][11] ),
    .B(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__o21a_1 _31400_ (.A1(_01527_),
    .A2(_03125_),
    .B1(_03127_),
    .X(_03129_));
 sky130_fd_sc_hd__inv_2 _31401_ (.A(net402),
    .Y(_03130_));
 sky130_fd_sc_hd__clkbuf_2 _31402_ (.A(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__or3b_1 _31403_ (.A(_03125_),
    .B(_03131_),
    .C_N(_00121_),
    .X(_03132_));
 sky130_fd_sc_hd__and3_1 _31404_ (.A(_25372_),
    .B(_03129_),
    .C(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__a21oi_1 _31405_ (.A1(_03129_),
    .A2(_03132_),
    .B1(_25372_),
    .Y(_03134_));
 sky130_fd_sc_hd__nor3b_1 _31406_ (.A(_03133_),
    .B(_03134_),
    .C_N(_00099_),
    .Y(_03135_));
 sky130_fd_sc_hd__o21ba_1 _31407_ (.A1(_03133_),
    .A2(_03134_),
    .B1_N(_00099_),
    .X(_03136_));
 sky130_fd_sc_hd__nor3_1 _31408_ (.A(_03124_),
    .B(_03135_),
    .C(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__o21a_1 _31409_ (.A1(_03135_),
    .A2(_03136_),
    .B1(_03124_),
    .X(_03138_));
 sky130_fd_sc_hd__or2_1 _31410_ (.A(_03137_),
    .B(_03138_),
    .X(_03140_));
 sky130_fd_sc_hd__a21oi_1 _31411_ (.A1(_00130_),
    .A2(_03123_),
    .B1(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__and3_1 _31412_ (.A(_03140_),
    .B(_00130_),
    .C(_03123_),
    .X(_03142_));
 sky130_fd_sc_hd__o21ai_2 _31413_ (.A1(_01636_),
    .A2(_01625_),
    .B1(_01638_),
    .Y(_03143_));
 sky130_fd_sc_hd__nor2_1 _31414_ (.A(_00075_),
    .B(\delay_line[13][13] ),
    .Y(_03144_));
 sky130_fd_sc_hd__buf_1 _31415_ (.A(\delay_line[13][13] ),
    .X(_03145_));
 sky130_fd_sc_hd__nand2_1 _31416_ (.A(_00075_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__and4b_2 _31417_ (.A_N(_03144_),
    .B(_01547_),
    .C(_22343_),
    .D(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__buf_2 _31418_ (.A(_01547_),
    .X(_03148_));
 sky130_fd_sc_hd__and2_1 _31419_ (.A(_00075_),
    .B(_03145_),
    .X(_03149_));
 sky130_fd_sc_hd__o2bb2a_1 _31420_ (.A1_N(_22343_),
    .A2_N(_03148_),
    .B1(_03149_),
    .B2(_03144_),
    .X(_03151_));
 sky130_fd_sc_hd__or4_2 _31421_ (.A(_01557_),
    .B(_25431_),
    .C(_01554_),
    .D(_25437_),
    .X(_03152_));
 sky130_fd_sc_hd__xnor2_4 _31422_ (.A(_22308_),
    .B(net410),
    .Y(_03153_));
 sky130_fd_sc_hd__o21a_1 _31423_ (.A1(_21718_),
    .A2(\delay_line[11][10] ),
    .B1(_01558_),
    .X(_03154_));
 sky130_fd_sc_hd__a211o_1 _31424_ (.A1(_21728_),
    .A2(_01555_),
    .B1(_03153_),
    .C1(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__o21ai_1 _31425_ (.A1(_01554_),
    .A2(_03154_),
    .B1(_03153_),
    .Y(_03156_));
 sky130_fd_sc_hd__nand2_1 _31426_ (.A(_03155_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__a21oi_2 _31427_ (.A1(_01599_),
    .A2(_03152_),
    .B1(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__o211a_1 _31428_ (.A1(_01564_),
    .A2(_01570_),
    .B1(_03157_),
    .C1(_03152_),
    .X(_03159_));
 sky130_fd_sc_hd__clkbuf_2 _31429_ (.A(\delay_line[4][10] ),
    .X(_03160_));
 sky130_fd_sc_hd__and2b_1 _31430_ (.A_N(_25416_),
    .B(_03160_),
    .X(_03162_));
 sky130_fd_sc_hd__and2b_1 _31431_ (.A_N(\delay_line[4][10] ),
    .B(\delay_line[4][8] ),
    .X(_03163_));
 sky130_fd_sc_hd__nand2_1 _31432_ (.A(_01573_),
    .B(_01579_),
    .Y(_03164_));
 sky130_fd_sc_hd__clkbuf_2 _31433_ (.A(_01575_),
    .X(_03165_));
 sky130_fd_sc_hd__a2bb2o_1 _31434_ (.A1_N(_03162_),
    .A2_N(_03163_),
    .B1(_03164_),
    .B2(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__nor2_1 _31435_ (.A(_03162_),
    .B(_03163_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand3_2 _31436_ (.A(_03165_),
    .B(_03164_),
    .C(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__clkbuf_2 _31437_ (.A(\delay_line[4][9] ),
    .X(_03169_));
 sky130_fd_sc_hd__and2_1 _31438_ (.A(_25417_),
    .B(_25418_),
    .X(_03170_));
 sky130_fd_sc_hd__a32oi_4 _31439_ (.A1(_03169_),
    .A2(_25419_),
    .A3(_03170_),
    .B1(_01581_),
    .B2(_01582_),
    .Y(_03171_));
 sky130_fd_sc_hd__a22oi_4 _31440_ (.A1(_03166_),
    .A2(_03168_),
    .B1(_01604_),
    .B2(_03171_),
    .Y(_03173_));
 sky130_fd_sc_hd__a21oi_2 _31441_ (.A1(_03165_),
    .A2(_03164_),
    .B1(_03167_),
    .Y(_03174_));
 sky130_fd_sc_hd__and3_1 _31442_ (.A(_03165_),
    .B(_03164_),
    .C(_03167_),
    .X(_03175_));
 sky130_fd_sc_hd__nor2_1 _31443_ (.A(_03174_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__inv_2 _31444_ (.A(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__a32o_2 _31445_ (.A1(_03169_),
    .A2(_25419_),
    .A3(_03170_),
    .B1(_01581_),
    .B2(_01582_),
    .X(_03178_));
 sky130_fd_sc_hd__a21oi_4 _31446_ (.A1(_25411_),
    .A2(_25415_),
    .B1(_01586_),
    .Y(_03179_));
 sky130_fd_sc_hd__nor3_2 _31447_ (.A(_03177_),
    .B(_03178_),
    .C(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__o22ai_4 _31448_ (.A1(_03158_),
    .A2(_03159_),
    .B1(_03173_),
    .B2(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__a21o_1 _31449_ (.A1(_01599_),
    .A2(_03152_),
    .B1(_03157_),
    .X(_03182_));
 sky130_fd_sc_hd__o211ai_2 _31450_ (.A1(_01564_),
    .A2(_01570_),
    .B1(_03157_),
    .C1(_03152_),
    .Y(_03184_));
 sky130_fd_sc_hd__o22ai_4 _31451_ (.A1(_03174_),
    .A2(_03175_),
    .B1(_03178_),
    .B2(_03179_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand3_1 _31452_ (.A(_01604_),
    .B(_03176_),
    .C(_03171_),
    .Y(_03186_));
 sky130_fd_sc_hd__nand4_4 _31453_ (.A(_03182_),
    .B(_03184_),
    .C(_03185_),
    .D(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__a21oi_4 _31454_ (.A1(_03181_),
    .A2(_03187_),
    .B1(net453),
    .Y(_03188_));
 sky130_fd_sc_hd__nand3_2 _31455_ (.A(_03181_),
    .B(_03187_),
    .C(net453),
    .Y(_03189_));
 sky130_fd_sc_hd__o21ai_2 _31456_ (.A1(_01602_),
    .A2(_01627_),
    .B1(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__clkbuf_4 _31457_ (.A(\delay_line[0][12] ),
    .X(_03191_));
 sky130_fd_sc_hd__and3_1 _31458_ (.A(_03181_),
    .B(_03187_),
    .C(net453),
    .X(_03192_));
 sky130_fd_sc_hd__a21oi_1 _31459_ (.A1(_01626_),
    .A2(_01609_),
    .B1(_01590_),
    .Y(_03193_));
 sky130_fd_sc_hd__o21bai_4 _31460_ (.A1(_03188_),
    .A2(_03192_),
    .B1_N(_03193_),
    .Y(_03195_));
 sky130_fd_sc_hd__o211ai_4 _31461_ (.A1(_03188_),
    .A2(_03190_),
    .B1(_03191_),
    .C1(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__nor2_1 _31462_ (.A(_03188_),
    .B(_03190_),
    .Y(_03197_));
 sky130_fd_sc_hd__clkbuf_2 _31463_ (.A(net453),
    .X(_03198_));
 sky130_fd_sc_hd__a21o_1 _31464_ (.A1(_03181_),
    .A2(_03187_),
    .B1(_03198_),
    .X(_03199_));
 sky130_fd_sc_hd__a21oi_2 _31465_ (.A1(_03199_),
    .A2(_03189_),
    .B1(_03193_),
    .Y(_03200_));
 sky130_fd_sc_hd__o21bai_1 _31466_ (.A1(_03197_),
    .A2(_03200_),
    .B1_N(_03191_),
    .Y(_03201_));
 sky130_fd_sc_hd__a21o_1 _31467_ (.A1(_01620_),
    .A2(_01630_),
    .B1(_01616_),
    .X(_03202_));
 sky130_fd_sc_hd__a21oi_2 _31468_ (.A1(_03196_),
    .A2(_03201_),
    .B1(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__o2111ai_4 _31469_ (.A1(_03191_),
    .A2(_01602_),
    .B1(_03199_),
    .C1(_03189_),
    .D1(_01607_),
    .Y(_03204_));
 sky130_fd_sc_hd__buf_2 _31470_ (.A(_03191_),
    .X(_03206_));
 sky130_fd_sc_hd__a21oi_4 _31471_ (.A1(_03204_),
    .A2(_03195_),
    .B1(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__nand2_2 _31472_ (.A(_03202_),
    .B(_03196_),
    .Y(_03208_));
 sky130_fd_sc_hd__nor2_2 _31473_ (.A(_03207_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__o22ai_4 _31474_ (.A1(_03147_),
    .A2(_03151_),
    .B1(_03203_),
    .B2(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__nor2_1 _31475_ (.A(_03147_),
    .B(_03151_),
    .Y(_03211_));
 sky130_fd_sc_hd__a21o_1 _31476_ (.A1(_03196_),
    .A2(_03201_),
    .B1(_03202_),
    .X(_03212_));
 sky130_fd_sc_hd__o211ai_4 _31477_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03211_),
    .C1(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__nand3_2 _31478_ (.A(_03143_),
    .B(_03210_),
    .C(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__o21ai_1 _31479_ (.A1(_03203_),
    .A2(_03209_),
    .B1(_03211_),
    .Y(_03215_));
 sky130_fd_sc_hd__o31a_1 _31480_ (.A1(_01550_),
    .A2(_01552_),
    .A3(_01625_),
    .B1(_01638_),
    .X(_03217_));
 sky130_fd_sc_hd__o221ai_1 _31481_ (.A1(_03147_),
    .A2(_03151_),
    .B1(_03207_),
    .B2(_03208_),
    .C1(_03212_),
    .Y(_03218_));
 sky130_fd_sc_hd__nand3_1 _31482_ (.A(_03215_),
    .B(_03217_),
    .C(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__clkbuf_2 _31483_ (.A(_18918_),
    .X(_03220_));
 sky130_fd_sc_hd__buf_2 _31484_ (.A(_00096_),
    .X(_03221_));
 sky130_fd_sc_hd__xnor2_2 _31485_ (.A(_20046_),
    .B(\delay_line[13][11] ),
    .Y(_03222_));
 sky130_fd_sc_hd__nor2_1 _31486_ (.A(_23811_),
    .B(_01635_),
    .Y(_03223_));
 sky130_fd_sc_hd__a221oi_4 _31487_ (.A1(_03220_),
    .A2(_03221_),
    .B1(_01635_),
    .B2(_03222_),
    .C1(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__a21oi_1 _31488_ (.A1(_01635_),
    .A2(_03222_),
    .B1(_03223_),
    .Y(_03225_));
 sky130_fd_sc_hd__nor2_1 _31489_ (.A(_01647_),
    .B(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__o2bb2ai_1 _31490_ (.A1_N(_03214_),
    .A2_N(_03219_),
    .B1(_03224_),
    .B2(_03226_),
    .Y(_03228_));
 sky130_fd_sc_hd__nor2_1 _31491_ (.A(_01657_),
    .B(_01658_),
    .Y(_03229_));
 sky130_fd_sc_hd__a32oi_1 _31492_ (.A1(_01544_),
    .A2(_01634_),
    .A3(_01639_),
    .B1(_01659_),
    .B2(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__and3_1 _31493_ (.A(_03220_),
    .B(_03221_),
    .C(_03225_),
    .X(_03231_));
 sky130_fd_sc_hd__a21oi_1 _31494_ (.A1(_03220_),
    .A2(_03221_),
    .B1(_03225_),
    .Y(_03232_));
 sky130_fd_sc_hd__clkbuf_2 _31495_ (.A(_03219_),
    .X(_03233_));
 sky130_fd_sc_hd__o211ai_1 _31496_ (.A1(_03231_),
    .A2(_03232_),
    .B1(_03214_),
    .C1(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand3_1 _31497_ (.A(_03228_),
    .B(_03230_),
    .C(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__buf_4 _31498_ (.A(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__o21ai_2 _31499_ (.A1(_03141_),
    .A2(_03142_),
    .B1(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__a32o_2 _31500_ (.A1(_01544_),
    .A2(_01634_),
    .A3(_01639_),
    .B1(_01659_),
    .B2(_03229_),
    .X(_03239_));
 sky130_fd_sc_hd__o2bb2ai_2 _31501_ (.A1_N(_03214_),
    .A2_N(_03233_),
    .B1(_03231_),
    .B2(_03232_),
    .Y(_03240_));
 sky130_fd_sc_hd__o211ai_4 _31502_ (.A1(_03224_),
    .A2(_03226_),
    .B1(_03214_),
    .C1(_03233_),
    .Y(_03241_));
 sky130_fd_sc_hd__and3_1 _31503_ (.A(_03239_),
    .B(_03240_),
    .C(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__nor2_1 _31504_ (.A(_01672_),
    .B(_01673_),
    .Y(_03243_));
 sky130_fd_sc_hd__a32o_1 _31505_ (.A1(_01664_),
    .A2(_01665_),
    .A3(_01667_),
    .B1(_01662_),
    .B2(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__nand3_2 _31506_ (.A(_03239_),
    .B(_03240_),
    .C(_03241_),
    .Y(_03245_));
 sky130_fd_sc_hd__and2_1 _31507_ (.A(_03123_),
    .B(_00130_),
    .X(_03246_));
 sky130_fd_sc_hd__inv_2 _31508_ (.A(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__nor2_2 _31509_ (.A(_03247_),
    .B(_03140_),
    .Y(_03248_));
 sky130_fd_sc_hd__and2_1 _31510_ (.A(_03247_),
    .B(_03140_),
    .X(_03250_));
 sky130_fd_sc_hd__o2bb2ai_2 _31511_ (.A1_N(_03245_),
    .A2_N(_03236_),
    .B1(_03248_),
    .B2(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__o211ai_4 _31512_ (.A1(_03237_),
    .A2(_03242_),
    .B1(_03244_),
    .C1(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__o2bb2ai_1 _31513_ (.A1_N(_03245_),
    .A2_N(_03235_),
    .B1(_03141_),
    .B2(_03142_),
    .Y(_03253_));
 sky130_fd_sc_hd__a21oi_1 _31514_ (.A1(_01662_),
    .A2(_03243_),
    .B1(_01668_),
    .Y(_03254_));
 sky130_fd_sc_hd__o211ai_1 _31515_ (.A1(_03248_),
    .A2(_03250_),
    .B1(_03245_),
    .C1(_03236_),
    .Y(_03255_));
 sky130_fd_sc_hd__nand3_1 _31516_ (.A(_03253_),
    .B(_03254_),
    .C(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__clkbuf_2 _31517_ (.A(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__a21o_1 _31518_ (.A1(_01671_),
    .A2(_01539_),
    .B1(_01538_),
    .X(_03258_));
 sky130_fd_sc_hd__or2b_1 _31519_ (.A(_17918_),
    .B_N(net416),
    .X(_03259_));
 sky130_fd_sc_hd__or2b_1 _31520_ (.A(net416),
    .B_N(_17918_),
    .X(_03261_));
 sky130_fd_sc_hd__nand4_1 _31521_ (.A(_03259_),
    .B(_03261_),
    .C(_19964_),
    .D(_25392_),
    .Y(_03262_));
 sky130_fd_sc_hd__a22o_1 _31522_ (.A1(_22447_),
    .A2(_25392_),
    .B1(_03259_),
    .B2(_03261_),
    .X(_03263_));
 sky130_fd_sc_hd__and3b_1 _31523_ (.A_N(_01683_),
    .B(_03262_),
    .C(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__clkbuf_2 _31524_ (.A(_01682_),
    .X(_03265_));
 sky130_fd_sc_hd__o2bb2a_1 _31525_ (.A1_N(_03262_),
    .A2_N(_03263_),
    .B1(_25396_),
    .B2(_03265_),
    .X(_03266_));
 sky130_fd_sc_hd__nor2_1 _31526_ (.A(_19956_),
    .B(_21800_),
    .Y(_03267_));
 sky130_fd_sc_hd__and2_1 _31527_ (.A(net412),
    .B(_21800_),
    .X(_03268_));
 sky130_fd_sc_hd__o21ai_1 _31528_ (.A1(_03267_),
    .A2(_03268_),
    .B1(_23762_),
    .Y(_03269_));
 sky130_fd_sc_hd__or3_1 _31529_ (.A(_23758_),
    .B(_03267_),
    .C(_03268_),
    .X(_03270_));
 sky130_fd_sc_hd__and3b_1 _31530_ (.A_N(_01693_),
    .B(_03269_),
    .C(_03270_),
    .X(_03272_));
 sky130_fd_sc_hd__a32oi_2 _31531_ (.A1(_01694_),
    .A2(_01690_),
    .A3(_01691_),
    .B1(_03269_),
    .B2(_03270_),
    .Y(_03273_));
 sky130_fd_sc_hd__or4_1 _31532_ (.A(_03264_),
    .B(_03266_),
    .C(_03272_),
    .D(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__o22ai_2 _31533_ (.A1(_03264_),
    .A2(_03266_),
    .B1(_03272_),
    .B2(_03273_),
    .Y(_03275_));
 sky130_fd_sc_hd__and3_1 _31534_ (.A(_03130_),
    .B(_01526_),
    .C(_23800_),
    .X(_03276_));
 sky130_fd_sc_hd__a31o_1 _31535_ (.A1(_01528_),
    .A2(_01530_),
    .A3(_21805_),
    .B1(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__and2_1 _31536_ (.A(_20060_),
    .B(net411),
    .X(_03278_));
 sky130_fd_sc_hd__nor2_1 _31537_ (.A(_20062_),
    .B(net411),
    .Y(_03279_));
 sky130_fd_sc_hd__or3b_2 _31538_ (.A(_03278_),
    .B(_03279_),
    .C_N(_01705_),
    .X(_03280_));
 sky130_fd_sc_hd__buf_1 _31539_ (.A(\delay_line[10][12] ),
    .X(_03281_));
 sky130_fd_sc_hd__clkbuf_2 _31540_ (.A(_03281_),
    .X(_03283_));
 sky130_fd_sc_hd__a2bb2o_1 _31541_ (.A1_N(_03278_),
    .A2_N(_03279_),
    .B1(_18985_),
    .B2(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__and3_1 _31542_ (.A(_03277_),
    .B(_03280_),
    .C(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__a21oi_1 _31543_ (.A1(_03280_),
    .A2(_03284_),
    .B1(_03277_),
    .Y(_03286_));
 sky130_fd_sc_hd__o21ai_1 _31544_ (.A1(_03285_),
    .A2(_03286_),
    .B1(_01711_),
    .Y(_03287_));
 sky130_fd_sc_hd__or3_1 _31545_ (.A(_03286_),
    .B(_01711_),
    .C(_03285_),
    .X(_03288_));
 sky130_fd_sc_hd__or2b_1 _31546_ (.A(_01709_),
    .B_N(_01713_),
    .X(_03289_));
 sky130_fd_sc_hd__a21o_1 _31547_ (.A1(_03287_),
    .A2(_03288_),
    .B1(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__nand2_1 _31548_ (.A(_03289_),
    .B(_03287_),
    .Y(_03291_));
 sky130_fd_sc_hd__and4_1 _31549_ (.A(_03274_),
    .B(_03275_),
    .C(_03290_),
    .D(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__a22oi_1 _31550_ (.A1(_03274_),
    .A2(_03275_),
    .B1(_03290_),
    .B2(_03291_),
    .Y(_03294_));
 sky130_fd_sc_hd__nor2_1 _31551_ (.A(_03292_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__xnor2_1 _31552_ (.A(_03258_),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__a31o_1 _31553_ (.A1(_01718_),
    .A2(_01700_),
    .A3(_01698_),
    .B1(_01717_),
    .X(_03297_));
 sky130_fd_sc_hd__nor2_1 _31554_ (.A(_03296_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__and2_1 _31555_ (.A(_03296_),
    .B(_03297_),
    .X(_03299_));
 sky130_fd_sc_hd__o2bb2ai_1 _31556_ (.A1_N(_03252_),
    .A2_N(_03257_),
    .B1(_03298_),
    .B2(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__inv_2 _31557_ (.A(_03297_),
    .Y(_03301_));
 sky130_fd_sc_hd__nor2_2 _31558_ (.A(_03301_),
    .B(_03296_),
    .Y(_03302_));
 sky130_fd_sc_hd__and2_1 _31559_ (.A(_03296_),
    .B(_03301_),
    .X(_03303_));
 sky130_fd_sc_hd__o211ai_2 _31560_ (.A1(_03302_),
    .A2(_03303_),
    .B1(_03252_),
    .C1(_03257_),
    .Y(_03305_));
 sky130_fd_sc_hd__a21oi_1 _31561_ (.A1(_01734_),
    .A2(_01824_),
    .B1(_01826_),
    .Y(_03306_));
 sky130_fd_sc_hd__nand3_4 _31562_ (.A(_03300_),
    .B(_03305_),
    .C(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__o21a_1 _31563_ (.A1(_01784_),
    .A2(_01814_),
    .B1(_01812_),
    .X(_03308_));
 sky130_fd_sc_hd__a21o_1 _31564_ (.A1(_01723_),
    .A2(_01722_),
    .B1(_01720_),
    .X(_03309_));
 sky130_fd_sc_hd__or2b_1 _31565_ (.A(_01696_),
    .B_N(_01698_),
    .X(_03310_));
 sky130_fd_sc_hd__buf_1 _31566_ (.A(net418),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_2 _31567_ (.A(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__or2_1 _31568_ (.A(_03311_),
    .B(net417),
    .X(_03313_));
 sky130_fd_sc_hd__nand2_2 _31569_ (.A(_03311_),
    .B(net417),
    .Y(_03314_));
 sky130_fd_sc_hd__a22o_1 _31570_ (.A1(_25341_),
    .A2(_03312_),
    .B1(_03313_),
    .B2(_03314_),
    .X(_03316_));
 sky130_fd_sc_hd__nand3_1 _31571_ (.A(_03265_),
    .B(_03312_),
    .C(_25341_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21o_1 _31572_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_01788_),
    .X(_03318_));
 sky130_fd_sc_hd__nand3_1 _31573_ (.A(_03316_),
    .B(_03317_),
    .C(_23969_),
    .Y(_03319_));
 sky130_fd_sc_hd__a211o_1 _31574_ (.A1(_03318_),
    .A2(_03319_),
    .B1(_01686_),
    .C1(_01687_),
    .X(_03320_));
 sky130_fd_sc_hd__o211ai_2 _31575_ (.A1(_01686_),
    .A2(_01687_),
    .B1(_03318_),
    .C1(_03319_),
    .Y(_03321_));
 sky130_fd_sc_hd__buf_2 _31576_ (.A(_03312_),
    .X(_03322_));
 sky130_fd_sc_hd__nor2_1 _31577_ (.A(_03322_),
    .B(_25339_),
    .Y(_03323_));
 sky130_fd_sc_hd__a221o_1 _31578_ (.A1(_01794_),
    .A2(_20123_),
    .B1(_03320_),
    .B2(_03321_),
    .C1(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__o211ai_2 _31579_ (.A1(_03323_),
    .A2(_01797_),
    .B1(_03321_),
    .C1(_03320_),
    .Y(_03325_));
 sky130_fd_sc_hd__nand3_2 _31580_ (.A(_03310_),
    .B(_03324_),
    .C(_03325_),
    .Y(_03327_));
 sky130_fd_sc_hd__a21o_1 _31581_ (.A1(_03324_),
    .A2(_03325_),
    .B1(_03310_),
    .X(_03328_));
 sky130_fd_sc_hd__a211o_1 _31582_ (.A1(_03327_),
    .A2(_03328_),
    .B1(_01799_),
    .C1(net231),
    .X(_03329_));
 sky130_fd_sc_hd__o211ai_4 _31583_ (.A1(_01799_),
    .A2(net231),
    .B1(_03327_),
    .C1(_03328_),
    .Y(_03330_));
 sky130_fd_sc_hd__a221oi_2 _31584_ (.A1(_01791_),
    .A2(_01803_),
    .B1(_03329_),
    .B2(_03330_),
    .C1(_01807_),
    .Y(_03331_));
 sky130_fd_sc_hd__inv_2 _31585_ (.A(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__o211ai_4 _31586_ (.A1(_01805_),
    .A2(_01807_),
    .B1(_03329_),
    .C1(_03330_),
    .Y(_03333_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31587_ (.A(\delay_line[7][13] ),
    .X(_03334_));
 sky130_fd_sc_hd__nor2b_1 _31588_ (.A(_18040_),
    .B_N(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__buf_1 _31589_ (.A(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_2 _31590_ (.A(_03334_),
    .X(_03338_));
 sky130_fd_sc_hd__and2b_1 _31591_ (.A_N(_03338_),
    .B(_18044_),
    .X(_03339_));
 sky130_fd_sc_hd__nor3_1 _31592_ (.A(_03336_),
    .B(_03339_),
    .C(_01748_),
    .Y(_03340_));
 sky130_fd_sc_hd__clkbuf_2 _31593_ (.A(_01744_),
    .X(_03341_));
 sky130_fd_sc_hd__o2bb2a_1 _31594_ (.A1_N(_11866_),
    .A2_N(_03341_),
    .B1(_03336_),
    .B2(_03339_),
    .X(_03342_));
 sky130_fd_sc_hd__o211a_1 _31595_ (.A1(_03340_),
    .A2(_03342_),
    .B1(_01766_),
    .C1(_01769_),
    .X(_03343_));
 sky130_fd_sc_hd__a211oi_2 _31596_ (.A1(_01766_),
    .A2(_01769_),
    .B1(_03340_),
    .C1(_03342_),
    .Y(_03344_));
 sky130_fd_sc_hd__nor3_2 _31597_ (.A(_01749_),
    .B(_03343_),
    .C(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__o21a_1 _31598_ (.A1(_03343_),
    .A2(_03344_),
    .B1(_01749_),
    .X(_03346_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31599_ (.A(_01771_),
    .X(_03347_));
 sky130_fd_sc_hd__clkbuf_2 _31600_ (.A(_03347_),
    .X(_03349_));
 sky130_fd_sc_hd__a31o_1 _31601_ (.A1(_03349_),
    .A2(_18054_),
    .A3(_01773_),
    .B1(_01778_),
    .X(_03350_));
 sky130_fd_sc_hd__and2_1 _31602_ (.A(_25308_),
    .B(_01770_),
    .X(_03351_));
 sky130_fd_sc_hd__o21ai_2 _31603_ (.A1(_01757_),
    .A2(_01771_),
    .B1(_01760_),
    .Y(_03352_));
 sky130_fd_sc_hd__nor2_1 _31604_ (.A(_25311_),
    .B(_01770_),
    .Y(_03353_));
 sky130_fd_sc_hd__inv_2 _31605_ (.A(_01760_),
    .Y(_03354_));
 sky130_fd_sc_hd__o21ai_2 _31606_ (.A1(_03351_),
    .A2(_03353_),
    .B1(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__a21bo_1 _31607_ (.A1(_01760_),
    .A2(_01757_),
    .B1_N(_01758_),
    .X(_03356_));
 sky130_fd_sc_hd__o211ai_4 _31608_ (.A1(_03351_),
    .A2(_03352_),
    .B1(_03355_),
    .C1(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__inv_2 _31609_ (.A(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31610_ (.A(_25311_),
    .X(_03360_));
 sky130_fd_sc_hd__a21o_1 _31611_ (.A1(_03360_),
    .A2(_01771_),
    .B1(_03352_),
    .X(_03361_));
 sky130_fd_sc_hd__a21oi_1 _31612_ (.A1(_03361_),
    .A2(_03355_),
    .B1(_03356_),
    .Y(_03362_));
 sky130_fd_sc_hd__o21bai_1 _31613_ (.A1(_03358_),
    .A2(_03362_),
    .B1_N(_23954_),
    .Y(_03363_));
 sky130_fd_sc_hd__nand3b_1 _31614_ (.A_N(_03362_),
    .B(_23954_),
    .C(_03357_),
    .Y(_03364_));
 sky130_fd_sc_hd__or2b_1 _31615_ (.A(_18052_),
    .B_N(_03347_),
    .X(_03365_));
 sky130_fd_sc_hd__nand2_1 _31616_ (.A(_25310_),
    .B(_01772_),
    .Y(_03366_));
 sky130_fd_sc_hd__clkbuf_2 _31617_ (.A(\delay_line[8][13] ),
    .X(_03367_));
 sky130_fd_sc_hd__buf_1 _31618_ (.A(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_2 _31619_ (.A(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__xnor2_2 _31620_ (.A(_17916_),
    .B(_03369_),
    .Y(_03371_));
 sky130_fd_sc_hd__and3_1 _31621_ (.A(_03365_),
    .B(_03366_),
    .C(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__a21oi_1 _31622_ (.A1(_03365_),
    .A2(_03366_),
    .B1(_03371_),
    .Y(_03373_));
 sky130_fd_sc_hd__a211oi_1 _31623_ (.A1(_03363_),
    .A2(_03364_),
    .B1(_03372_),
    .C1(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__o211a_1 _31624_ (.A1(_03372_),
    .A2(_03373_),
    .B1(_03363_),
    .C1(_03364_),
    .X(_03375_));
 sky130_fd_sc_hd__nor2_2 _31625_ (.A(_03374_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__xnor2_1 _31626_ (.A(_03350_),
    .B(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__nor3_2 _31627_ (.A(_03345_),
    .B(_03346_),
    .C(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__o21a_1 _31628_ (.A1(_03345_),
    .A2(_03346_),
    .B1(_03377_),
    .X(_03379_));
 sky130_fd_sc_hd__nor2_1 _31629_ (.A(_03378_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand3_1 _31630_ (.A(_03332_),
    .B(_03333_),
    .C(_03380_),
    .Y(_03382_));
 sky130_fd_sc_hd__a21o_1 _31631_ (.A1(_03332_),
    .A2(_03333_),
    .B1(_03380_),
    .X(_03383_));
 sky130_fd_sc_hd__and3_1 _31632_ (.A(_03309_),
    .B(_03382_),
    .C(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_2 _31633_ (.A(_03382_),
    .X(_03385_));
 sky130_fd_sc_hd__a21oi_2 _31634_ (.A1(_03385_),
    .A2(_03383_),
    .B1(_03309_),
    .Y(_03386_));
 sky130_fd_sc_hd__nor3_2 _31635_ (.A(_03308_),
    .B(_03384_),
    .C(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__a21boi_1 _31636_ (.A1(_03385_),
    .A2(_03383_),
    .B1_N(_03309_),
    .Y(_03388_));
 sky130_fd_sc_hd__nand4bb_1 _31637_ (.A_N(_01720_),
    .B_N(_01731_),
    .C(_03382_),
    .D(_03383_),
    .Y(_03389_));
 sky130_fd_sc_hd__and3b_1 _31638_ (.A_N(_03388_),
    .B(_03308_),
    .C(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__nor2_1 _31639_ (.A(_03387_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__nand2_2 _31640_ (.A(_03307_),
    .B(_03391_),
    .Y(_03393_));
 sky130_fd_sc_hd__nor2_1 _31641_ (.A(_03302_),
    .B(_03303_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand2_1 _31642_ (.A(_03257_),
    .B(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__o211a_2 _31643_ (.A1(_03237_),
    .A2(_03242_),
    .B1(_03244_),
    .C1(_03251_),
    .X(_03396_));
 sky130_fd_sc_hd__a21o_1 _31644_ (.A1(_01734_),
    .A2(_01824_),
    .B1(_01826_),
    .X(_03397_));
 sky130_fd_sc_hd__o2bb2ai_2 _31645_ (.A1_N(_03252_),
    .A2_N(_03257_),
    .B1(_03302_),
    .B2(_03303_),
    .Y(_03398_));
 sky130_fd_sc_hd__o211a_4 _31646_ (.A1(_03395_),
    .A2(_03396_),
    .B1(_03397_),
    .C1(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__a21o_2 _31647_ (.A1(_01737_),
    .A2(_01822_),
    .B1(_01829_),
    .X(_03400_));
 sky130_fd_sc_hd__o211ai_4 _31648_ (.A1(_03395_),
    .A2(_03396_),
    .B1(_03397_),
    .C1(_03398_),
    .Y(_03401_));
 sky130_fd_sc_hd__o2bb2ai_2 _31649_ (.A1_N(_03401_),
    .A2_N(_03307_),
    .B1(_03387_),
    .B2(_03390_),
    .Y(_03402_));
 sky130_fd_sc_hd__o211ai_4 _31650_ (.A1(_03393_),
    .A2(_03399_),
    .B1(_03400_),
    .C1(_03402_),
    .Y(_03404_));
 sky130_fd_sc_hd__a21bo_1 _31651_ (.A1(_03401_),
    .A2(_03307_),
    .B1_N(_03391_),
    .X(_03405_));
 sky130_fd_sc_hd__o211ai_4 _31652_ (.A1(_03387_),
    .A2(_03390_),
    .B1(_03401_),
    .C1(_03307_),
    .Y(_03406_));
 sky130_fd_sc_hd__a21oi_4 _31653_ (.A1(_01737_),
    .A2(_01822_),
    .B1(_01829_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand3_2 _31654_ (.A(_03405_),
    .B(_03406_),
    .C(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__o21a_1 _31655_ (.A1(_25327_),
    .A2(_25330_),
    .B1(_01935_),
    .X(_03409_));
 sky130_fd_sc_hd__nor2_1 _31656_ (.A(_01932_),
    .B(_01933_),
    .Y(_03410_));
 sky130_fd_sc_hd__a21oi_1 _31657_ (.A1(_01910_),
    .A2(_00272_),
    .B1(_01934_),
    .Y(_03411_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31658_ (.A(_21862_),
    .X(_03412_));
 sky130_fd_sc_hd__buf_1 _31659_ (.A(net425),
    .X(_03413_));
 sky130_fd_sc_hd__nor2_1 _31660_ (.A(_03412_),
    .B(_03413_),
    .Y(_03415_));
 sky130_fd_sc_hd__and2_1 _31661_ (.A(_21862_),
    .B(_22525_),
    .X(_03416_));
 sky130_fd_sc_hd__or3b_2 _31662_ (.A(_03415_),
    .B(_03416_),
    .C_N(_01912_),
    .X(_03417_));
 sky130_fd_sc_hd__o21bai_2 _31663_ (.A1(_03415_),
    .A2(_03416_),
    .B1_N(_01912_),
    .Y(_03418_));
 sky130_fd_sc_hd__o21ai_1 _31664_ (.A1(_00265_),
    .A2(_22527_),
    .B1(_00253_),
    .Y(_03419_));
 sky130_fd_sc_hd__and2b_1 _31665_ (.A_N(_00252_),
    .B(net426),
    .X(_03420_));
 sky130_fd_sc_hd__and2b_1 _31666_ (.A_N(net426),
    .B(_00252_),
    .X(_03421_));
 sky130_fd_sc_hd__a211o_2 _31667_ (.A1(_01914_),
    .A2(_03419_),
    .B1(_03420_),
    .C1(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__o211ai_2 _31668_ (.A1(_03420_),
    .A2(_03421_),
    .B1(_01914_),
    .C1(_03419_),
    .Y(_03423_));
 sky130_fd_sc_hd__clkbuf_2 _31669_ (.A(_01920_),
    .X(_03424_));
 sky130_fd_sc_hd__nand4_4 _31670_ (.A(_21910_),
    .B(_03422_),
    .C(_03423_),
    .D(_03424_),
    .Y(_03426_));
 sky130_fd_sc_hd__a22o_1 _31671_ (.A1(_21910_),
    .A2(_03424_),
    .B1(_03422_),
    .B2(_03423_),
    .X(_03427_));
 sky130_fd_sc_hd__nand4_4 _31672_ (.A(_03417_),
    .B(_03418_),
    .C(_03426_),
    .D(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__a22o_1 _31673_ (.A1(_03417_),
    .A2(_03418_),
    .B1(_03426_),
    .B2(_03427_),
    .X(_03429_));
 sky130_fd_sc_hd__a211o_1 _31674_ (.A1(_03428_),
    .A2(_03429_),
    .B1(_01751_),
    .C1(net180),
    .X(_03430_));
 sky130_fd_sc_hd__o211ai_1 _31675_ (.A1(_01751_),
    .A2(net180),
    .B1(_03428_),
    .C1(_03429_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _31676_ (.A(_03430_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__xor2_1 _31677_ (.A(_01929_),
    .B(_03432_),
    .X(_03433_));
 sky130_fd_sc_hd__a21bo_1 _31678_ (.A1(_01782_),
    .A2(_01756_),
    .B1_N(_01781_),
    .X(_03434_));
 sky130_fd_sc_hd__xor2_1 _31679_ (.A(_03433_),
    .B(_03434_),
    .X(_03435_));
 sky130_fd_sc_hd__o21a_1 _31680_ (.A1(_03410_),
    .A2(_03411_),
    .B1(_03435_),
    .X(_03437_));
 sky130_fd_sc_hd__nor3_1 _31681_ (.A(_03410_),
    .B(_03411_),
    .C(_03435_),
    .Y(_03438_));
 sky130_fd_sc_hd__nor2_1 _31682_ (.A(_03437_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nor3_2 _31683_ (.A(_03409_),
    .B(_01938_),
    .C(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21a_1 _31684_ (.A1(_03409_),
    .A2(_01938_),
    .B1(_03439_),
    .X(_03441_));
 sky130_fd_sc_hd__nand2_1 _31685_ (.A(_01896_),
    .B(_01899_),
    .Y(_03442_));
 sky130_fd_sc_hd__or2b_1 _31686_ (.A(_21978_),
    .B_N(\delay_line[5][13] ),
    .X(_03443_));
 sky130_fd_sc_hd__or2b_1 _31687_ (.A(\delay_line[5][13] ),
    .B_N(_24058_),
    .X(_03444_));
 sky130_fd_sc_hd__and3_1 _31688_ (.A(_03443_),
    .B(_03444_),
    .C(_01869_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_2 _31689_ (.A(_03443_),
    .X(_03446_));
 sky130_fd_sc_hd__a21oi_2 _31690_ (.A1(_03446_),
    .A2(_03444_),
    .B1(_01869_),
    .Y(_03448_));
 sky130_fd_sc_hd__a211oi_4 _31691_ (.A1(_01871_),
    .A2(_01873_),
    .B1(_03445_),
    .C1(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__o211a_1 _31692_ (.A1(_03445_),
    .A2(_03448_),
    .B1(_01871_),
    .C1(_01873_),
    .X(_03450_));
 sky130_fd_sc_hd__a2111oi_4 _31693_ (.A1(_00196_),
    .A2(_00201_),
    .B1(_01876_),
    .C1(_03449_),
    .D1(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__o21a_1 _31694_ (.A1(_03449_),
    .A2(_03450_),
    .B1(_01878_),
    .X(_03452_));
 sky130_fd_sc_hd__nor2_1 _31695_ (.A(_03451_),
    .B(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31696_ (.A(\delay_line[3][13] ),
    .X(_03454_));
 sky130_fd_sc_hd__and2_1 _31697_ (.A(_22642_),
    .B(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__nor2_1 _31698_ (.A(_03454_),
    .B(_22643_),
    .Y(_03456_));
 sky130_fd_sc_hd__clkbuf_2 _31699_ (.A(_01872_),
    .X(_03457_));
 sky130_fd_sc_hd__or3b_1 _31700_ (.A(_03455_),
    .B(_03456_),
    .C_N(_03457_),
    .X(_03459_));
 sky130_fd_sc_hd__o21bai_1 _31701_ (.A1(_03455_),
    .A2(_03456_),
    .B1_N(_03457_),
    .Y(_03460_));
 sky130_fd_sc_hd__and3_1 _31702_ (.A(_03453_),
    .B(_03459_),
    .C(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__o2bb2a_1 _31703_ (.A1_N(_03460_),
    .A2_N(_03459_),
    .B1(_03451_),
    .B2(_03452_),
    .X(_03462_));
 sky130_fd_sc_hd__nor2_1 _31704_ (.A(_03461_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__clkbuf_2 _31705_ (.A(_01888_),
    .X(_03464_));
 sky130_fd_sc_hd__o21ai_2 _31706_ (.A1(_01885_),
    .A2(_03464_),
    .B1(_00211_),
    .Y(_03465_));
 sky130_fd_sc_hd__o21ai_1 _31707_ (.A1(_01885_),
    .A2(_01888_),
    .B1(_01924_),
    .Y(_03466_));
 sky130_fd_sc_hd__or3_1 _31708_ (.A(_01884_),
    .B(_24062_),
    .C(net427),
    .X(_03467_));
 sky130_fd_sc_hd__nand2_1 _31709_ (.A(_03466_),
    .B(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand3_1 _31710_ (.A(_01923_),
    .B(_01926_),
    .C(_03468_),
    .Y(_03470_));
 sky130_fd_sc_hd__a21o_1 _31711_ (.A1(_01923_),
    .A2(_01926_),
    .B1(_03468_),
    .X(_03471_));
 sky130_fd_sc_hd__nand2_1 _31712_ (.A(_03470_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__xor2_1 _31713_ (.A(_03465_),
    .B(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__and2b_1 _31714_ (.A_N(_01893_),
    .B(_01894_),
    .X(_03474_));
 sky130_fd_sc_hd__and2b_1 _31715_ (.A_N(_03473_),
    .B(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__and2b_1 _31716_ (.A_N(_03474_),
    .B(_03473_),
    .X(_03476_));
 sky130_fd_sc_hd__nor2_1 _31717_ (.A(_03475_),
    .B(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__xnor2_2 _31718_ (.A(_03463_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__xnor2_2 _31719_ (.A(_03442_),
    .B(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__o21bai_2 _31720_ (.A1(_00234_),
    .A2(_01851_),
    .B1_N(_01850_),
    .Y(_03481_));
 sky130_fd_sc_hd__and2b_1 _31721_ (.A_N(\delay_line[3][11] ),
    .B(net439),
    .X(_03482_));
 sky130_fd_sc_hd__or2b_1 _31722_ (.A(net439),
    .B_N(_00207_),
    .X(_03483_));
 sky130_fd_sc_hd__or3b_1 _31723_ (.A(_01860_),
    .B(_03482_),
    .C_N(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__or2b_1 _31724_ (.A(_00207_),
    .B_N(net439),
    .X(_03485_));
 sky130_fd_sc_hd__a21bo_1 _31725_ (.A1(_03485_),
    .A2(_03483_),
    .B1_N(_01860_),
    .X(_03486_));
 sky130_fd_sc_hd__a21boi_1 _31726_ (.A1(_03484_),
    .A2(_03486_),
    .B1_N(_01843_),
    .Y(_03487_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31727_ (.A(\delay_line[2][12] ),
    .X(_03488_));
 sky130_fd_sc_hd__and4b_2 _31728_ (.A_N(_24016_),
    .B(_03484_),
    .C(_03486_),
    .D(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__nor3_2 _31729_ (.A(_03487_),
    .B(_01867_),
    .C(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__o21a_1 _31730_ (.A1(_03489_),
    .A2(_03487_),
    .B1(_01867_),
    .X(_03492_));
 sky130_fd_sc_hd__a211oi_2 _31731_ (.A1(_01846_),
    .A2(_01849_),
    .B1(_03490_),
    .C1(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__o211a_1 _31732_ (.A1(_03490_),
    .A2(_03492_),
    .B1(_01846_),
    .C1(_01849_),
    .X(_03494_));
 sky130_fd_sc_hd__a211oi_1 _31733_ (.A1(_01880_),
    .A2(_01881_),
    .B1(_03493_),
    .C1(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__o211a_1 _31734_ (.A1(_03493_),
    .A2(_03494_),
    .B1(_01880_),
    .C1(_01881_),
    .X(_03496_));
 sky130_fd_sc_hd__nor2_1 _31735_ (.A(_03495_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__xor2_2 _31736_ (.A(_03481_),
    .B(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__xnor2_1 _31737_ (.A(_03479_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__o21ai_2 _31738_ (.A1(_03440_),
    .A2(_03441_),
    .B1(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__or3_1 _31739_ (.A(_03440_),
    .B(_03441_),
    .C(_03499_),
    .X(_03501_));
 sky130_fd_sc_hd__o21a_2 _31740_ (.A1(_01738_),
    .A2(_01815_),
    .B1(_01816_),
    .X(_03503_));
 sky130_fd_sc_hd__a21boi_2 _31741_ (.A1(_03500_),
    .A2(_03501_),
    .B1_N(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__nand3b_2 _31742_ (.A_N(_03503_),
    .B(_03500_),
    .C(_03501_),
    .Y(_03505_));
 sky130_fd_sc_hd__inv_2 _31743_ (.A(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__or2b_2 _31744_ (.A(_01905_),
    .B_N(_01942_),
    .X(_03507_));
 sky130_fd_sc_hd__o211a_2 _31745_ (.A1(_03504_),
    .A2(_03506_),
    .B1(_01940_),
    .C1(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__a211oi_4 _31746_ (.A1(_01940_),
    .A2(_03507_),
    .B1(_03504_),
    .C1(_03506_),
    .Y(_03509_));
 sky130_fd_sc_hd__o2bb2ai_4 _31747_ (.A1_N(_03404_),
    .A2_N(_03408_),
    .B1(_03508_),
    .B2(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__nor2_1 _31748_ (.A(_03508_),
    .B(_03509_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand3_1 _31749_ (.A(_03404_),
    .B(_03408_),
    .C(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__a21o_2 _31750_ (.A1(_01838_),
    .A2(_01954_),
    .B1(_01970_),
    .X(_03514_));
 sky130_fd_sc_hd__a21o_1 _31751_ (.A1(_03510_),
    .A2(_03512_),
    .B1(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__o211a_4 _31752_ (.A1(_03393_),
    .A2(_03399_),
    .B1(_03400_),
    .C1(_03402_),
    .X(_03516_));
 sky130_fd_sc_hd__nand2_1 _31753_ (.A(_03408_),
    .B(_03511_),
    .Y(_03517_));
 sky130_fd_sc_hd__o211ai_4 _31754_ (.A1(_03516_),
    .A2(_03517_),
    .B1(_03510_),
    .C1(_03514_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand3_2 _31755_ (.A(_03122_),
    .B(_03515_),
    .C(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__a21oi_2 _31756_ (.A1(_03510_),
    .A2(_03512_),
    .B1(_03514_),
    .Y(_03520_));
 sky130_fd_sc_hd__o211a_1 _31757_ (.A1(_03517_),
    .A2(_03516_),
    .B1(_03514_),
    .C1(_03510_),
    .X(_03521_));
 sky130_fd_sc_hd__xor2_2 _31758_ (.A(_03075_),
    .B(_03121_),
    .X(_03522_));
 sky130_fd_sc_hd__o21ai_2 _31759_ (.A1(_03520_),
    .A2(_03521_),
    .B1(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__o211ai_4 _31760_ (.A1(_01972_),
    .A2(_03074_),
    .B1(_03519_),
    .C1(_03523_),
    .Y(_03525_));
 sky130_fd_sc_hd__o21a_1 _31761_ (.A1(_01522_),
    .A2(_01967_),
    .B1(_01958_),
    .X(_03526_));
 sky130_fd_sc_hd__nor3_1 _31762_ (.A(_03522_),
    .B(_03520_),
    .C(_03521_),
    .Y(_03527_));
 sky130_fd_sc_hd__a21oi_1 _31763_ (.A1(_03515_),
    .A2(_03518_),
    .B1(_03122_),
    .Y(_03528_));
 sky130_fd_sc_hd__o22ai_4 _31764_ (.A1(_01969_),
    .A2(_03526_),
    .B1(net69),
    .B2(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__o21ai_2 _31765_ (.A1(_00354_),
    .A2(_01966_),
    .B1(_01521_),
    .Y(_03530_));
 sky130_fd_sc_hd__clkbuf_2 _31766_ (.A(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__a21oi_1 _31767_ (.A1(_03525_),
    .A2(_03529_),
    .B1(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__a211oi_2 _31768_ (.A1(_01960_),
    .A2(_01962_),
    .B1(_01987_),
    .C1(_01976_),
    .Y(_03533_));
 sky130_fd_sc_hd__o211ai_2 _31769_ (.A1(_01519_),
    .A2(_01967_),
    .B1(_03525_),
    .C1(_03529_),
    .Y(_03534_));
 sky130_fd_sc_hd__o21ai_1 _31770_ (.A1(_01978_),
    .A2(_03533_),
    .B1(_03534_),
    .Y(_03536_));
 sky130_fd_sc_hd__o21ai_1 _31771_ (.A1(_01524_),
    .A2(_01969_),
    .B1(_01958_),
    .Y(_03537_));
 sky130_fd_sc_hd__a21oi_1 _31772_ (.A1(_03519_),
    .A2(_03523_),
    .B1(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__clkbuf_2 _31773_ (.A(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__a31o_1 _31774_ (.A1(_03523_),
    .A2(_03537_),
    .A3(_03519_),
    .B1(_03531_),
    .X(_03540_));
 sky130_fd_sc_hd__o22a_2 _31775_ (.A1(_01983_),
    .A2(_01982_),
    .B1(_01987_),
    .B2(_01976_),
    .X(_03541_));
 sky130_fd_sc_hd__o211a_2 _31776_ (.A1(_01972_),
    .A2(_03074_),
    .B1(_03519_),
    .C1(_03523_),
    .X(_03542_));
 sky130_fd_sc_hd__o21ai_2 _31777_ (.A1(_03542_),
    .A2(_03539_),
    .B1(_03531_),
    .Y(_03543_));
 sky130_fd_sc_hd__o211ai_4 _31778_ (.A1(_03539_),
    .A2(_03540_),
    .B1(_03541_),
    .C1(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__o21a_1 _31779_ (.A1(_03532_),
    .A2(_03536_),
    .B1(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__nand2_1 _31780_ (.A(_03072_),
    .B(_03545_),
    .Y(_03547_));
 sky130_fd_sc_hd__inv_2 _31781_ (.A(_03530_),
    .Y(_03548_));
 sky130_fd_sc_hd__o21ai_1 _31782_ (.A1(_03542_),
    .A2(_03538_),
    .B1(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__o211a_1 _31783_ (.A1(_01978_),
    .A2(_03533_),
    .B1(_03534_),
    .C1(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__o211a_1 _31784_ (.A1(_03539_),
    .A2(_03540_),
    .B1(_03541_),
    .C1(_03543_),
    .X(_03551_));
 sky130_fd_sc_hd__buf_2 _31785_ (.A(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__o221ai_4 _31786_ (.A1(_03070_),
    .A2(_03069_),
    .B1(_03550_),
    .B2(_03552_),
    .C1(_02000_),
    .Y(_03553_));
 sky130_fd_sc_hd__o211ai_2 _31787_ (.A1(_03067_),
    .A2(_03068_),
    .B1(_03547_),
    .C1(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__o21a_2 _31788_ (.A1(_02728_),
    .A2(_02715_),
    .B1(_02713_),
    .X(_03555_));
 sky130_fd_sc_hd__a31oi_1 _31789_ (.A1(_03530_),
    .A2(_03525_),
    .A3(_03529_),
    .B1(_03541_),
    .Y(_03556_));
 sky130_fd_sc_hd__a2bb2oi_2 _31790_ (.A1_N(_03069_),
    .A2_N(_03070_),
    .B1(_03549_),
    .B2(_03556_),
    .Y(_03558_));
 sky130_fd_sc_hd__o21ai_4 _31791_ (.A1(_01990_),
    .A2(_03071_),
    .B1(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__nor2_2 _31792_ (.A(_03067_),
    .B(_03068_),
    .Y(_03560_));
 sky130_fd_sc_hd__o2bb2ai_2 _31793_ (.A1_N(_01989_),
    .A2_N(_02000_),
    .B1(_03551_),
    .B2(_03550_),
    .Y(_03561_));
 sky130_fd_sc_hd__o211ai_2 _31794_ (.A1(_03552_),
    .A2(_03559_),
    .B1(_03560_),
    .C1(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__nand3_4 _31795_ (.A(_03554_),
    .B(_03555_),
    .C(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__buf_2 _31796_ (.A(\delay_line[23][12] ),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_2 _31797_ (.A(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__nand2_2 _31798_ (.A(_02016_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__a21oi_2 _31799_ (.A1(_03566_),
    .A2(_02001_),
    .B1(_02003_),
    .Y(_03567_));
 sky130_fd_sc_hd__nand2_1 _31800_ (.A(_03563_),
    .B(_03567_),
    .Y(_03569_));
 sky130_fd_sc_hd__o21ai_2 _31801_ (.A1(_02728_),
    .A2(_02715_),
    .B1(_02713_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand3_1 _31802_ (.A(_03547_),
    .B(_03553_),
    .C(_03560_),
    .Y(_03571_));
 sky130_fd_sc_hd__o221ai_4 _31803_ (.A1(_03067_),
    .A2(_03068_),
    .B1(_03552_),
    .B2(_03559_),
    .C1(_03561_),
    .Y(_03572_));
 sky130_fd_sc_hd__and3_2 _31804_ (.A(_03570_),
    .B(_03571_),
    .C(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__a21o_1 _31805_ (.A1(_02731_),
    .A2(_02785_),
    .B1(_02784_),
    .X(_03574_));
 sky130_fd_sc_hd__nand3_2 _31806_ (.A(_03570_),
    .B(_03571_),
    .C(_03572_),
    .Y(_03575_));
 sky130_fd_sc_hd__a21o_1 _31807_ (.A1(_03575_),
    .A2(_03563_),
    .B1(_03567_),
    .X(_03576_));
 sky130_fd_sc_hd__o211ai_2 _31808_ (.A1(_03569_),
    .A2(_03573_),
    .B1(_03574_),
    .C1(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__a21bo_1 _31809_ (.A1(_03575_),
    .A2(_03563_),
    .B1_N(_03567_),
    .X(_03578_));
 sky130_fd_sc_hd__nand3b_1 _31810_ (.A_N(_03567_),
    .B(_03575_),
    .C(_03563_),
    .Y(_03580_));
 sky130_fd_sc_hd__inv_2 _31811_ (.A(_03574_),
    .Y(_03581_));
 sky130_fd_sc_hd__nand3_2 _31812_ (.A(_03578_),
    .B(_03580_),
    .C(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__a21oi_2 _31813_ (.A1(_02021_),
    .A2(_02014_),
    .B1(_02011_),
    .Y(_03583_));
 sky130_fd_sc_hd__a21oi_1 _31814_ (.A1(_03577_),
    .A2(_03582_),
    .B1(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__and3_1 _31815_ (.A(_03577_),
    .B(_03582_),
    .C(_03583_),
    .X(_03585_));
 sky130_fd_sc_hd__a21bo_1 _31816_ (.A1(_02033_),
    .A2(_02027_),
    .B1_N(_02032_),
    .X(_03586_));
 sky130_fd_sc_hd__o21bai_2 _31817_ (.A1(_03584_),
    .A2(_03585_),
    .B1_N(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__buf_1 _31818_ (.A(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__and2_1 _31819_ (.A(_22761_),
    .B(\delay_line[23][11] ),
    .X(_03589_));
 sky130_fd_sc_hd__nor2_1 _31820_ (.A(_22761_),
    .B(_02002_),
    .Y(_03591_));
 sky130_fd_sc_hd__or3b_1 _31821_ (.A(_03589_),
    .B(_03591_),
    .C_N(_02042_),
    .X(_03592_));
 sky130_fd_sc_hd__a2bb2o_1 _31822_ (.A1_N(_03589_),
    .A2_N(_03591_),
    .B1(_24286_),
    .B2(_02019_),
    .X(_03593_));
 sky130_fd_sc_hd__nand2_1 _31823_ (.A(_03592_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__or3b_1 _31824_ (.A(_15394_),
    .B(_19848_),
    .C_N(_17897_),
    .X(_03595_));
 sky130_fd_sc_hd__o21ai_2 _31825_ (.A1(_10361_),
    .A2(_15053_),
    .B1(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__xor2_2 _31826_ (.A(_03594_),
    .B(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__nand2_1 _31827_ (.A(_03588_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__nand2_2 _31828_ (.A(_03582_),
    .B(_03583_),
    .Y(_03599_));
 sky130_fd_sc_hd__o211a_2 _31829_ (.A1(_03569_),
    .A2(_03573_),
    .B1(_03574_),
    .C1(_03576_),
    .X(_03600_));
 sky130_fd_sc_hd__a22o_1 _31830_ (.A1(_02024_),
    .A2(_02022_),
    .B1(_03577_),
    .B2(_03582_),
    .X(_03602_));
 sky130_fd_sc_hd__o211a_2 _31831_ (.A1(_03599_),
    .A2(_03600_),
    .B1(_03586_),
    .C1(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__o21ai_4 _31832_ (.A1(_02681_),
    .A2(_02919_),
    .B1(_02923_),
    .Y(_03604_));
 sky130_fd_sc_hd__o211ai_4 _31833_ (.A1(_03599_),
    .A2(_03600_),
    .B1(_03586_),
    .C1(_03602_),
    .Y(_03605_));
 sky130_fd_sc_hd__a21o_1 _31834_ (.A1(_03587_),
    .A2(_03605_),
    .B1(_03597_),
    .X(_03606_));
 sky130_fd_sc_hd__o211ai_2 _31835_ (.A1(_03598_),
    .A2(_03603_),
    .B1(_03604_),
    .C1(_03606_),
    .Y(_03607_));
 sky130_fd_sc_hd__buf_1 _31836_ (.A(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__inv_2 _31837_ (.A(_03597_),
    .Y(_03609_));
 sky130_fd_sc_hd__a21o_1 _31838_ (.A1(_03588_),
    .A2(_03605_),
    .B1(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__inv_2 _31839_ (.A(_03604_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand3_1 _31840_ (.A(_03588_),
    .B(_03605_),
    .C(_03609_),
    .Y(_03613_));
 sky130_fd_sc_hd__nand3_2 _31841_ (.A(_03610_),
    .B(_03611_),
    .C(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__o21a_1 _31842_ (.A1(_02047_),
    .A2(_02048_),
    .B1(_02049_),
    .X(_03615_));
 sky130_fd_sc_hd__a31o_1 _31843_ (.A1(_02054_),
    .A2(_02052_),
    .A3(_02053_),
    .B1(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__a21oi_1 _31844_ (.A1(_03608_),
    .A2(_03614_),
    .B1(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__o211a_1 _31845_ (.A1(_02037_),
    .A2(_03615_),
    .B1(_03607_),
    .C1(_03614_),
    .X(_03618_));
 sky130_fd_sc_hd__a2bb2o_1 _31846_ (.A1_N(_02679_),
    .A2_N(_02924_),
    .B1(_02071_),
    .B2(_02677_),
    .X(_03619_));
 sky130_fd_sc_hd__o21ai_2 _31847_ (.A1(_02786_),
    .A2(_02918_),
    .B1(_02917_),
    .Y(_03620_));
 sky130_fd_sc_hd__o21ba_1 _31848_ (.A1(_01240_),
    .A2(_01241_),
    .B1_N(_02705_),
    .X(_03621_));
 sky130_fd_sc_hd__buf_1 _31849_ (.A(_01233_),
    .X(_03622_));
 sky130_fd_sc_hd__buf_1 _31850_ (.A(\delay_line[39][12] ),
    .X(_03624_));
 sky130_fd_sc_hd__nand2_1 _31851_ (.A(_03622_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__nor2_1 _31852_ (.A(_03624_),
    .B(\delay_line[39][13] ),
    .Y(_03626_));
 sky130_fd_sc_hd__nand2_1 _31853_ (.A(\delay_line[39][12] ),
    .B(\delay_line[39][13] ),
    .Y(_03627_));
 sky130_fd_sc_hd__and2b_1 _31854_ (.A_N(_03626_),
    .B(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__xnor2_1 _31855_ (.A(_03622_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__a21oi_1 _31856_ (.A1(_03625_),
    .A2(_02697_),
    .B1(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__nand3_1 _31857_ (.A(_03625_),
    .B(_02697_),
    .C(_03629_),
    .Y(_03631_));
 sky130_fd_sc_hd__and2b_1 _31858_ (.A_N(_03630_),
    .B(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__xnor2_1 _31859_ (.A(_02693_),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__nor3b_1 _31860_ (.A(_02701_),
    .B(_02702_),
    .C_N(_03633_),
    .Y(_03635_));
 sky130_fd_sc_hd__o21ba_1 _31861_ (.A1(_02701_),
    .A2(_02702_),
    .B1_N(_03633_),
    .X(_03636_));
 sky130_fd_sc_hd__nor2_1 _31862_ (.A(_03635_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__nor3_1 _31863_ (.A(_03621_),
    .B(_02708_),
    .C(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__o21a_1 _31864_ (.A1(_03621_),
    .A2(_02708_),
    .B1(_03637_),
    .X(_03639_));
 sky130_fd_sc_hd__nor2_1 _31865_ (.A(_03638_),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__nor2_1 _31866_ (.A(_02682_),
    .B(_02684_),
    .Y(_03641_));
 sky130_fd_sc_hd__buf_1 _31867_ (.A(\delay_line[38][11] ),
    .X(_03642_));
 sky130_fd_sc_hd__nor2_1 _31868_ (.A(_02686_),
    .B(\delay_line[38][13] ),
    .Y(_03643_));
 sky130_fd_sc_hd__and2_1 _31869_ (.A(_02686_),
    .B(\delay_line[38][13] ),
    .X(_03644_));
 sky130_fd_sc_hd__nor2_1 _31870_ (.A(_03643_),
    .B(_03644_),
    .Y(_03646_));
 sky130_fd_sc_hd__a311o_1 _31871_ (.A1(_01215_),
    .A2(_03642_),
    .A3(_03641_),
    .B1(_03646_),
    .C1(_02684_),
    .X(_03647_));
 sky130_fd_sc_hd__a31o_1 _31872_ (.A1(_01215_),
    .A2(_03642_),
    .A3(_03641_),
    .B1(_02684_),
    .X(_03648_));
 sky130_fd_sc_hd__or3b_1 _31873_ (.A(_03643_),
    .B(_03644_),
    .C_N(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__a221o_1 _31874_ (.A1(_03641_),
    .A2(_02687_),
    .B1(_03647_),
    .B2(_03649_),
    .C1(_02692_),
    .X(_03650_));
 sky130_fd_sc_hd__a31o_1 _31875_ (.A1(_25032_),
    .A2(_01224_),
    .A3(_03641_),
    .B1(_02692_),
    .X(_03651_));
 sky130_fd_sc_hd__and3_1 _31876_ (.A(_03647_),
    .B(_03649_),
    .C(_03651_),
    .X(_03652_));
 sky130_fd_sc_hd__inv_2 _31877_ (.A(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__and3_1 _31878_ (.A(_03640_),
    .B(_03650_),
    .C(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__a21o_1 _31879_ (.A1(_03653_),
    .A2(_03650_),
    .B1(_03640_),
    .X(_03655_));
 sky130_fd_sc_hd__and2b_1 _31880_ (.A_N(_03654_),
    .B(_03655_),
    .X(_03657_));
 sky130_fd_sc_hd__buf_1 _31881_ (.A(_01254_),
    .X(_03658_));
 sky130_fd_sc_hd__clkbuf_2 _31882_ (.A(\delay_line[40][11] ),
    .X(_03659_));
 sky130_fd_sc_hd__nand2_1 _31883_ (.A(_03658_),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__buf_1 _31884_ (.A(\delay_line[40][12] ),
    .X(_03661_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31885_ (.A(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_2 _31886_ (.A(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__nor2_1 _31887_ (.A(_03661_),
    .B(\delay_line[40][13] ),
    .Y(_03664_));
 sky130_fd_sc_hd__and2_1 _31888_ (.A(_03661_),
    .B(\delay_line[40][13] ),
    .X(_03665_));
 sky130_fd_sc_hd__a2bb2o_1 _31889_ (.A1_N(_03664_),
    .A2_N(_03665_),
    .B1(_03659_),
    .B2(_03661_),
    .X(_03666_));
 sky130_fd_sc_hd__or3b_1 _31890_ (.A(_02719_),
    .B(\delay_line[40][13] ),
    .C_N(_03661_),
    .X(_03668_));
 sky130_fd_sc_hd__a21oi_1 _31891_ (.A1(_03666_),
    .A2(_03668_),
    .B1(_23465_),
    .Y(_03669_));
 sky130_fd_sc_hd__and3_1 _31892_ (.A(_03666_),
    .B(_03668_),
    .C(_23465_),
    .X(_03670_));
 sky130_fd_sc_hd__nand2_1 _31893_ (.A(_23464_),
    .B(_02721_),
    .Y(_03671_));
 sky130_fd_sc_hd__o221a_1 _31894_ (.A1(_03660_),
    .A2(_03663_),
    .B1(_03669_),
    .B2(_03670_),
    .C1(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__or3b_1 _31895_ (.A(_03662_),
    .B(_02719_),
    .C_N(_03658_),
    .X(_03673_));
 sky130_fd_sc_hd__a211oi_1 _31896_ (.A1(_03671_),
    .A2(_03673_),
    .B1(_03670_),
    .C1(_03669_),
    .Y(_03674_));
 sky130_fd_sc_hd__a21o_1 _31897_ (.A1(_02723_),
    .A2(_02724_),
    .B1(_02726_),
    .X(_03675_));
 sky130_fd_sc_hd__or3_1 _31898_ (.A(_03672_),
    .B(_03674_),
    .C(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__o21ai_1 _31899_ (.A1(_03672_),
    .A2(_03674_),
    .B1(_03675_),
    .Y(_03677_));
 sky130_fd_sc_hd__and2_2 _31900_ (.A(_03676_),
    .B(_03677_),
    .X(_03679_));
 sky130_fd_sc_hd__xnor2_4 _31901_ (.A(_03657_),
    .B(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__xnor2_1 _31902_ (.A(_02732_),
    .B(\delay_line[37][13] ),
    .Y(_03681_));
 sky130_fd_sc_hd__inv_2 _31903_ (.A(\delay_line[37][12] ),
    .Y(_03682_));
 sky130_fd_sc_hd__and3b_1 _31904_ (.A_N(_23521_),
    .B(\delay_line[37][11] ),
    .C(_02736_),
    .X(_03683_));
 sky130_fd_sc_hd__o21ba_1 _31905_ (.A1(_01269_),
    .A2(_03682_),
    .B1_N(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__xnor2_1 _31906_ (.A(_03681_),
    .B(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__o22a_1 _31907_ (.A1(_03682_),
    .A2(_02735_),
    .B1(_02739_),
    .B2(_02740_),
    .X(_03686_));
 sky130_fd_sc_hd__xor2_1 _31908_ (.A(_03685_),
    .B(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__or2b_1 _31909_ (.A(_02764_),
    .B_N(\delay_line[36][10] ),
    .X(_03688_));
 sky130_fd_sc_hd__or2b_1 _31910_ (.A(\delay_line[36][10] ),
    .B_N(_02764_),
    .X(_03690_));
 sky130_fd_sc_hd__nor3_1 _31911_ (.A(_02768_),
    .B(_02769_),
    .C(_01278_),
    .Y(_03691_));
 sky130_fd_sc_hd__buf_1 _31912_ (.A(_02768_),
    .X(_03692_));
 sky130_fd_sc_hd__o2bb2a_1 _31913_ (.A1_N(_03688_),
    .A2_N(_03690_),
    .B1(_03691_),
    .B2(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__a21oi_1 _31914_ (.A1(_02767_),
    .A2(_02770_),
    .B1(_03692_),
    .Y(_03694_));
 sky130_fd_sc_hd__and3_1 _31915_ (.A(_03694_),
    .B(_03690_),
    .C(_03688_),
    .X(_03695_));
 sky130_fd_sc_hd__and4_1 _31916_ (.A(\delay_line[36][9] ),
    .B(_01278_),
    .C(_01279_),
    .D(_01281_),
    .X(_03696_));
 sky130_fd_sc_hd__or4_1 _31917_ (.A(_02774_),
    .B(_03693_),
    .C(_03695_),
    .D(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__o22ai_2 _31918_ (.A1(_03693_),
    .A2(_03695_),
    .B1(_03696_),
    .B2(_02774_),
    .Y(_03698_));
 sky130_fd_sc_hd__nand2_1 _31919_ (.A(_03697_),
    .B(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__o31a_1 _31920_ (.A1(_01298_),
    .A2(_02750_),
    .A3(_02751_),
    .B1(_02756_),
    .X(_03701_));
 sky130_fd_sc_hd__buf_1 _31921_ (.A(_02745_),
    .X(_03702_));
 sky130_fd_sc_hd__buf_1 _31922_ (.A(net301),
    .X(_03703_));
 sky130_fd_sc_hd__and2_1 _31923_ (.A(net301),
    .B(net300),
    .X(_03704_));
 sky130_fd_sc_hd__nor2_1 _31924_ (.A(net301),
    .B(\delay_line[35][13] ),
    .Y(_03705_));
 sky130_fd_sc_hd__or3b_1 _31925_ (.A(_03704_),
    .B(_03705_),
    .C_N(_02745_),
    .X(_03706_));
 sky130_fd_sc_hd__o21bai_1 _31926_ (.A1(_03704_),
    .A2(_03705_),
    .B1_N(_02745_),
    .Y(_03707_));
 sky130_fd_sc_hd__nor3b_1 _31927_ (.A(_02746_),
    .B(_02747_),
    .C_N(_01290_),
    .Y(_03708_));
 sky130_fd_sc_hd__a221o_1 _31928_ (.A1(_03702_),
    .A2(_03703_),
    .B1(_03706_),
    .B2(_03707_),
    .C1(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__o211ai_2 _31929_ (.A1(_02747_),
    .A2(_03708_),
    .B1(_03706_),
    .C1(_03707_),
    .Y(_03710_));
 sky130_fd_sc_hd__nand3_1 _31930_ (.A(_03709_),
    .B(_02750_),
    .C(_03710_),
    .Y(_03712_));
 sky130_fd_sc_hd__a21o_1 _31931_ (.A1(_03710_),
    .A2(_03709_),
    .B1(_02750_),
    .X(_03713_));
 sky130_fd_sc_hd__nand2_1 _31932_ (.A(_03712_),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__or2_1 _31933_ (.A(_20842_),
    .B(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__nand2_1 _31934_ (.A(_03714_),
    .B(_20842_),
    .Y(_03716_));
 sky130_fd_sc_hd__and3b_1 _31935_ (.A_N(_03701_),
    .B(_03715_),
    .C(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__a21boi_1 _31936_ (.A1(_03715_),
    .A2(_03716_),
    .B1_N(_03701_),
    .Y(_03718_));
 sky130_fd_sc_hd__or2_1 _31937_ (.A(_03717_),
    .B(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__o21ai_2 _31938_ (.A1(_02761_),
    .A2(_02762_),
    .B1(_02758_),
    .Y(_03720_));
 sky130_fd_sc_hd__xor2_1 _31939_ (.A(_03719_),
    .B(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__nand2_1 _31940_ (.A(_03699_),
    .B(_03721_),
    .Y(_03723_));
 sky130_fd_sc_hd__or2_1 _31941_ (.A(_03699_),
    .B(_03721_),
    .X(_03724_));
 sky130_fd_sc_hd__nand2_1 _31942_ (.A(_03723_),
    .B(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__nor2_1 _31943_ (.A(_03687_),
    .B(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__and2_1 _31944_ (.A(_03687_),
    .B(_03725_),
    .X(_03727_));
 sky130_fd_sc_hd__or3b_1 _31945_ (.A(_02741_),
    .B(_02778_),
    .C_N(_02779_),
    .X(_03728_));
 sky130_fd_sc_hd__o211a_1 _31946_ (.A1(_03726_),
    .A2(_03727_),
    .B1(_02779_),
    .C1(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__a211o_1 _31947_ (.A1(_02779_),
    .A2(_03728_),
    .B1(_03726_),
    .C1(_03727_),
    .X(_03730_));
 sky130_fd_sc_hd__and2b_1 _31948_ (.A_N(_03729_),
    .B(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__xnor2_4 _31949_ (.A(_03680_),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__a21oi_1 _31950_ (.A1(_02787_),
    .A2(_02910_),
    .B1(_02913_),
    .Y(_03734_));
 sky130_fd_sc_hd__buf_1 _31951_ (.A(\delay_line[34][10] ),
    .X(_03735_));
 sky130_fd_sc_hd__or2_1 _31952_ (.A(_01078_),
    .B(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__nand2_1 _31953_ (.A(_01078_),
    .B(_03735_),
    .Y(_03737_));
 sky130_fd_sc_hd__nor2_1 _31954_ (.A(net306),
    .B(\delay_line[34][13] ),
    .Y(_03738_));
 sky130_fd_sc_hd__and2_1 _31955_ (.A(net306),
    .B(\delay_line[34][13] ),
    .X(_03739_));
 sky130_fd_sc_hd__or4bb_2 _31956_ (.A(_03738_),
    .B(_03739_),
    .C_N(_24880_),
    .D_N(net305),
    .X(_03740_));
 sky130_fd_sc_hd__a2bb2o_1 _31957_ (.A1_N(_03738_),
    .A2_N(_03739_),
    .B1(_24880_),
    .B2(_02883_),
    .X(_03741_));
 sky130_fd_sc_hd__a22o_1 _31958_ (.A1(_03736_),
    .A2(_03737_),
    .B1(_03740_),
    .B2(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__nand4_1 _31959_ (.A(_03736_),
    .B(_03737_),
    .C(_03740_),
    .D(_03741_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand2_1 _31960_ (.A(_03742_),
    .B(_03743_),
    .Y(_03745_));
 sky130_fd_sc_hd__nand3_1 _31961_ (.A(_02886_),
    .B(_02890_),
    .C(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__a21oi_2 _31962_ (.A1(_02886_),
    .A2(_02890_),
    .B1(_03745_),
    .Y(_03747_));
 sky130_fd_sc_hd__inv_2 _31963_ (.A(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__xor2_1 _31964_ (.A(_24876_),
    .B(_02882_),
    .X(_03749_));
 sky130_fd_sc_hd__a21o_1 _31965_ (.A1(_03746_),
    .A2(_03748_),
    .B1(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__nand3_1 _31966_ (.A(_03748_),
    .B(_03749_),
    .C(_03746_),
    .Y(_03751_));
 sky130_fd_sc_hd__and3_1 _31967_ (.A(_02891_),
    .B(_02889_),
    .C(_02890_),
    .X(_03752_));
 sky130_fd_sc_hd__a211oi_1 _31968_ (.A1(_03750_),
    .A2(_03751_),
    .B1(_03752_),
    .C1(_02895_),
    .Y(_03753_));
 sky130_fd_sc_hd__o211a_1 _31969_ (.A1(_03752_),
    .A2(_02895_),
    .B1(_03750_),
    .C1(_03751_),
    .X(_03754_));
 sky130_fd_sc_hd__nor2_1 _31970_ (.A(_03753_),
    .B(_03754_),
    .Y(_03756_));
 sky130_fd_sc_hd__xnor2_1 _31971_ (.A(_02879_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__and2b_1 _31972_ (.A_N(_02896_),
    .B(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__a21oi_2 _31973_ (.A1(_02900_),
    .A2(_02899_),
    .B1(_03757_),
    .Y(_03759_));
 sky130_fd_sc_hd__a21o_1 _31974_ (.A1(_03758_),
    .A2(_02899_),
    .B1(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__nand2_1 _31975_ (.A(_02904_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__inv_2 _31976_ (.A(_02904_),
    .Y(_03762_));
 sky130_fd_sc_hd__o21ba_1 _31977_ (.A1(_03762_),
    .A2(_02906_),
    .B1_N(_03760_),
    .X(_03763_));
 sky130_fd_sc_hd__o21bai_1 _31978_ (.A1(_02906_),
    .A2(_03761_),
    .B1_N(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__inv_2 _31979_ (.A(_02861_),
    .Y(_03765_));
 sky130_fd_sc_hd__nor2_1 _31980_ (.A(_03765_),
    .B(_02862_),
    .Y(_03767_));
 sky130_fd_sc_hd__buf_1 _31981_ (.A(_20666_),
    .X(_03768_));
 sky130_fd_sc_hd__clkbuf_2 _31982_ (.A(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__a21oi_1 _31983_ (.A1(_17825_),
    .A2(_01164_),
    .B1(_02851_),
    .Y(_03770_));
 sky130_fd_sc_hd__a31o_1 _31984_ (.A1(_17825_),
    .A2(_02836_),
    .A3(_03769_),
    .B1(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__nor2_1 _31985_ (.A(_02840_),
    .B(_02848_),
    .Y(_03772_));
 sky130_fd_sc_hd__nor2_1 _31986_ (.A(_03768_),
    .B(_23357_),
    .Y(_03773_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _31987_ (.A(\delay_line[33][12] ),
    .X(_03774_));
 sky130_fd_sc_hd__nand3b_2 _31988_ (.A_N(_23347_),
    .B(_24921_),
    .C(net311),
    .Y(_03775_));
 sky130_fd_sc_hd__o21bai_1 _31989_ (.A1(_23347_),
    .A2(_23358_),
    .B1_N(net311),
    .Y(_03776_));
 sky130_fd_sc_hd__o2111a_1 _31990_ (.A1(_03772_),
    .A2(_03773_),
    .B1(_03774_),
    .C1(_03775_),
    .D1(_03776_),
    .X(_03778_));
 sky130_fd_sc_hd__a21oi_1 _31991_ (.A1(_23364_),
    .A2(_03768_),
    .B1(_18651_),
    .Y(_03779_));
 sky130_fd_sc_hd__buf_1 _31992_ (.A(_19574_),
    .X(_03780_));
 sky130_fd_sc_hd__a311o_1 _31993_ (.A1(_18651_),
    .A2(_23364_),
    .A3(_03768_),
    .B1(_17823_),
    .C1(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__and3_1 _31994_ (.A(_18651_),
    .B(_23364_),
    .C(_03768_),
    .X(_03782_));
 sky130_fd_sc_hd__o22ai_1 _31995_ (.A1(_03780_),
    .A2(_17823_),
    .B1(_03779_),
    .B2(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__o21ai_1 _31996_ (.A1(_03779_),
    .A2(_03781_),
    .B1(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__a21boi_1 _31997_ (.A1(_03775_),
    .A2(_03776_),
    .B1_N(_02844_),
    .Y(_03785_));
 sky130_fd_sc_hd__or3_1 _31998_ (.A(_03778_),
    .B(_03784_),
    .C(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__o21ai_1 _31999_ (.A1(_03785_),
    .A2(_03778_),
    .B1(_03784_),
    .Y(_03787_));
 sky130_fd_sc_hd__a211o_1 _32000_ (.A1(_03786_),
    .A2(_03787_),
    .B1(_02856_),
    .C1(_02857_),
    .X(_03789_));
 sky130_fd_sc_hd__o211ai_2 _32001_ (.A1(_02856_),
    .A2(_02857_),
    .B1(_03786_),
    .C1(_03787_),
    .Y(_03790_));
 sky130_fd_sc_hd__nand3_1 _32002_ (.A(_03771_),
    .B(_03789_),
    .C(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__a21o_1 _32003_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03771_),
    .X(_03792_));
 sky130_fd_sc_hd__nand2_1 _32004_ (.A(_03791_),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__xnor2_1 _32005_ (.A(_03767_),
    .B(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__nor2_1 _32006_ (.A(_02864_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__and2_1 _32007_ (.A(_02864_),
    .B(_03794_),
    .X(_03796_));
 sky130_fd_sc_hd__nor2_1 _32008_ (.A(_03795_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__o21bai_2 _32009_ (.A1(_02869_),
    .A2(_02871_),
    .B1_N(_02868_),
    .Y(_03798_));
 sky130_fd_sc_hd__xor2_1 _32010_ (.A(_03797_),
    .B(_03798_),
    .X(_03800_));
 sky130_fd_sc_hd__xnor2_1 _32011_ (.A(_01146_),
    .B(_02830_),
    .Y(_03801_));
 sky130_fd_sc_hd__xor2_1 _32012_ (.A(_24948_),
    .B(_24986_),
    .X(_03802_));
 sky130_fd_sc_hd__a21oi_1 _32013_ (.A1(_23413_),
    .A2(_23409_),
    .B1(_24946_),
    .Y(_03803_));
 sky130_fd_sc_hd__o2bb2ai_1 _32014_ (.A1_N(_01154_),
    .A2_N(_01151_),
    .B1(_03802_),
    .B2(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__a21oi_1 _32015_ (.A1(_03804_),
    .A2(_01152_),
    .B1(_02790_),
    .Y(_03805_));
 sky130_fd_sc_hd__and4_1 _32016_ (.A(_02830_),
    .B(_01144_),
    .C(_01142_),
    .D(_01110_),
    .X(_03806_));
 sky130_fd_sc_hd__o21bai_2 _32017_ (.A1(_03801_),
    .A2(_03805_),
    .B1_N(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__clkbuf_2 _32018_ (.A(_02828_),
    .X(_03808_));
 sky130_fd_sc_hd__buf_1 _32019_ (.A(_02793_),
    .X(_03809_));
 sky130_fd_sc_hd__buf_1 _32020_ (.A(\delay_line[32][13] ),
    .X(_03811_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32021_ (.A(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__o21ai_1 _32022_ (.A1(_03809_),
    .A2(_03811_),
    .B1(_01113_),
    .Y(_03813_));
 sky130_fd_sc_hd__a21oi_1 _32023_ (.A1(_03809_),
    .A2(_03812_),
    .B1(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__nand2_1 _32024_ (.A(_03809_),
    .B(_03812_),
    .Y(_03815_));
 sky130_fd_sc_hd__or2_1 _32025_ (.A(_02793_),
    .B(_03811_),
    .X(_03816_));
 sky130_fd_sc_hd__a21oi_1 _32026_ (.A1(_03815_),
    .A2(_03816_),
    .B1(_01113_),
    .Y(_03817_));
 sky130_fd_sc_hd__a211o_2 _32027_ (.A1(_02794_),
    .A2(_02796_),
    .B1(_03814_),
    .C1(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__o211ai_2 _32028_ (.A1(_03814_),
    .A2(_03817_),
    .B1(_02794_),
    .C1(_02796_),
    .Y(_03819_));
 sky130_fd_sc_hd__nand3_2 _32029_ (.A(_03818_),
    .B(_03819_),
    .C(_02795_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21o_1 _32030_ (.A1(_03818_),
    .A2(_03819_),
    .B1(_02795_),
    .X(_03822_));
 sky130_fd_sc_hd__o211a_1 _32031_ (.A1(_02803_),
    .A2(_02804_),
    .B1(_03820_),
    .C1(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__or2_1 _32032_ (.A(_01132_),
    .B(_24969_),
    .X(_03824_));
 sky130_fd_sc_hd__nand2_1 _32033_ (.A(_24969_),
    .B(_01132_),
    .Y(_03825_));
 sky130_fd_sc_hd__clkbuf_2 _32034_ (.A(_20699_),
    .X(_03826_));
 sky130_fd_sc_hd__nand4_2 _32035_ (.A(_19611_),
    .B(_03824_),
    .C(_03825_),
    .D(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__a22o_1 _32036_ (.A1(_19611_),
    .A2(_03826_),
    .B1(_03824_),
    .B2(_03825_),
    .X(_03828_));
 sky130_fd_sc_hd__nand2_1 _32037_ (.A(_03827_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__a211oi_1 _32038_ (.A1(_03820_),
    .A2(_03822_),
    .B1(_02803_),
    .C1(_02804_),
    .Y(_03830_));
 sky130_fd_sc_hd__nor3_2 _32039_ (.A(_03823_),
    .B(_03829_),
    .C(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__o2bb2a_1 _32040_ (.A1_N(_03827_),
    .A2_N(_03828_),
    .B1(_03830_),
    .B2(_03823_),
    .X(_03833_));
 sky130_fd_sc_hd__inv_2 _32041_ (.A(_02819_),
    .Y(_03834_));
 sky130_fd_sc_hd__o211a_1 _32042_ (.A1(_03831_),
    .A2(_03833_),
    .B1(_02814_),
    .C1(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__a211oi_2 _32043_ (.A1(_02814_),
    .A2(_03834_),
    .B1(_03831_),
    .C1(_03833_),
    .Y(_03836_));
 sky130_fd_sc_hd__nor2_1 _32044_ (.A(_03835_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__a21oi_1 _32045_ (.A1(_02826_),
    .A2(_02817_),
    .B1(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__and3_1 _32046_ (.A(_02826_),
    .B(_02817_),
    .C(_03837_),
    .X(_03839_));
 sky130_fd_sc_hd__o221a_1 _32047_ (.A1(_02822_),
    .A2(_02791_),
    .B1(_03838_),
    .B2(_03839_),
    .C1(_02823_),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _32048_ (.A(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__o21a_1 _32049_ (.A1(_02791_),
    .A2(_02822_),
    .B1(_02823_),
    .X(_03842_));
 sky130_fd_sc_hd__or3_4 _32050_ (.A(_03842_),
    .B(_03839_),
    .C(_03838_),
    .X(_03844_));
 sky130_fd_sc_hd__a21oi_2 _32051_ (.A1(_03841_),
    .A2(_03844_),
    .B1(_03808_),
    .Y(_03845_));
 sky130_fd_sc_hd__a21oi_1 _32052_ (.A1(_03808_),
    .A2(_03841_),
    .B1(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__xor2_2 _32053_ (.A(_03807_),
    .B(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__xnor2_1 _32054_ (.A(_03800_),
    .B(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__or2_1 _32055_ (.A(_03764_),
    .B(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__nand2_1 _32056_ (.A(_03764_),
    .B(_03848_),
    .Y(_03850_));
 sky130_fd_sc_hd__and2b_2 _32057_ (.A_N(_02085_),
    .B(_02124_),
    .X(_03851_));
 sky130_fd_sc_hd__a211oi_2 _32058_ (.A1(_03849_),
    .A2(_03850_),
    .B1(_03851_),
    .C1(_02165_),
    .Y(_03852_));
 sky130_fd_sc_hd__o211a_2 _32059_ (.A1(_03851_),
    .A2(_02165_),
    .B1(_03849_),
    .C1(_03850_),
    .X(_03853_));
 sky130_fd_sc_hd__o221a_1 _32060_ (.A1(_02875_),
    .A2(_02908_),
    .B1(_03852_),
    .B2(_03853_),
    .C1(_02874_),
    .X(_03855_));
 sky130_fd_sc_hd__or3b_1 _32061_ (.A(_02875_),
    .B(_02906_),
    .C_N(_02907_),
    .X(_03856_));
 sky130_fd_sc_hd__a211oi_4 _32062_ (.A1(_02874_),
    .A2(_03856_),
    .B1(_03852_),
    .C1(_03853_),
    .Y(_03857_));
 sky130_fd_sc_hd__or3_1 _32063_ (.A(_03734_),
    .B(_03855_),
    .C(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__o21ai_1 _32064_ (.A1(_03855_),
    .A2(_03857_),
    .B1(_03734_),
    .Y(_03859_));
 sky130_fd_sc_hd__nand2_1 _32065_ (.A(_03858_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__nand2_1 _32066_ (.A(_03732_),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__or2_1 _32067_ (.A(_03860_),
    .B(_03732_),
    .X(_03862_));
 sky130_fd_sc_hd__nand2_1 _32068_ (.A(_03861_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__nand3_2 _32069_ (.A(_02261_),
    .B(_02263_),
    .C(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__a21oi_4 _32070_ (.A1(_02261_),
    .A2(_02263_),
    .B1(_03863_),
    .Y(_03866_));
 sky130_fd_sc_hd__inv_2 _32071_ (.A(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__and3_2 _32072_ (.A(_03620_),
    .B(_03864_),
    .C(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__a21oi_2 _32073_ (.A1(_03864_),
    .A2(_03867_),
    .B1(_03620_),
    .Y(_03869_));
 sky130_fd_sc_hd__and2b_1 _32074_ (.A_N(_02265_),
    .B(_02676_),
    .X(_03870_));
 sky130_fd_sc_hd__a21oi_2 _32075_ (.A1(_02266_),
    .A2(_02675_),
    .B1(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__o21bai_2 _32076_ (.A1(_24844_),
    .A2(_24847_),
    .B1_N(_24845_),
    .Y(_03872_));
 sky130_fd_sc_hd__and4b_1 _32077_ (.A_N(_02528_),
    .B(_00863_),
    .C(_03872_),
    .D(_02529_),
    .X(_03873_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32078_ (.A(_20630_),
    .X(_03874_));
 sky130_fd_sc_hd__o21a_1 _32079_ (.A1(_21517_),
    .A2(_23024_),
    .B1(_20630_),
    .X(_03875_));
 sky130_fd_sc_hd__o21bai_1 _32080_ (.A1(_03874_),
    .A2(_02487_),
    .B1_N(_03875_),
    .Y(_03877_));
 sky130_fd_sc_hd__and2_2 _32081_ (.A(net383),
    .B(_24819_),
    .X(_03878_));
 sky130_fd_sc_hd__o21ai_4 _32082_ (.A1(_23023_),
    .A2(_24819_),
    .B1(_21516_),
    .Y(_03879_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32083_ (.A(\delay_line[16][12] ),
    .X(_03880_));
 sky130_fd_sc_hd__nor2_1 _32084_ (.A(_23023_),
    .B(_24821_),
    .Y(_03881_));
 sky130_fd_sc_hd__o21bai_2 _32085_ (.A1(_03878_),
    .A2(_03881_),
    .B1_N(_21517_),
    .Y(_03882_));
 sky130_fd_sc_hd__o211a_1 _32086_ (.A1(_03878_),
    .A2(_03879_),
    .B1(_03880_),
    .C1(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__a21o_1 _32087_ (.A1(_23024_),
    .A2(_24821_),
    .B1(_03879_),
    .X(_03884_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32088_ (.A(_03880_),
    .X(_03885_));
 sky130_fd_sc_hd__a21oi_1 _32089_ (.A1(_03884_),
    .A2(_03882_),
    .B1(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__and3_1 _32090_ (.A(_02488_),
    .B(_02494_),
    .C(_02492_),
    .X(_03888_));
 sky130_fd_sc_hd__o21ai_1 _32091_ (.A1(_03883_),
    .A2(_03886_),
    .B1(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__o211ai_2 _32092_ (.A1(_03878_),
    .A2(_03879_),
    .B1(_03880_),
    .C1(_03882_),
    .Y(_03890_));
 sky130_fd_sc_hd__a21o_1 _32093_ (.A1(_03884_),
    .A2(_03882_),
    .B1(_03880_),
    .X(_03891_));
 sky130_fd_sc_hd__nand3_1 _32094_ (.A(_02500_),
    .B(_03890_),
    .C(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand3_1 _32095_ (.A(_03877_),
    .B(_03889_),
    .C(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__nand3_1 _32096_ (.A(_03891_),
    .B(_03888_),
    .C(_03890_),
    .Y(_03894_));
 sky130_fd_sc_hd__o21ai_1 _32097_ (.A1(_03883_),
    .A2(_03886_),
    .B1(_02500_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand3b_2 _32098_ (.A_N(_03877_),
    .B(_03894_),
    .C(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__a21oi_1 _32099_ (.A1(_02500_),
    .A2(_02495_),
    .B1(_00831_),
    .Y(_03897_));
 sky130_fd_sc_hd__o21ai_1 _32100_ (.A1(_02485_),
    .A2(_03897_),
    .B1(_02504_),
    .Y(_03899_));
 sky130_fd_sc_hd__a21o_1 _32101_ (.A1(_03893_),
    .A2(_03896_),
    .B1(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32102_ (.A(_19441_),
    .X(_03901_));
 sky130_fd_sc_hd__o211a_1 _32103_ (.A1(_03874_),
    .A2(_21518_),
    .B1(_16601_),
    .C1(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__nand2_1 _32104_ (.A(_16667_),
    .B(_00837_),
    .Y(_03903_));
 sky130_fd_sc_hd__and2b_1 _32105_ (.A_N(_03902_),
    .B(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__nand3_1 _32106_ (.A(_03899_),
    .B(_03893_),
    .C(_03896_),
    .Y(_03905_));
 sky130_fd_sc_hd__nand3_2 _32107_ (.A(_03900_),
    .B(_03904_),
    .C(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__a21o_1 _32108_ (.A1(_03905_),
    .A2(_03900_),
    .B1(_03904_),
    .X(_03907_));
 sky130_fd_sc_hd__o21ai_1 _32109_ (.A1(_02508_),
    .A2(_02507_),
    .B1(_02516_),
    .Y(_03908_));
 sky130_fd_sc_hd__a21o_1 _32110_ (.A1(_03906_),
    .A2(_03907_),
    .B1(_03908_),
    .X(_03910_));
 sky130_fd_sc_hd__nand3_2 _32111_ (.A(_03908_),
    .B(_03906_),
    .C(_03907_),
    .Y(_03911_));
 sky130_fd_sc_hd__nand3_2 _32112_ (.A(_03910_),
    .B(_03911_),
    .C(_02510_),
    .Y(_03912_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32113_ (.A(_24835_),
    .X(_03913_));
 sky130_fd_sc_hd__a32o_1 _32114_ (.A1(_21536_),
    .A2(_03913_),
    .A3(_24814_),
    .B1(_03910_),
    .B2(_03911_),
    .X(_03914_));
 sky130_fd_sc_hd__nand2_1 _32115_ (.A(_02518_),
    .B(_02523_),
    .Y(_03915_));
 sky130_fd_sc_hd__a21o_1 _32116_ (.A1(_03912_),
    .A2(_03914_),
    .B1(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__nand3_2 _32117_ (.A(_03915_),
    .B(_03912_),
    .C(_03914_),
    .Y(_03917_));
 sky130_fd_sc_hd__o211a_1 _32118_ (.A1(_02528_),
    .A2(_03873_),
    .B1(_03916_),
    .C1(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__and2_1 _32119_ (.A(_03916_),
    .B(_03917_),
    .X(_03919_));
 sky130_fd_sc_hd__a311oi_2 _32120_ (.A1(_00863_),
    .A2(_03872_),
    .A3(_02529_),
    .B1(_03919_),
    .C1(_02528_),
    .Y(_03921_));
 sky130_fd_sc_hd__buf_1 _32121_ (.A(_20589_),
    .X(_03922_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32122_ (.A(_21497_),
    .X(_03923_));
 sky130_fd_sc_hd__a21oi_1 _32123_ (.A1(_03922_),
    .A2(_03923_),
    .B1(_18407_),
    .Y(_03924_));
 sky130_fd_sc_hd__and3_1 _32124_ (.A(_18407_),
    .B(_20589_),
    .C(_21497_),
    .X(_03925_));
 sky130_fd_sc_hd__inv_2 _32125_ (.A(\delay_line[14][12] ),
    .Y(_03926_));
 sky130_fd_sc_hd__nor2_1 _32126_ (.A(_21492_),
    .B(net390),
    .Y(_03927_));
 sky130_fd_sc_hd__and2_1 _32127_ (.A(\delay_line[14][7] ),
    .B(net390),
    .X(_03928_));
 sky130_fd_sc_hd__or3_1 _32128_ (.A(_03926_),
    .B(_03927_),
    .C(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__o21bai_1 _32129_ (.A1(_03927_),
    .A2(_03928_),
    .B1_N(\delay_line[14][12] ),
    .Y(_03930_));
 sky130_fd_sc_hd__nand3b_2 _32130_ (.A_N(_02409_),
    .B(_03929_),
    .C(_03930_),
    .Y(_03932_));
 sky130_fd_sc_hd__inv_2 _32131_ (.A(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__a21boi_1 _32132_ (.A1(_03929_),
    .A2(_03930_),
    .B1_N(_02409_),
    .Y(_03934_));
 sky130_fd_sc_hd__or4_2 _32133_ (.A(_03924_),
    .B(_03925_),
    .C(_03933_),
    .D(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__o22ai_2 _32134_ (.A1(_03924_),
    .A2(_03925_),
    .B1(_03933_),
    .B2(_03934_),
    .Y(_03936_));
 sky130_fd_sc_hd__nor4_1 _32135_ (.A(_02413_),
    .B(_02415_),
    .C(_02419_),
    .D(_02412_),
    .Y(_03937_));
 sky130_fd_sc_hd__a211oi_1 _32136_ (.A1(_03935_),
    .A2(_03936_),
    .B1(_02419_),
    .C1(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__o211ai_2 _32137_ (.A1(_02419_),
    .A2(net229),
    .B1(_03935_),
    .C1(_03936_),
    .Y(_03939_));
 sky130_fd_sc_hd__inv_2 _32138_ (.A(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__or3b_4 _32139_ (.A(_03938_),
    .B(_03940_),
    .C_N(_02415_),
    .X(_03941_));
 sky130_fd_sc_hd__a2bb2o_1 _32140_ (.A1_N(_03938_),
    .A2_N(_03940_),
    .B1(_16843_),
    .B2(_00745_),
    .X(_03943_));
 sky130_fd_sc_hd__a21bo_1 _32141_ (.A1(_02421_),
    .A2(_00742_),
    .B1_N(_02422_),
    .X(_03944_));
 sky130_fd_sc_hd__a21oi_2 _32142_ (.A1(_03941_),
    .A2(_03943_),
    .B1(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__and3_1 _32143_ (.A(_03944_),
    .B(_03941_),
    .C(_03943_),
    .X(_03946_));
 sky130_fd_sc_hd__or2_2 _32144_ (.A(_03945_),
    .B(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__o21bai_2 _32145_ (.A1(_00761_),
    .A2(_00763_),
    .B1_N(_00762_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2_1 _32146_ (.A(_02424_),
    .B(_02426_),
    .Y(_03949_));
 sky130_fd_sc_hd__a21boi_4 _32147_ (.A1(_03948_),
    .A2(_02427_),
    .B1_N(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__xnor2_4 _32148_ (.A(_03947_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__o22ai_4 _32149_ (.A1(_02471_),
    .A2(_02474_),
    .B1(_02475_),
    .B2(_02479_),
    .Y(_03952_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32150_ (.A(\delay_line[15][13] ),
    .X(_03954_));
 sky130_fd_sc_hd__nor2_1 _32151_ (.A(_00781_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__and2_1 _32152_ (.A(_00781_),
    .B(\delay_line[15][13] ),
    .X(_03956_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32153_ (.A(_02431_),
    .X(_03957_));
 sky130_fd_sc_hd__nand2_1 _32154_ (.A(_24737_),
    .B(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__o21ai_2 _32155_ (.A1(_03955_),
    .A2(_03956_),
    .B1(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__buf_1 _32156_ (.A(_21459_),
    .X(_03960_));
 sky130_fd_sc_hd__nand2_1 _32157_ (.A(_00781_),
    .B(_03954_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand3b_1 _32158_ (.A_N(_03955_),
    .B(_03961_),
    .C(_02430_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand3_1 _32159_ (.A(_03959_),
    .B(_03960_),
    .C(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__a21o_1 _32160_ (.A1(_03962_),
    .A2(_03959_),
    .B1(_21459_),
    .X(_03965_));
 sky130_fd_sc_hd__o2bb2ai_1 _32161_ (.A1_N(_02433_),
    .A2_N(_02437_),
    .B1(_02432_),
    .B2(_02430_),
    .Y(_03966_));
 sky130_fd_sc_hd__nand3_2 _32162_ (.A(_03963_),
    .B(_03965_),
    .C(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__and3_1 _32163_ (.A(_03959_),
    .B(_21459_),
    .C(_03962_),
    .X(_03968_));
 sky130_fd_sc_hd__a21oi_1 _32164_ (.A1(_03962_),
    .A2(_03959_),
    .B1(_03960_),
    .Y(_03969_));
 sky130_fd_sc_hd__o21bai_2 _32165_ (.A1(_03968_),
    .A2(_03969_),
    .B1_N(_03966_),
    .Y(_03970_));
 sky130_fd_sc_hd__buf_1 _32166_ (.A(_21458_),
    .X(_03971_));
 sky130_fd_sc_hd__a21oi_1 _32167_ (.A1(_16689_),
    .A2(_18423_),
    .B1(_03971_),
    .Y(_03972_));
 sky130_fd_sc_hd__and3_1 _32168_ (.A(_16689_),
    .B(_18423_),
    .C(_03971_),
    .X(_03973_));
 sky130_fd_sc_hd__nor2_1 _32169_ (.A(_03972_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand3_2 _32170_ (.A(_03967_),
    .B(_03970_),
    .C(_03974_),
    .Y(_03976_));
 sky130_fd_sc_hd__o2bb2ai_1 _32171_ (.A1_N(_03967_),
    .A2_N(_03970_),
    .B1(_03972_),
    .B2(_03973_),
    .Y(_03977_));
 sky130_fd_sc_hd__nand2_1 _32172_ (.A(_02443_),
    .B(_02456_),
    .Y(_03978_));
 sky130_fd_sc_hd__a21oi_1 _32173_ (.A1(_03976_),
    .A2(_03977_),
    .B1(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__or3b_1 _32174_ (.A(_18429_),
    .B(_19467_),
    .C_N(_07107_),
    .X(_03980_));
 sky130_fd_sc_hd__clkbuf_2 _32175_ (.A(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__nand3_1 _32176_ (.A(_03978_),
    .B(_03976_),
    .C(_03977_),
    .Y(_03982_));
 sky130_fd_sc_hd__nand4b_2 _32177_ (.A_N(_03979_),
    .B(_18413_),
    .C(_03981_),
    .D(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__a21o_1 _32178_ (.A1(_18429_),
    .A2(_19467_),
    .B1(_02448_),
    .X(_03984_));
 sky130_fd_sc_hd__a21boi_1 _32179_ (.A1(_02445_),
    .A2(_03984_),
    .B1_N(_02443_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _32180_ (.A(_03976_),
    .B(_03977_),
    .Y(_03987_));
 sky130_fd_sc_hd__nor2_1 _32181_ (.A(_03985_),
    .B(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__o2bb2ai_1 _32182_ (.A1_N(_18413_),
    .A2_N(_03981_),
    .B1(_03979_),
    .B2(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__o21ai_1 _32183_ (.A1(_02460_),
    .A2(_02465_),
    .B1(_02459_),
    .Y(_03990_));
 sky130_fd_sc_hd__a21o_1 _32184_ (.A1(_03983_),
    .A2(_03989_),
    .B1(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__nand3_1 _32185_ (.A(_03990_),
    .B(_03983_),
    .C(_03989_),
    .Y(_03992_));
 sky130_fd_sc_hd__nand2_1 _32186_ (.A(_03991_),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__xnor2_1 _32187_ (.A(_02467_),
    .B(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__o21bai_1 _32188_ (.A1(_02470_),
    .A2(_02473_),
    .B1_N(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__o211ai_1 _32189_ (.A1(_00800_),
    .A2(_02463_),
    .B1(_02472_),
    .C1(_03994_),
    .Y(_03996_));
 sky130_fd_sc_hd__and2_1 _32190_ (.A(_03995_),
    .B(_03996_),
    .X(_03998_));
 sky130_fd_sc_hd__xnor2_2 _32191_ (.A(_03952_),
    .B(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__xnor2_1 _32192_ (.A(_03951_),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__o21ai_2 _32193_ (.A1(_03918_),
    .A2(_03921_),
    .B1(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__or3_2 _32194_ (.A(_03918_),
    .B(_03921_),
    .C(_04000_),
    .X(_04002_));
 sky130_fd_sc_hd__a21bo_1 _32195_ (.A1(_02531_),
    .A2(_02482_),
    .B1_N(_02532_),
    .X(_04003_));
 sky130_fd_sc_hd__a21o_1 _32196_ (.A1(_04001_),
    .A2(_04002_),
    .B1(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__nand3_4 _32197_ (.A(_04003_),
    .B(_04001_),
    .C(_04002_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand2_2 _32198_ (.A(_04004_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__and3_1 _32199_ (.A(_02648_),
    .B(_02643_),
    .C(_02647_),
    .X(_04007_));
 sky130_fd_sc_hd__a31oi_1 _32200_ (.A1(_02649_),
    .A2(_07525_),
    .A3(_02650_),
    .B1(_04007_),
    .Y(_04009_));
 sky130_fd_sc_hd__and3_1 _32201_ (.A(_18388_),
    .B(_07525_),
    .C(_24704_),
    .X(_04010_));
 sky130_fd_sc_hd__o21ai_1 _32202_ (.A1(_24704_),
    .A2(_18388_),
    .B1(_19395_),
    .Y(_04011_));
 sky130_fd_sc_hd__nand3_1 _32203_ (.A(_16338_),
    .B(_18384_),
    .C(_19391_),
    .Y(_04012_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32204_ (.A(\delay_line[18][12] ),
    .X(_04013_));
 sky130_fd_sc_hd__nor2_1 _32205_ (.A(_22925_),
    .B(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__nand2_1 _32206_ (.A(_22931_),
    .B(_04013_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand3b_2 _32207_ (.A_N(_04014_),
    .B(_02639_),
    .C(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__and2_1 _32208_ (.A(_22925_),
    .B(\delay_line[18][12] ),
    .X(_04017_));
 sky130_fd_sc_hd__o21ai_1 _32209_ (.A1(_04017_),
    .A2(_04014_),
    .B1(_02636_),
    .Y(_04018_));
 sky130_fd_sc_hd__nand4_2 _32210_ (.A(_04011_),
    .B(_04012_),
    .C(_04016_),
    .D(_04018_),
    .Y(_04020_));
 sky130_fd_sc_hd__a22o_1 _32211_ (.A1(_04011_),
    .A2(_04012_),
    .B1(_04016_),
    .B2(_04018_),
    .X(_04021_));
 sky130_fd_sc_hd__o21ai_1 _32212_ (.A1(_02646_),
    .A2(_02644_),
    .B1(_02637_),
    .Y(_04022_));
 sky130_fd_sc_hd__a21oi_1 _32213_ (.A1(_04020_),
    .A2(_04021_),
    .B1(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__and3_1 _32214_ (.A(_04022_),
    .B(_04020_),
    .C(_04021_),
    .X(_04024_));
 sky130_fd_sc_hd__nor4_2 _32215_ (.A(_16338_),
    .B(_04010_),
    .C(_04023_),
    .D(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__o22a_1 _32216_ (.A1(_16349_),
    .A2(_04010_),
    .B1(_04023_),
    .B2(_04024_),
    .X(_04026_));
 sky130_fd_sc_hd__or3_2 _32217_ (.A(_04009_),
    .B(_04025_),
    .C(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__o21ai_1 _32218_ (.A1(_04025_),
    .A2(_04026_),
    .B1(_04009_),
    .Y(_04028_));
 sky130_fd_sc_hd__and3_1 _32219_ (.A(_16349_),
    .B(_07536_),
    .C(_01688_),
    .X(_04029_));
 sky130_fd_sc_hd__nand3_1 _32220_ (.A(_04027_),
    .B(_04028_),
    .C(_04029_),
    .Y(_04031_));
 sky130_fd_sc_hd__a32o_1 _32221_ (.A1(_01688_),
    .A2(_16349_),
    .A3(_07536_),
    .B1(_04027_),
    .B2(_04028_),
    .X(_04032_));
 sky130_fd_sc_hd__nand2_1 _32222_ (.A(_02654_),
    .B(_02661_),
    .Y(_04033_));
 sky130_fd_sc_hd__a21oi_2 _32223_ (.A1(_04031_),
    .A2(_04032_),
    .B1(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__and3_1 _32224_ (.A(_04033_),
    .B(_04031_),
    .C(_04032_),
    .X(_04035_));
 sky130_fd_sc_hd__a211oi_4 _32225_ (.A1(_02662_),
    .A2(_02660_),
    .B1(_04034_),
    .C1(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__o211a_1 _32226_ (.A1(_04034_),
    .A2(_04035_),
    .B1(_02662_),
    .C1(_02660_),
    .X(_04037_));
 sky130_fd_sc_hd__o21ai_1 _32227_ (.A1(_07426_),
    .A2(_20575_),
    .B1(_07470_),
    .Y(_04038_));
 sky130_fd_sc_hd__nand2_1 _32228_ (.A(_22956_),
    .B(_00668_),
    .Y(_04039_));
 sky130_fd_sc_hd__o2111ai_4 _32229_ (.A1(_19400_),
    .A2(_18368_),
    .B1(_20554_),
    .C1(_20552_),
    .D1(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__a22o_1 _32230_ (.A1(_20552_),
    .A2(_20554_),
    .B1(_04039_),
    .B2(_18372_),
    .X(_04042_));
 sky130_fd_sc_hd__buf_2 _32231_ (.A(_02587_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_1 _32232_ (.A(_02586_),
    .B(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__clkbuf_2 _32233_ (.A(\delay_line[19][12] ),
    .X(_04045_));
 sky130_fd_sc_hd__nand2_2 _32234_ (.A(_00658_),
    .B(_02585_),
    .Y(_04046_));
 sky130_fd_sc_hd__nor2_2 _32235_ (.A(_02585_),
    .B(\delay_line[19][12] ),
    .Y(_04047_));
 sky130_fd_sc_hd__and2_1 _32236_ (.A(\delay_line[19][11] ),
    .B(\delay_line[19][12] ),
    .X(_04048_));
 sky130_fd_sc_hd__o21ai_2 _32237_ (.A1(_04047_),
    .A2(_04048_),
    .B1(_04046_),
    .Y(_04049_));
 sky130_fd_sc_hd__o211ai_4 _32238_ (.A1(_04045_),
    .A2(_04046_),
    .B1(_21382_),
    .C1(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__or2_1 _32239_ (.A(_04045_),
    .B(_04046_),
    .X(_04051_));
 sky130_fd_sc_hd__a21o_1 _32240_ (.A1(_04049_),
    .A2(_04051_),
    .B1(_21382_),
    .X(_04053_));
 sky130_fd_sc_hd__o211ai_4 _32241_ (.A1(_04044_),
    .A2(_02597_),
    .B1(_04050_),
    .C1(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__clkbuf_2 _32242_ (.A(_21381_),
    .X(_04055_));
 sky130_fd_sc_hd__a21oi_1 _32243_ (.A1(_04049_),
    .A2(_04051_),
    .B1(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__and3_1 _32244_ (.A(_04049_),
    .B(_04051_),
    .C(_21382_),
    .X(_04057_));
 sky130_fd_sc_hd__o221ai_4 _32245_ (.A1(_04043_),
    .A2(_02586_),
    .B1(_04056_),
    .B2(_04057_),
    .C1(_02592_),
    .Y(_04058_));
 sky130_fd_sc_hd__nand4_1 _32246_ (.A(_04040_),
    .B(_04042_),
    .C(_04054_),
    .D(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__a22o_1 _32247_ (.A1(_04040_),
    .A2(_04042_),
    .B1(_04054_),
    .B2(_04058_),
    .X(_04060_));
 sky130_fd_sc_hd__nand4_1 _32248_ (.A(_02596_),
    .B(_02610_),
    .C(_04059_),
    .D(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__a22o_1 _32249_ (.A1(_02596_),
    .A2(_02610_),
    .B1(_04059_),
    .B2(_04060_),
    .X(_04062_));
 sky130_fd_sc_hd__o22a_1 _32250_ (.A1(_07459_),
    .A2(_20569_),
    .B1(_19401_),
    .B2(_19403_),
    .X(_04064_));
 sky130_fd_sc_hd__a21oi_1 _32251_ (.A1(_07470_),
    .A2(_20569_),
    .B1(_18380_),
    .Y(_04065_));
 sky130_fd_sc_hd__or2_1 _32252_ (.A(_04064_),
    .B(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__a21oi_1 _32253_ (.A1(_04061_),
    .A2(_04062_),
    .B1(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__nand2_1 _32254_ (.A(_02613_),
    .B(_02618_),
    .Y(_04068_));
 sky130_fd_sc_hd__and3_1 _32255_ (.A(_04066_),
    .B(_04061_),
    .C(_04062_),
    .X(_04069_));
 sky130_fd_sc_hd__nor3_1 _32256_ (.A(_04067_),
    .B(_04068_),
    .C(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__o2bb2a_1 _32257_ (.A1_N(_02613_),
    .A2_N(_02618_),
    .B1(_04069_),
    .B2(_04067_),
    .X(_04071_));
 sky130_fd_sc_hd__nor4_1 _32258_ (.A(_18373_),
    .B(_04038_),
    .C(_04070_),
    .D(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__o22a_1 _32259_ (.A1(_18373_),
    .A2(_04038_),
    .B1(_04070_),
    .B2(_04071_),
    .X(_04073_));
 sky130_fd_sc_hd__nor2_1 _32260_ (.A(_02621_),
    .B(_02622_),
    .Y(_04075_));
 sky130_fd_sc_hd__o21ai_1 _32261_ (.A1(net132),
    .A2(_04073_),
    .B1(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__or3_1 _32262_ (.A(_04075_),
    .B(net132),
    .C(_04073_),
    .X(_04077_));
 sky130_fd_sc_hd__o21ai_1 _32263_ (.A1(_02628_),
    .A2(_02583_),
    .B1(_02625_),
    .Y(_04078_));
 sky130_fd_sc_hd__and3_2 _32264_ (.A(_04076_),
    .B(_04077_),
    .C(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__or2_1 _32265_ (.A(_04075_),
    .B(net132),
    .X(_04080_));
 sky130_fd_sc_hd__o21ai_1 _32266_ (.A1(_04073_),
    .A2(_04080_),
    .B1(_04076_),
    .Y(_04081_));
 sky130_fd_sc_hd__o311a_2 _32267_ (.A1(net140),
    .A2(_02624_),
    .A3(_02626_),
    .B1(_02630_),
    .C1(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__o22ai_4 _32268_ (.A1(_04036_),
    .A2(_04037_),
    .B1(_04079_),
    .B2(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__or4_4 _32269_ (.A(_04036_),
    .B(_04037_),
    .C(_04079_),
    .D(_04082_),
    .X(_04084_));
 sky130_fd_sc_hd__o22a_1 _32270_ (.A1(_07591_),
    .A2(_18350_),
    .B1(_19418_),
    .B2(_19419_),
    .X(_04086_));
 sky130_fd_sc_hd__o21bai_1 _32271_ (.A1(_18361_),
    .A2(_00605_),
    .B1_N(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__o211ai_2 _32272_ (.A1(_02553_),
    .A2(_02554_),
    .B1(_02549_),
    .C1(_02551_),
    .Y(_04088_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32273_ (.A(_21423_),
    .X(_04089_));
 sky130_fd_sc_hd__buf_1 _32274_ (.A(_21412_),
    .X(_04090_));
 sky130_fd_sc_hd__a21boi_1 _32275_ (.A1(_18352_),
    .A2(_04090_),
    .B1_N(_18356_),
    .Y(_04091_));
 sky130_fd_sc_hd__o211ai_2 _32276_ (.A1(_04089_),
    .A2(_20517_),
    .B1(_20518_),
    .C1(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__a21o_1 _32277_ (.A1(_20518_),
    .A2(_20519_),
    .B1(_04091_),
    .X(_04093_));
 sky130_fd_sc_hd__buf_2 _32278_ (.A(net357),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_2 _32279_ (.A(\delay_line[21][11] ),
    .X(_04095_));
 sky130_fd_sc_hd__nand2_4 _32280_ (.A(_00613_),
    .B(_04095_),
    .Y(_04097_));
 sky130_fd_sc_hd__clkbuf_2 _32281_ (.A(_21418_),
    .X(_04098_));
 sky130_fd_sc_hd__nor2_2 _32282_ (.A(_04095_),
    .B(net357),
    .Y(_04099_));
 sky130_fd_sc_hd__and2_1 _32283_ (.A(_04095_),
    .B(net357),
    .X(_04100_));
 sky130_fd_sc_hd__o21ai_2 _32284_ (.A1(_04099_),
    .A2(_04100_),
    .B1(_04097_),
    .Y(_04101_));
 sky130_fd_sc_hd__o211ai_4 _32285_ (.A1(_04094_),
    .A2(_04097_),
    .B1(_04098_),
    .C1(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__clkbuf_2 _32286_ (.A(net357),
    .X(_04103_));
 sky130_fd_sc_hd__or2_1 _32287_ (.A(_04103_),
    .B(_04097_),
    .X(_04104_));
 sky130_fd_sc_hd__a21o_1 _32288_ (.A1(_04101_),
    .A2(_04104_),
    .B1(_04098_),
    .X(_04105_));
 sky130_fd_sc_hd__buf_1 _32289_ (.A(_04095_),
    .X(_04106_));
 sky130_fd_sc_hd__a2bb2o_1 _32290_ (.A1_N(_04106_),
    .A2_N(_02542_),
    .B1(_21423_),
    .B2(_02543_),
    .X(_04108_));
 sky130_fd_sc_hd__nand3_1 _32291_ (.A(_04102_),
    .B(_04105_),
    .C(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__a21o_1 _32292_ (.A1(_04102_),
    .A2(_04105_),
    .B1(_04108_),
    .X(_04110_));
 sky130_fd_sc_hd__nand4_1 _32293_ (.A(_04092_),
    .B(_04093_),
    .C(_04109_),
    .D(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__a22o_1 _32294_ (.A1(_04092_),
    .A2(_04093_),
    .B1(_04109_),
    .B2(_04110_),
    .X(_04112_));
 sky130_fd_sc_hd__nand4_1 _32295_ (.A(_02549_),
    .B(_04088_),
    .C(_04111_),
    .D(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__a22o_1 _32296_ (.A1(_02549_),
    .A2(_04088_),
    .B1(_04111_),
    .B2(_04112_),
    .X(_04114_));
 sky130_fd_sc_hd__and3_1 _32297_ (.A(_04087_),
    .B(_04113_),
    .C(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__a21oi_1 _32298_ (.A1(_04113_),
    .A2(_04114_),
    .B1(_04087_),
    .Y(_04116_));
 sky130_fd_sc_hd__nand2_1 _32299_ (.A(_02562_),
    .B(_02570_),
    .Y(_04117_));
 sky130_fd_sc_hd__or3_1 _32300_ (.A(_04115_),
    .B(_04116_),
    .C(_04117_),
    .X(_04119_));
 sky130_fd_sc_hd__o21ai_1 _32301_ (.A1(_04115_),
    .A2(_04116_),
    .B1(_04117_),
    .Y(_04120_));
 sky130_fd_sc_hd__and3_1 _32302_ (.A(_04119_),
    .B(_04120_),
    .C(_18362_),
    .X(_04121_));
 sky130_fd_sc_hd__a21oi_1 _32303_ (.A1(_04119_),
    .A2(_04120_),
    .B1(_18362_),
    .Y(_04122_));
 sky130_fd_sc_hd__a211oi_1 _32304_ (.A1(_02571_),
    .A2(_02573_),
    .B1(_04121_),
    .C1(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__o221a_1 _32305_ (.A1(_16536_),
    .A2(_02572_),
    .B1(_04121_),
    .B2(_04122_),
    .C1(_02571_),
    .X(_04124_));
 sky130_fd_sc_hd__nor2_1 _32306_ (.A(_04123_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__a21boi_2 _32307_ (.A1(_02580_),
    .A2(_02577_),
    .B1_N(_02576_),
    .Y(_04126_));
 sky130_fd_sc_hd__xnor2_2 _32308_ (.A(_04125_),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__a21o_1 _32309_ (.A1(_04083_),
    .A2(_04084_),
    .B1(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__nand3_4 _32310_ (.A(_04084_),
    .B(_04127_),
    .C(_04083_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand3b_4 _32311_ (.A_N(_04006_),
    .B(_04128_),
    .C(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__a21bo_1 _32312_ (.A1(_04128_),
    .A2(_04130_),
    .B1_N(_04006_),
    .X(_04132_));
 sky130_fd_sc_hd__o211ai_4 _32313_ (.A1(_02538_),
    .A2(_02670_),
    .B1(_04131_),
    .C1(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__inv_2 _32314_ (.A(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__and2_1 _32315_ (.A(_02669_),
    .B(_02668_),
    .X(_04135_));
 sky130_fd_sc_hd__a221oi_4 _32316_ (.A1(_04135_),
    .A2(_02539_),
    .B1(_04131_),
    .B2(_04132_),
    .C1(_02538_),
    .Y(_04136_));
 sky130_fd_sc_hd__nor2_1 _32317_ (.A(_04134_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__o21a_1 _32318_ (.A1(_02358_),
    .A2(_02393_),
    .B1(_02395_),
    .X(_04138_));
 sky130_fd_sc_hd__a22o_1 _32319_ (.A1(_00500_),
    .A2(_00503_),
    .B1(_02306_),
    .B2(_02307_),
    .X(_04139_));
 sky130_fd_sc_hd__o21ai_4 _32320_ (.A1(_02309_),
    .A2(_02269_),
    .B1(_04139_),
    .Y(_04141_));
 sky130_fd_sc_hd__nor2_1 _32321_ (.A(_00474_),
    .B(\delay_line[25][13] ),
    .Y(_04142_));
 sky130_fd_sc_hd__and2_1 _32322_ (.A(_00474_),
    .B(\delay_line[25][13] ),
    .X(_04143_));
 sky130_fd_sc_hd__nor2_1 _32323_ (.A(_04142_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__nand2_1 _32324_ (.A(_02277_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__o21ai_2 _32325_ (.A1(_04142_),
    .A2(_04143_),
    .B1(_02279_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand3_1 _32326_ (.A(_04145_),
    .B(_04146_),
    .C(_21570_),
    .Y(_04147_));
 sky130_fd_sc_hd__a21o_1 _32327_ (.A1(_04145_),
    .A2(_04146_),
    .B1(_21570_),
    .X(_04148_));
 sky130_fd_sc_hd__nand2_1 _32328_ (.A(_02280_),
    .B(_02281_),
    .Y(_04149_));
 sky130_fd_sc_hd__nand3_1 _32329_ (.A(_04147_),
    .B(_04148_),
    .C(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__a21o_1 _32330_ (.A1(_04147_),
    .A2(_04148_),
    .B1(_04149_),
    .X(_04152_));
 sky130_fd_sc_hd__xor2_1 _32331_ (.A(_00484_),
    .B(_02273_),
    .X(_04153_));
 sky130_fd_sc_hd__nand3_1 _32332_ (.A(_04150_),
    .B(_04152_),
    .C(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__a21o_1 _32333_ (.A1(_04150_),
    .A2(_04152_),
    .B1(_04153_),
    .X(_04155_));
 sky130_fd_sc_hd__a31o_1 _32334_ (.A1(_02281_),
    .A2(_02283_),
    .A3(_02284_),
    .B1(_02287_),
    .X(_04156_));
 sky130_fd_sc_hd__a21o_1 _32335_ (.A1(_04154_),
    .A2(_04155_),
    .B1(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__nand3b_2 _32336_ (.A_N(_24507_),
    .B(_00465_),
    .C(_17215_),
    .Y(_04158_));
 sky130_fd_sc_hd__nand3_2 _32337_ (.A(_04156_),
    .B(_04154_),
    .C(_04155_),
    .Y(_04159_));
 sky130_fd_sc_hd__nand4_2 _32338_ (.A(_04157_),
    .B(_18322_),
    .C(_04158_),
    .D(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__inv_2 _32339_ (.A(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__a22oi_2 _32340_ (.A1(_18322_),
    .A2(_04158_),
    .B1(_04157_),
    .B2(_04159_),
    .Y(_04163_));
 sky130_fd_sc_hd__a211oi_2 _32341_ (.A1(_02296_),
    .A2(_02302_),
    .B1(_04161_),
    .C1(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__o211a_1 _32342_ (.A1(_04161_),
    .A2(_04163_),
    .B1(_02296_),
    .C1(_02302_),
    .X(_04165_));
 sky130_fd_sc_hd__nor3_2 _32343_ (.A(_04164_),
    .B(_00470_),
    .C(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__o21a_1 _32344_ (.A1(_04165_),
    .A2(_04164_),
    .B1(_00470_),
    .X(_04167_));
 sky130_fd_sc_hd__a31o_1 _32345_ (.A1(_02298_),
    .A2(_02299_),
    .A3(_02301_),
    .B1(_02272_),
    .X(_04168_));
 sky130_fd_sc_hd__o211a_1 _32346_ (.A1(_04166_),
    .A2(_04167_),
    .B1(_02305_),
    .C1(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__a211oi_1 _32347_ (.A1(_02305_),
    .A2(_04168_),
    .B1(_04166_),
    .C1(_04167_),
    .Y(_04170_));
 sky130_fd_sc_hd__or2_2 _32348_ (.A(_04169_),
    .B(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__xnor2_4 _32349_ (.A(_04141_),
    .B(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32350_ (.A(_02371_),
    .X(_04174_));
 sky130_fd_sc_hd__o21ai_1 _32351_ (.A1(_02360_),
    .A2(_04174_),
    .B1(_00517_),
    .Y(_04175_));
 sky130_fd_sc_hd__nand3_1 _32352_ (.A(_17084_),
    .B(_18316_),
    .C(_00512_),
    .Y(_04176_));
 sky130_fd_sc_hd__buf_1 _32353_ (.A(\delay_line[22][8] ),
    .X(_04177_));
 sky130_fd_sc_hd__nor2_1 _32354_ (.A(_04177_),
    .B(\delay_line[22][12] ),
    .Y(_04178_));
 sky130_fd_sc_hd__buf_1 _32355_ (.A(\delay_line[22][12] ),
    .X(_04179_));
 sky130_fd_sc_hd__nand2_1 _32356_ (.A(_04177_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__nand3b_2 _32357_ (.A_N(_04178_),
    .B(_02368_),
    .C(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__and2_1 _32358_ (.A(_04177_),
    .B(\delay_line[22][12] ),
    .X(_04182_));
 sky130_fd_sc_hd__o21ai_1 _32359_ (.A1(_04182_),
    .A2(_04178_),
    .B1(_02365_),
    .Y(_04183_));
 sky130_fd_sc_hd__nand4_2 _32360_ (.A(_04175_),
    .B(_04176_),
    .C(_04181_),
    .D(_04183_),
    .Y(_04185_));
 sky130_fd_sc_hd__a22o_1 _32361_ (.A1(_04175_),
    .A2(_04176_),
    .B1(_04181_),
    .B2(_04183_),
    .X(_04186_));
 sky130_fd_sc_hd__nand2_1 _32362_ (.A(_02366_),
    .B(_02374_),
    .Y(_04187_));
 sky130_fd_sc_hd__a21o_1 _32363_ (.A1(_04185_),
    .A2(_04186_),
    .B1(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__nand3_2 _32364_ (.A(_04187_),
    .B(_04185_),
    .C(_04186_),
    .Y(_04189_));
 sky130_fd_sc_hd__nand2_1 _32365_ (.A(_04188_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__and2_1 _32366_ (.A(_02376_),
    .B(_02378_),
    .X(_04191_));
 sky130_fd_sc_hd__or3b_2 _32367_ (.A(_17095_),
    .B(_18317_),
    .C_N(_06865_),
    .X(_04192_));
 sky130_fd_sc_hd__and4_1 _32368_ (.A(_04188_),
    .B(_02360_),
    .C(_04192_),
    .D(_04189_),
    .X(_04193_));
 sky130_fd_sc_hd__a22oi_1 _32369_ (.A1(_02360_),
    .A2(_04192_),
    .B1(_04188_),
    .B2(_04189_),
    .Y(_04194_));
 sky130_fd_sc_hd__o21ai_1 _32370_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04191_),
    .Y(_04196_));
 sky130_fd_sc_hd__o2111a_1 _32371_ (.A1(_04190_),
    .A2(_04191_),
    .B1(_24549_),
    .C1(_17095_),
    .D1(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__a211o_1 _32372_ (.A1(_02376_),
    .A2(_02378_),
    .B1(_04193_),
    .C1(_04194_),
    .X(_04198_));
 sky130_fd_sc_hd__o2bb2a_1 _32373_ (.A1_N(_04196_),
    .A2_N(_04198_),
    .B1(_02360_),
    .B2(_02361_),
    .X(_04199_));
 sky130_fd_sc_hd__o211ai_2 _32374_ (.A1(_04197_),
    .A2(_04199_),
    .B1(_02384_),
    .C1(_02385_),
    .Y(_04200_));
 sky130_fd_sc_hd__a211o_1 _32375_ (.A1(_02384_),
    .A2(_02385_),
    .B1(_04197_),
    .C1(_04199_),
    .X(_04201_));
 sky130_fd_sc_hd__o21bai_1 _32376_ (.A1(_02387_),
    .A2(_02389_),
    .B1_N(_02390_),
    .Y(_04202_));
 sky130_fd_sc_hd__a21oi_1 _32377_ (.A1(_04200_),
    .A2(_04201_),
    .B1(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__and3_1 _32378_ (.A(_04202_),
    .B(_04200_),
    .C(_04201_),
    .X(_04204_));
 sky130_fd_sc_hd__a31oi_2 _32379_ (.A1(_00584_),
    .A2(_00583_),
    .A3(_02356_),
    .B1(_02355_),
    .Y(_04205_));
 sky130_fd_sc_hd__nor2_1 _32380_ (.A(\delay_line[24][8] ),
    .B(\delay_line[24][9] ),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_1 _32381_ (.A(_22883_),
    .B(_24579_),
    .Y(_04208_));
 sky130_fd_sc_hd__nand3b_1 _32382_ (.A_N(_04207_),
    .B(_04208_),
    .C(_21620_),
    .Y(_04209_));
 sky130_fd_sc_hd__and2_1 _32383_ (.A(net342),
    .B(\delay_line[24][9] ),
    .X(_04210_));
 sky130_fd_sc_hd__inv_2 _32384_ (.A(_21619_),
    .Y(_04211_));
 sky130_fd_sc_hd__o21ai_1 _32385_ (.A1(_04207_),
    .A2(_04210_),
    .B1(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__clkbuf_2 _32386_ (.A(net341),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_2 _32387_ (.A(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__a21o_1 _32388_ (.A1(_04209_),
    .A2(_04212_),
    .B1(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__nand3_2 _32389_ (.A(_04212_),
    .B(_04214_),
    .C(_04209_),
    .Y(_04216_));
 sky130_fd_sc_hd__nand3_2 _32390_ (.A(_04215_),
    .B(_02320_),
    .C(_04216_),
    .Y(_04218_));
 sky130_fd_sc_hd__a21o_1 _32391_ (.A1(_04216_),
    .A2(_04215_),
    .B1(_02320_),
    .X(_04219_));
 sky130_fd_sc_hd__o21a_1 _32392_ (.A1(_20464_),
    .A2(_02314_),
    .B1(_02316_),
    .X(_04220_));
 sky130_fd_sc_hd__a21oi_1 _32393_ (.A1(_04218_),
    .A2(_04219_),
    .B1(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__and3_1 _32394_ (.A(_04219_),
    .B(_04220_),
    .C(_04218_),
    .X(_04222_));
 sky130_fd_sc_hd__a21boi_1 _32395_ (.A1(_02331_),
    .A2(_02313_),
    .B1_N(_02330_),
    .Y(_04223_));
 sky130_fd_sc_hd__o21ai_1 _32396_ (.A1(_04221_),
    .A2(_04222_),
    .B1(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__clkbuf_2 _32397_ (.A(_20464_),
    .X(_04225_));
 sky130_fd_sc_hd__o211a_1 _32398_ (.A1(_04225_),
    .A2(_21628_),
    .B1(_17029_),
    .C1(_19519_),
    .X(_04226_));
 sky130_fd_sc_hd__o21ba_1 _32399_ (.A1(_02336_),
    .A2(_00552_),
    .B1_N(_17029_),
    .X(_04227_));
 sky130_fd_sc_hd__nor2_1 _32400_ (.A(_04226_),
    .B(_04227_),
    .Y(_04229_));
 sky130_fd_sc_hd__a21o_1 _32401_ (.A1(_04218_),
    .A2(_04219_),
    .B1(_04220_),
    .X(_04230_));
 sky130_fd_sc_hd__o2111ai_1 _32402_ (.A1(_04225_),
    .A2(_02314_),
    .B1(_02316_),
    .C1(_04218_),
    .D1(_04219_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand3b_1 _32403_ (.A_N(_04223_),
    .B(_04230_),
    .C(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__nand3_1 _32404_ (.A(_04224_),
    .B(_04229_),
    .C(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__a2bb2o_1 _32405_ (.A1_N(_04226_),
    .A2_N(_04227_),
    .B1(_04232_),
    .B2(_04224_),
    .X(_04234_));
 sky130_fd_sc_hd__nand2_1 _32406_ (.A(_02342_),
    .B(_02343_),
    .Y(_04235_));
 sky130_fd_sc_hd__a21o_1 _32407_ (.A1(_04233_),
    .A2(_04234_),
    .B1(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__nand3_1 _32408_ (.A(_04235_),
    .B(_04233_),
    .C(_04234_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand3_1 _32409_ (.A(_04236_),
    .B(_04237_),
    .C(_02339_),
    .Y(_04238_));
 sky130_fd_sc_hd__a21o_1 _32410_ (.A1(_04236_),
    .A2(_04237_),
    .B1(_02339_),
    .X(_04240_));
 sky130_fd_sc_hd__nand2_1 _32411_ (.A(_04238_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__o311a_1 _32412_ (.A1(_19508_),
    .A2(_24572_),
    .A3(_02352_),
    .B1(_04241_),
    .C1(_02346_),
    .X(_04242_));
 sky130_fd_sc_hd__a21oi_1 _32413_ (.A1(_02346_),
    .A2(_02351_),
    .B1(_04241_),
    .Y(_04243_));
 sky130_fd_sc_hd__or2_1 _32414_ (.A(_04242_),
    .B(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__nor2_1 _32415_ (.A(_04205_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__o221a_1 _32416_ (.A1(_02354_),
    .A2(_02311_),
    .B1(_02357_),
    .B2(_00586_),
    .C1(_04244_),
    .X(_04246_));
 sky130_fd_sc_hd__or4_1 _32417_ (.A(_04203_),
    .B(_04204_),
    .C(_04245_),
    .D(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__inv_2 _32418_ (.A(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__o22a_1 _32419_ (.A1(_04203_),
    .A2(_04204_),
    .B1(_04245_),
    .B2(_04246_),
    .X(_04249_));
 sky130_fd_sc_hd__nor2_2 _32420_ (.A(_04248_),
    .B(_04249_),
    .Y(_04251_));
 sky130_fd_sc_hd__xnor2_4 _32421_ (.A(_04172_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__o311a_1 _32422_ (.A1(_02581_),
    .A2(_02582_),
    .A3(_02666_),
    .B1(_04252_),
    .C1(_02664_),
    .X(_04253_));
 sky130_fd_sc_hd__a21oi_4 _32423_ (.A1(_02664_),
    .A2(_02669_),
    .B1(_04252_),
    .Y(_04254_));
 sky130_fd_sc_hd__nor2_2 _32424_ (.A(_04253_),
    .B(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__and2b_1 _32425_ (.A_N(_04138_),
    .B(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__and2b_1 _32426_ (.A_N(_04255_),
    .B(_04138_),
    .X(_04257_));
 sky130_fd_sc_hd__or2_1 _32427_ (.A(_04256_),
    .B(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__xor2_1 _32428_ (.A(_04137_),
    .B(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__o32a_2 _32429_ (.A1(_02670_),
    .A2(_02671_),
    .A3(_02673_),
    .B1(_02674_),
    .B2(_02404_),
    .X(_04260_));
 sky130_fd_sc_hd__nand2_1 _32430_ (.A(_04259_),
    .B(_04260_),
    .Y(_04262_));
 sky130_fd_sc_hd__or2_1 _32431_ (.A(_04260_),
    .B(_04259_),
    .X(_04263_));
 sky130_fd_sc_hd__nand2_1 _32432_ (.A(_04262_),
    .B(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__or3b_1 _32433_ (.A(_02170_),
    .B(_02171_),
    .C_N(_02173_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_2 _32434_ (.A(net325),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_2 _32435_ (.A(_01032_),
    .X(_04267_));
 sky130_fd_sc_hd__or3b_1 _32436_ (.A(_01028_),
    .B(_04266_),
    .C_N(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__buf_1 _32437_ (.A(_23177_),
    .X(_04269_));
 sky130_fd_sc_hd__inv_2 _32438_ (.A(net325),
    .Y(_04270_));
 sky130_fd_sc_hd__or3b_1 _32439_ (.A(net326),
    .B(_04270_),
    .C_N(net324),
    .X(_04271_));
 sky130_fd_sc_hd__o21a_1 _32440_ (.A1(\delay_line[28][12] ),
    .A2(net324),
    .B1(_04271_),
    .X(_04273_));
 sky130_fd_sc_hd__or3b_2 _32441_ (.A(net324),
    .B(_04270_),
    .C_N(_01032_),
    .X(_04274_));
 sky130_fd_sc_hd__and3_1 _32442_ (.A(_04269_),
    .B(_04273_),
    .C(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__a21oi_1 _32443_ (.A1(_04273_),
    .A2(_04274_),
    .B1(_04269_),
    .Y(_04276_));
 sky130_fd_sc_hd__a211oi_1 _32444_ (.A1(_04265_),
    .A2(_04268_),
    .B1(_04275_),
    .C1(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__o211a_1 _32445_ (.A1(_04275_),
    .A2(_04276_),
    .B1(_04265_),
    .C1(_04268_),
    .X(_04278_));
 sky130_fd_sc_hd__o21bai_1 _32446_ (.A1(_04277_),
    .A2(_04278_),
    .B1_N(_02173_),
    .Y(_04279_));
 sky130_fd_sc_hd__or3b_1 _32447_ (.A(_04277_),
    .B(_04278_),
    .C_N(_02173_),
    .X(_04280_));
 sky130_fd_sc_hd__o211a_1 _32448_ (.A1(_02176_),
    .A2(net230),
    .B1(_04279_),
    .C1(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__a211oi_1 _32449_ (.A1(_04279_),
    .A2(_04280_),
    .B1(_02176_),
    .C1(net230),
    .Y(_04282_));
 sky130_fd_sc_hd__nor2_1 _32450_ (.A(_04281_),
    .B(_04282_),
    .Y(_04284_));
 sky130_fd_sc_hd__xor2_1 _32451_ (.A(_02182_),
    .B(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__a21oi_1 _32452_ (.A1(_02168_),
    .A2(_02186_),
    .B1(_02185_),
    .Y(_04286_));
 sky130_fd_sc_hd__nor2_1 _32453_ (.A(_04285_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__and2_1 _32454_ (.A(_04286_),
    .B(_04285_),
    .X(_04288_));
 sky130_fd_sc_hd__or2_1 _32455_ (.A(_04287_),
    .B(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__inv_2 _32456_ (.A(net336),
    .Y(_04290_));
 sky130_fd_sc_hd__nor2_1 _32457_ (.A(_02191_),
    .B(\delay_line[26][8] ),
    .Y(_04291_));
 sky130_fd_sc_hd__nand2_1 _32458_ (.A(_02191_),
    .B(_23140_),
    .Y(_04292_));
 sky130_fd_sc_hd__nand3b_1 _32459_ (.A_N(_04291_),
    .B(_04292_),
    .C(_19271_),
    .Y(_04293_));
 sky130_fd_sc_hd__and2_1 _32460_ (.A(_02191_),
    .B(\delay_line[26][8] ),
    .X(_04295_));
 sky130_fd_sc_hd__o21bai_1 _32461_ (.A1(_04291_),
    .A2(_04295_),
    .B1_N(_19271_),
    .Y(_04296_));
 sky130_fd_sc_hd__o21ai_1 _32462_ (.A1(_21223_),
    .A2(_02192_),
    .B1(_02193_),
    .Y(_04297_));
 sky130_fd_sc_hd__and3_1 _32463_ (.A(_04293_),
    .B(_04296_),
    .C(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__buf_1 _32464_ (.A(_04293_),
    .X(_04299_));
 sky130_fd_sc_hd__a21oi_1 _32465_ (.A1(_04299_),
    .A2(_04296_),
    .B1(_04297_),
    .Y(_04300_));
 sky130_fd_sc_hd__nor2_1 _32466_ (.A(_04298_),
    .B(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__o21bai_1 _32467_ (.A1(_02190_),
    .A2(_02200_),
    .B1_N(_02203_),
    .Y(_04302_));
 sky130_fd_sc_hd__xnor2_1 _32468_ (.A(_04301_),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__xor2_1 _32469_ (.A(_04290_),
    .B(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__a31oi_2 _32470_ (.A1(_24350_),
    .A2(_02188_),
    .A3(_02201_),
    .B1(_02208_),
    .Y(_04306_));
 sky130_fd_sc_hd__xnor2_1 _32471_ (.A(_04304_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21boi_1 _32472_ (.A1(_01014_),
    .A2(_01019_),
    .B1_N(_01015_),
    .Y(_04308_));
 sky130_fd_sc_hd__o21bai_1 _32473_ (.A1(_02211_),
    .A2(_04308_),
    .B1_N(_02210_),
    .Y(_04309_));
 sky130_fd_sc_hd__xnor2_1 _32474_ (.A(_04307_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32475_ (.A(_02237_),
    .X(_04311_));
 sky130_fd_sc_hd__o32a_1 _32476_ (.A1(net274),
    .A2(_19286_),
    .A3(_02229_),
    .B1(_02214_),
    .B2(_02223_),
    .X(_04312_));
 sky130_fd_sc_hd__nand2_1 _32477_ (.A(_20377_),
    .B(_23147_),
    .Y(_04313_));
 sky130_fd_sc_hd__inv_2 _32478_ (.A(net330),
    .Y(_04314_));
 sky130_fd_sc_hd__inv_2 _32479_ (.A(\delay_line[27][13] ),
    .Y(_04315_));
 sky130_fd_sc_hd__nand2_1 _32480_ (.A(_04314_),
    .B(_04315_),
    .Y(_04317_));
 sky130_fd_sc_hd__buf_1 _32481_ (.A(\delay_line[27][13] ),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _32482_ (.A(_00971_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__nand4_1 _32483_ (.A(_04317_),
    .B(_02223_),
    .C(_24366_),
    .D(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__a22o_1 _32484_ (.A1(_24366_),
    .A2(_02217_),
    .B1(_04319_),
    .B2(_04317_),
    .X(_04321_));
 sky130_fd_sc_hd__and4b_1 _32485_ (.A_N(_02215_),
    .B(_02218_),
    .C(_04318_),
    .D(_00968_),
    .X(_04322_));
 sky130_fd_sc_hd__a31o_1 _32486_ (.A1(_02219_),
    .A2(_04320_),
    .A3(_04321_),
    .B1(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__xnor2_2 _32487_ (.A(_04313_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__xor2_2 _32488_ (.A(_04312_),
    .B(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__xor2_2 _32489_ (.A(net274),
    .B(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__a21o_1 _32490_ (.A1(_02236_),
    .A2(_04311_),
    .B1(_04326_),
    .X(_04328_));
 sky130_fd_sc_hd__nand3_1 _32491_ (.A(_02236_),
    .B(_04311_),
    .C(_04326_),
    .Y(_04329_));
 sky130_fd_sc_hd__and2_1 _32492_ (.A(_04328_),
    .B(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__and4_1 _32493_ (.A(_04330_),
    .B(_02241_),
    .C(_02239_),
    .D(_04311_),
    .X(_04331_));
 sky130_fd_sc_hd__a31oi_1 _32494_ (.A1(_04311_),
    .A2(_02239_),
    .A3(_02241_),
    .B1(_04330_),
    .Y(_04332_));
 sky130_fd_sc_hd__nor2_1 _32495_ (.A(_04331_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__o21bai_1 _32496_ (.A1(_00989_),
    .A2(_00991_),
    .B1_N(_00988_),
    .Y(_04334_));
 sky130_fd_sc_hd__a211o_1 _32497_ (.A1(_24374_),
    .A2(_24375_),
    .B1(_00983_),
    .C1(_02242_),
    .X(_04335_));
 sky130_fd_sc_hd__a21boi_1 _32498_ (.A1(_04334_),
    .A2(_02244_),
    .B1_N(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__xnor2_1 _32499_ (.A(_04333_),
    .B(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__xor2_1 _32500_ (.A(_04310_),
    .B(_04337_),
    .X(_04339_));
 sky130_fd_sc_hd__xnor2_1 _32501_ (.A(_04289_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__o311a_1 _32502_ (.A1(_02212_),
    .A2(_02213_),
    .A3(_02247_),
    .B1(_02252_),
    .C1(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__a21oi_2 _32503_ (.A1(_02248_),
    .A2(_02252_),
    .B1(_04340_),
    .Y(_04342_));
 sky130_fd_sc_hd__nor2_2 _32504_ (.A(_04341_),
    .B(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__inv_2 _32505_ (.A(_02157_),
    .Y(_04344_));
 sky130_fd_sc_hd__a21bo_2 _32506_ (.A1(_02153_),
    .A2(_00901_),
    .B1_N(_02152_),
    .X(_04345_));
 sky130_fd_sc_hd__nor2_1 _32507_ (.A(_02143_),
    .B(_23212_),
    .Y(_04346_));
 sky130_fd_sc_hd__and2_1 _32508_ (.A(_23212_),
    .B(_20307_),
    .X(_04347_));
 sky130_fd_sc_hd__or3_2 _32509_ (.A(_02145_),
    .B(_04346_),
    .C(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__a2bb2o_1 _32510_ (.A1_N(_04346_),
    .A2_N(_04347_),
    .B1(_24447_),
    .B2(_02144_),
    .X(_04350_));
 sky130_fd_sc_hd__buf_1 _32511_ (.A(\delay_line[31][12] ),
    .X(_04351_));
 sky130_fd_sc_hd__nor2_1 _32512_ (.A(_04351_),
    .B(\delay_line[31][13] ),
    .Y(_04352_));
 sky130_fd_sc_hd__inv_2 _32513_ (.A(_00885_),
    .Y(_04353_));
 sky130_fd_sc_hd__and2_1 _32514_ (.A(_02127_),
    .B(\delay_line[31][13] ),
    .X(_04354_));
 sky130_fd_sc_hd__nor3_1 _32515_ (.A(_04352_),
    .B(_04353_),
    .C(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__o21a_1 _32516_ (.A1(_04354_),
    .A2(_04352_),
    .B1(_04353_),
    .X(_04356_));
 sky130_fd_sc_hd__a211o_1 _32517_ (.A1(_02130_),
    .A2(_02136_),
    .B1(_04355_),
    .C1(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__o211ai_2 _32518_ (.A1(_04355_),
    .A2(_04356_),
    .B1(_02130_),
    .C1(_02136_),
    .Y(_04358_));
 sky130_fd_sc_hd__nand3_2 _32519_ (.A(_04357_),
    .B(_04358_),
    .C(_02135_),
    .Y(_04359_));
 sky130_fd_sc_hd__a32o_1 _32520_ (.A1(_02136_),
    .A2(_02133_),
    .A3(_02134_),
    .B1(_04357_),
    .B2(_04358_),
    .X(_04361_));
 sky130_fd_sc_hd__nand4_2 _32521_ (.A(_04348_),
    .B(_04350_),
    .C(_04359_),
    .D(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__a22o_1 _32522_ (.A1(_04348_),
    .A2(_04350_),
    .B1(_04359_),
    .B2(_04361_),
    .X(_04363_));
 sky130_fd_sc_hd__nand2_1 _32523_ (.A(_02138_),
    .B(_02149_),
    .Y(_04364_));
 sky130_fd_sc_hd__and3_1 _32524_ (.A(_04362_),
    .B(_04363_),
    .C(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__a21oi_1 _32525_ (.A1(_04362_),
    .A2(_04363_),
    .B1(_04364_),
    .Y(_04366_));
 sky130_fd_sc_hd__nor2_1 _32526_ (.A(_04365_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__and4b_1 _32527_ (.A_N(_00900_),
    .B(_04367_),
    .C(_02142_),
    .D(_02145_),
    .X(_04368_));
 sky130_fd_sc_hd__o21a_1 _32528_ (.A1(_04365_),
    .A2(_04366_),
    .B1(_02146_),
    .X(_04369_));
 sky130_fd_sc_hd__nor2_2 _32529_ (.A(_04368_),
    .B(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hd__xor2_4 _32530_ (.A(_04345_),
    .B(_04370_),
    .X(_04372_));
 sky130_fd_sc_hd__nor2_1 _32531_ (.A(_02126_),
    .B(_02158_),
    .Y(_04373_));
 sky130_fd_sc_hd__o21bai_4 _32532_ (.A1(_02159_),
    .A2(_02163_),
    .B1_N(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__xor2_2 _32533_ (.A(_04372_),
    .B(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__o21bai_2 _32534_ (.A1(_02159_),
    .A2(_02163_),
    .B1_N(_04372_),
    .Y(_04376_));
 sky130_fd_sc_hd__nand2_2 _32535_ (.A(_04376_),
    .B(_04344_),
    .Y(_04377_));
 sky130_fd_sc_hd__buf_2 _32536_ (.A(\delay_line[30][10] ),
    .X(_04378_));
 sky130_fd_sc_hd__xor2_1 _32537_ (.A(_23269_),
    .B(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__or2_1 _32538_ (.A(\delay_line[30][13] ),
    .B(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__nor2_1 _32539_ (.A(_02103_),
    .B(_02107_),
    .Y(_04381_));
 sky130_fd_sc_hd__clkbuf_2 _32540_ (.A(\delay_line[30][12] ),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_2 _32541_ (.A(_04379_),
    .X(_04384_));
 sky130_fd_sc_hd__nand2_1 _32542_ (.A(\delay_line[30][13] ),
    .B(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__and4_1 _32543_ (.A(_04380_),
    .B(_04381_),
    .C(_04383_),
    .D(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__a22oi_2 _32544_ (.A1(_04383_),
    .A2(_04381_),
    .B1(_04385_),
    .B2(_04380_),
    .Y(_04387_));
 sky130_fd_sc_hd__and3_1 _32545_ (.A(_18453_),
    .B(_00940_),
    .C(_02102_),
    .X(_04388_));
 sky130_fd_sc_hd__a21oi_1 _32546_ (.A1(_24394_),
    .A2(_24395_),
    .B1(_02107_),
    .Y(_04389_));
 sky130_fd_sc_hd__o22a_1 _32547_ (.A1(_20350_),
    .A2(_15580_),
    .B1(_04388_),
    .B2(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__a2111oi_1 _32548_ (.A1(_18453_),
    .A2(_02107_),
    .B1(_20350_),
    .C1(_15580_),
    .D1(_04389_),
    .Y(_04391_));
 sky130_fd_sc_hd__nor4_1 _32549_ (.A(_04386_),
    .B(_04387_),
    .C(_04390_),
    .D(net253),
    .Y(_04392_));
 sky130_fd_sc_hd__o22a_1 _32550_ (.A1(_04386_),
    .A2(_04387_),
    .B1(_04390_),
    .B2(net253),
    .X(_04394_));
 sky130_fd_sc_hd__a211oi_2 _32551_ (.A1(_02111_),
    .A2(_02112_),
    .B1(net202),
    .C1(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__o211a_1 _32552_ (.A1(net203),
    .A2(_04394_),
    .B1(_02111_),
    .C1(_02112_),
    .X(_04396_));
 sky130_fd_sc_hd__nor2_1 _32553_ (.A(_04395_),
    .B(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__o21a_2 _32554_ (.A1(_02096_),
    .A2(_02094_),
    .B1(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_2 _32555_ (.A(_23269_),
    .X(_04399_));
 sky130_fd_sc_hd__a311oi_2 _32556_ (.A1(_15580_),
    .A2(_19336_),
    .A3(_04399_),
    .B1(_02094_),
    .C1(_04397_),
    .Y(_04400_));
 sky130_fd_sc_hd__o21ba_1 _32557_ (.A1(_02091_),
    .A2(_02115_),
    .B1_N(_02116_),
    .X(_04401_));
 sky130_fd_sc_hd__o21a_1 _32558_ (.A1(_04398_),
    .A2(_04400_),
    .B1(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__nor3_2 _32559_ (.A(_04401_),
    .B(_04398_),
    .C(_04400_),
    .Y(_04403_));
 sky130_fd_sc_hd__o2bb2ai_1 _32560_ (.A1_N(_02121_),
    .A2_N(_02123_),
    .B1(_04402_),
    .B2(_04403_),
    .Y(_04405_));
 sky130_fd_sc_hd__and2_1 _32561_ (.A(_02088_),
    .B(_02119_),
    .X(_04406_));
 sky130_fd_sc_hd__buf_1 _32562_ (.A(_02076_),
    .X(_04407_));
 sky130_fd_sc_hd__and2b_1 _32563_ (.A_N(_00915_),
    .B(\delay_line[29][11] ),
    .X(_04408_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32564_ (.A(\delay_line[29][11] ),
    .X(_04409_));
 sky130_fd_sc_hd__or2b_1 _32565_ (.A(_04409_),
    .B_N(_00915_),
    .X(_04410_));
 sky130_fd_sc_hd__and2b_1 _32566_ (.A_N(_04408_),
    .B(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__a21oi_1 _32567_ (.A1(_00917_),
    .A2(_02078_),
    .B1(_04407_),
    .Y(_04412_));
 sky130_fd_sc_hd__xor2_1 _32568_ (.A(_04411_),
    .B(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__o311a_1 _32569_ (.A1(_04407_),
    .A2(_02077_),
    .A3(_02075_),
    .B1(_04413_),
    .C1(_02083_),
    .X(_04414_));
 sky130_fd_sc_hd__or2_1 _32570_ (.A(_04402_),
    .B(_04403_),
    .X(_04416_));
 sky130_fd_sc_hd__a32oi_4 _32571_ (.A1(_00927_),
    .A2(_00953_),
    .A3(_02120_),
    .B1(_02123_),
    .B2(_02121_),
    .Y(_04417_));
 sky130_fd_sc_hd__xor2_1 _32572_ (.A(_04416_),
    .B(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__a21oi_2 _32573_ (.A1(_02088_),
    .A2(_02119_),
    .B1(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__or3_1 _32574_ (.A(_04407_),
    .B(_02077_),
    .C(_02075_),
    .X(_04420_));
 sky130_fd_sc_hd__a21oi_2 _32575_ (.A1(_02083_),
    .A2(_04420_),
    .B1(_04413_),
    .Y(_04421_));
 sky130_fd_sc_hd__a2111oi_1 _32576_ (.A1(_04405_),
    .A2(_04406_),
    .B1(_04414_),
    .C1(_04419_),
    .D1(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__inv_2 _32577_ (.A(net90),
    .Y(_04423_));
 sky130_fd_sc_hd__and3_1 _32578_ (.A(_02088_),
    .B(_02119_),
    .C(_04405_),
    .X(_04424_));
 sky130_fd_sc_hd__o22ai_4 _32579_ (.A1(_04414_),
    .A2(_04421_),
    .B1(_04424_),
    .B2(_04419_),
    .Y(_04425_));
 sky130_fd_sc_hd__o2111ai_4 _32580_ (.A1(_04344_),
    .A2(_04375_),
    .B1(_04377_),
    .C1(_04423_),
    .D1(_04425_),
    .Y(_04427_));
 sky130_fd_sc_hd__o21a_1 _32581_ (.A1(_04344_),
    .A2(_04375_),
    .B1(_04377_),
    .X(_04428_));
 sky130_fd_sc_hd__a21o_1 _32582_ (.A1(_04423_),
    .A2(_04425_),
    .B1(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__and2_2 _32583_ (.A(_04427_),
    .B(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__xnor2_4 _32584_ (.A(_04343_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__a21oi_1 _32585_ (.A1(_02399_),
    .A2(_02400_),
    .B1(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__o211ai_1 _32586_ (.A1(_02401_),
    .A2(_02267_),
    .B1(_02399_),
    .C1(_04431_),
    .Y(_04433_));
 sky130_fd_sc_hd__or2b_1 _32587_ (.A(_04432_),
    .B_N(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__a21o_2 _32588_ (.A1(_02167_),
    .A2(_02257_),
    .B1(_02256_),
    .X(_04435_));
 sky130_fd_sc_hd__xor2_1 _32589_ (.A(_04434_),
    .B(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__nand2_1 _32590_ (.A(_04264_),
    .B(_04436_),
    .Y(_04438_));
 sky130_fd_sc_hd__or2_1 _32591_ (.A(_04264_),
    .B(_04436_),
    .X(_04439_));
 sky130_fd_sc_hd__nand2_1 _32592_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__xnor2_2 _32593_ (.A(_03871_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__o21ai_1 _32594_ (.A1(_03868_),
    .A2(_03869_),
    .B1(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__o31ai_1 _32595_ (.A1(_03868_),
    .A2(_03869_),
    .A3(_04441_),
    .B1(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__nor2_1 _32596_ (.A(_03619_),
    .B(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__and2_1 _32597_ (.A(_03619_),
    .B(_04443_),
    .X(_04445_));
 sky130_fd_sc_hd__or2_1 _32598_ (.A(_04444_),
    .B(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__o21bai_1 _32599_ (.A1(_03617_),
    .A2(_03618_),
    .B1_N(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__a21o_1 _32600_ (.A1(_03608_),
    .A2(_03614_),
    .B1(_03616_),
    .X(_04449_));
 sky130_fd_sc_hd__o211ai_2 _32601_ (.A1(_02037_),
    .A2(_03615_),
    .B1(_03607_),
    .C1(_03614_),
    .Y(_04450_));
 sky130_fd_sc_hd__clkbuf_2 _32602_ (.A(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__o211ai_1 _32603_ (.A1(_04444_),
    .A2(_04445_),
    .B1(_04449_),
    .C1(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__or2b_1 _32604_ (.A(_02925_),
    .B_N(_02070_),
    .X(_04453_));
 sky130_fd_sc_hd__o21ai_1 _32605_ (.A1(_02066_),
    .A2(_02927_),
    .B1(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__a21oi_1 _32606_ (.A1(_04447_),
    .A2(_04452_),
    .B1(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__o21ai_1 _32607_ (.A1(_04444_),
    .A2(_04445_),
    .B1(_04450_),
    .Y(_04456_));
 sky130_fd_sc_hd__o211a_1 _32608_ (.A1(_03617_),
    .A2(_04456_),
    .B1(_04447_),
    .C1(_04454_),
    .X(_04457_));
 sky130_fd_sc_hd__o22ai_4 _32609_ (.A1(_03064_),
    .A2(_03065_),
    .B1(_04455_),
    .B2(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__a21oi_1 _32610_ (.A1(_04449_),
    .A2(_04451_),
    .B1(_04446_),
    .Y(_04460_));
 sky130_fd_sc_hd__a32o_1 _32611_ (.A1(_04449_),
    .A2(_04451_),
    .A3(_04446_),
    .B1(_02935_),
    .B2(_04453_),
    .X(_04461_));
 sky130_fd_sc_hd__nor2_1 _32612_ (.A(_03064_),
    .B(_03065_),
    .Y(_04462_));
 sky130_fd_sc_hd__a21o_1 _32613_ (.A1(_04447_),
    .A2(_04452_),
    .B1(_04454_),
    .X(_04463_));
 sky130_fd_sc_hd__o211ai_2 _32614_ (.A1(_04460_),
    .A2(_04461_),
    .B1(_04462_),
    .C1(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand3_1 _32615_ (.A(_02993_),
    .B(_04458_),
    .C(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__a21o_1 _32616_ (.A1(_04458_),
    .A2(_04464_),
    .B1(_02993_),
    .X(_04466_));
 sky130_fd_sc_hd__o21ai_2 _32617_ (.A1(_01414_),
    .A2(_01437_),
    .B1(_01440_),
    .Y(_04467_));
 sky130_fd_sc_hd__and2_1 _32618_ (.A(_11328_),
    .B(_23602_),
    .X(_04468_));
 sky130_fd_sc_hd__nor2_1 _32619_ (.A(_23602_),
    .B(_11328_),
    .Y(_04469_));
 sky130_fd_sc_hd__a211o_1 _32620_ (.A1(_10833_),
    .A2(_02952_),
    .B1(_04468_),
    .C1(_04469_),
    .X(_04471_));
 sky130_fd_sc_hd__o211ai_4 _32621_ (.A1(_04468_),
    .A2(_04469_),
    .B1(_10833_),
    .C1(_02952_),
    .Y(_04472_));
 sky130_fd_sc_hd__clkbuf_2 _32622_ (.A(_01409_),
    .X(_04473_));
 sky130_fd_sc_hd__and3b_2 _32623_ (.A_N(_04473_),
    .B(_25255_),
    .C(_25236_),
    .X(_04474_));
 sky130_fd_sc_hd__a221oi_2 _32624_ (.A1(_04471_),
    .A2(_04472_),
    .B1(_01408_),
    .B2(_23724_),
    .C1(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__and3_1 _32625_ (.A(_01408_),
    .B(_25236_),
    .C(_25242_),
    .X(_04476_));
 sky130_fd_sc_hd__buf_2 _32626_ (.A(_04471_),
    .X(_04477_));
 sky130_fd_sc_hd__o211ai_4 _32627_ (.A1(_04474_),
    .A2(_04476_),
    .B1(_04472_),
    .C1(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__and3b_1 _32628_ (.A_N(_04475_),
    .B(_02954_),
    .C(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__o211a_1 _32629_ (.A1(_04474_),
    .A2(_04476_),
    .B1(_04472_),
    .C1(_04477_),
    .X(_04480_));
 sky130_fd_sc_hd__o21ba_1 _32630_ (.A1(_04480_),
    .A2(_04475_),
    .B1_N(_02954_),
    .X(_04482_));
 sky130_fd_sc_hd__nor2_1 _32631_ (.A(_04479_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__xnor2_1 _32632_ (.A(_04467_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__and3_1 _32633_ (.A(_02958_),
    .B(_02959_),
    .C(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__a21oi_2 _32634_ (.A1(_02958_),
    .A2(_02959_),
    .B1(_04484_),
    .Y(_04486_));
 sky130_fd_sc_hd__or2_2 _32635_ (.A(_04485_),
    .B(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__and3_1 _32636_ (.A(_02965_),
    .B(_02967_),
    .C(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__a21oi_2 _32637_ (.A1(_02965_),
    .A2(_02967_),
    .B1(_04487_),
    .Y(_04489_));
 sky130_fd_sc_hd__or2_1 _32638_ (.A(_04488_),
    .B(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__a21oi_1 _32639_ (.A1(_01472_),
    .A2(_01470_),
    .B1(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__nand3_1 _32640_ (.A(_01472_),
    .B(_01470_),
    .C(_04490_),
    .Y(_04493_));
 sky130_fd_sc_hd__or2b_1 _32641_ (.A(_04491_),
    .B_N(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__xor2_1 _32642_ (.A(_02970_),
    .B(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__a21bo_1 _32643_ (.A1(_04465_),
    .A2(_04466_),
    .B1_N(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__o21a_1 _32644_ (.A1(_02939_),
    .A2(_02940_),
    .B1(_02932_),
    .X(_04497_));
 sky130_fd_sc_hd__nand2_1 _32645_ (.A(_04458_),
    .B(_04464_),
    .Y(_04498_));
 sky130_fd_sc_hd__a21oi_1 _32646_ (.A1(_04497_),
    .A2(_04498_),
    .B1(_04495_),
    .Y(_04499_));
 sky130_fd_sc_hd__o21ai_1 _32647_ (.A1(_04497_),
    .A2(_04498_),
    .B1(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__and3_1 _32648_ (.A(_01404_),
    .B(_02937_),
    .C(_02941_),
    .X(_04501_));
 sky130_fd_sc_hd__o21ai_1 _32649_ (.A1(_02976_),
    .A2(_04501_),
    .B1(_02947_),
    .Y(_04502_));
 sky130_fd_sc_hd__a21boi_2 _32650_ (.A1(_04496_),
    .A2(_04500_),
    .B1_N(_04502_),
    .Y(_04504_));
 sky130_fd_sc_hd__a21boi_1 _32651_ (.A1(_04465_),
    .A2(_04466_),
    .B1_N(_04495_),
    .Y(_04505_));
 sky130_fd_sc_hd__a211oi_1 _32652_ (.A1(_04465_),
    .A2(_04499_),
    .B1(_04502_),
    .C1(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__a21oi_1 _32653_ (.A1(_01373_),
    .A2(_02973_),
    .B1(_02972_),
    .Y(_04507_));
 sky130_fd_sc_hd__o21a_1 _32654_ (.A1(_04504_),
    .A2(_04506_),
    .B1(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__o211a_1 _32655_ (.A1(_25169_),
    .A2(_25173_),
    .B1(_01372_),
    .C1(_02973_),
    .X(_04509_));
 sky130_fd_sc_hd__o2111ai_1 _32656_ (.A1(_02976_),
    .A2(_04501_),
    .B1(_02947_),
    .C1(_04496_),
    .D1(_04500_),
    .Y(_04510_));
 sky130_fd_sc_hd__o21ai_1 _32657_ (.A1(_02972_),
    .A2(_04509_),
    .B1(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__nor2_1 _32658_ (.A(_04504_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__a31o_1 _32659_ (.A1(_02977_),
    .A2(_02978_),
    .A3(_02980_),
    .B1(_02988_),
    .X(_04513_));
 sky130_fd_sc_hd__nand2_1 _32660_ (.A(_02982_),
    .B(_04513_),
    .Y(_04515_));
 sky130_fd_sc_hd__o21bai_1 _32661_ (.A1(_04508_),
    .A2(_04512_),
    .B1_N(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__o21ai_1 _32662_ (.A1(_04504_),
    .A2(_04506_),
    .B1(_04507_),
    .Y(_04517_));
 sky130_fd_sc_hd__o211ai_2 _32663_ (.A1(_04504_),
    .A2(_04511_),
    .B1(_04517_),
    .C1(_04515_),
    .Y(_04518_));
 sky130_fd_sc_hd__nand2_2 _32664_ (.A(_04516_),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__nand3_1 _32665_ (.A(_02983_),
    .B(_02984_),
    .C(_02985_),
    .Y(_04520_));
 sky130_fd_sc_hd__a22oi_4 _32666_ (.A1(_02990_),
    .A2(_02989_),
    .B1(_02992_),
    .B2(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__xor2_4 _32667_ (.A(_04519_),
    .B(_04521_),
    .X(_00007_));
 sky130_fd_sc_hd__a2bb2o_1 _32668_ (.A1_N(_04460_),
    .A2_N(_04461_),
    .B1(_04462_),
    .B2(_04463_),
    .X(_04522_));
 sky130_fd_sc_hd__nor4_1 _32669_ (.A(_22781_),
    .B(_02038_),
    .C(_03038_),
    .D(_03039_),
    .Y(_04523_));
 sky130_fd_sc_hd__clkbuf_2 _32670_ (.A(net363),
    .X(_04525_));
 sky130_fd_sc_hd__clkbuf_2 _32671_ (.A(net364),
    .X(_04526_));
 sky130_fd_sc_hd__and3b_2 _32672_ (.A_N(_04525_),
    .B(_04526_),
    .C(_03030_),
    .X(_04527_));
 sky130_fd_sc_hd__and2_1 _32673_ (.A(net364),
    .B(net363),
    .X(_04528_));
 sky130_fd_sc_hd__nor2_1 _32674_ (.A(net364),
    .B(\delay_line[20][14] ),
    .Y(_04529_));
 sky130_fd_sc_hd__o2bb2a_1 _32675_ (.A1_N(_03030_),
    .A2_N(_04526_),
    .B1(_04528_),
    .B2(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__xnor2_1 _32676_ (.A(_23682_),
    .B(_01448_),
    .Y(_04531_));
 sky130_fd_sc_hd__nor3_2 _32677_ (.A(_04527_),
    .B(_04530_),
    .C(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__clkbuf_2 _32678_ (.A(_04531_),
    .X(_04533_));
 sky130_fd_sc_hd__o21a_1 _32679_ (.A1(_04527_),
    .A2(_04530_),
    .B1(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__or4_1 _32680_ (.A(_19848_),
    .B(_15163_),
    .C(_04532_),
    .D(_04534_),
    .X(_04536_));
 sky130_fd_sc_hd__o21ai_1 _32681_ (.A1(_04532_),
    .A2(_04534_),
    .B1(_03595_),
    .Y(_04537_));
 sky130_fd_sc_hd__o211a_1 _32682_ (.A1(_03036_),
    .A2(_03038_),
    .B1(_04536_),
    .C1(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__a221oi_2 _32683_ (.A1(_01447_),
    .A2(_03035_),
    .B1(_04536_),
    .B2(_04537_),
    .C1(_03038_),
    .Y(_04539_));
 sky130_fd_sc_hd__o221a_1 _32684_ (.A1(_03594_),
    .A2(_03596_),
    .B1(_04538_),
    .B2(_04539_),
    .C1(_03592_),
    .X(_04540_));
 sky130_fd_sc_hd__o21a_1 _32685_ (.A1(_03594_),
    .A2(_03596_),
    .B1(_03592_),
    .X(_04541_));
 sky130_fd_sc_hd__nor3_1 _32686_ (.A(_04541_),
    .B(_04538_),
    .C(_04539_),
    .Y(_04542_));
 sky130_fd_sc_hd__or2_1 _32687_ (.A(_04540_),
    .B(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__or3b_1 _32688_ (.A(net228),
    .B(_03043_),
    .C_N(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__o21bai_2 _32689_ (.A1(net227),
    .A2(_03043_),
    .B1_N(_04543_),
    .Y(_04545_));
 sky130_fd_sc_hd__a211oi_2 _32690_ (.A1(_04544_),
    .A2(_04545_),
    .B1(_03048_),
    .C1(_03053_),
    .Y(_04547_));
 sky130_fd_sc_hd__o211a_1 _32691_ (.A1(_03048_),
    .A2(_03053_),
    .B1(_04544_),
    .C1(_04545_),
    .X(_04548_));
 sky130_fd_sc_hd__nor2_1 _32692_ (.A(_25264_),
    .B(_01429_),
    .Y(_04549_));
 sky130_fd_sc_hd__and2_1 _32693_ (.A(_01429_),
    .B(_25264_),
    .X(_04550_));
 sky130_fd_sc_hd__nor2_1 _32694_ (.A(_03001_),
    .B(\delay_line[17][14] ),
    .Y(_04551_));
 sky130_fd_sc_hd__and2_1 _32695_ (.A(\delay_line[17][13] ),
    .B(\delay_line[17][14] ),
    .X(_04552_));
 sky130_fd_sc_hd__nor2_1 _32696_ (.A(_04551_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__o21ai_1 _32697_ (.A1(_04549_),
    .A2(_04550_),
    .B1(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__or3_1 _32698_ (.A(_04553_),
    .B(_04549_),
    .C(_04550_),
    .X(_04555_));
 sky130_fd_sc_hd__and2_1 _32699_ (.A(_04554_),
    .B(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__buf_1 _32700_ (.A(_25260_),
    .X(_04558_));
 sky130_fd_sc_hd__a21oi_1 _32701_ (.A1(_23681_),
    .A2(_25220_),
    .B1(_25219_),
    .Y(_04559_));
 sky130_fd_sc_hd__nor2_1 _32702_ (.A(_04559_),
    .B(_25223_),
    .Y(_04560_));
 sky130_fd_sc_hd__and2_1 _32703_ (.A(_25223_),
    .B(_04559_),
    .X(_04561_));
 sky130_fd_sc_hd__or3_1 _32704_ (.A(_04558_),
    .B(_04560_),
    .C(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__o21ai_1 _32705_ (.A1(_04560_),
    .A2(_04561_),
    .B1(_04558_),
    .Y(_04563_));
 sky130_fd_sc_hd__a211oi_1 _32706_ (.A1(_04562_),
    .A2(_04563_),
    .B1(_03013_),
    .C1(_03015_),
    .Y(_04564_));
 sky130_fd_sc_hd__o211ai_1 _32707_ (.A1(_03013_),
    .A2(_03015_),
    .B1(_04562_),
    .C1(_04563_),
    .Y(_04565_));
 sky130_fd_sc_hd__and2b_1 _32708_ (.A_N(_04564_),
    .B(_04565_),
    .X(_04566_));
 sky130_fd_sc_hd__xor2_1 _32709_ (.A(_04556_),
    .B(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__o211a_1 _32710_ (.A1(_03010_),
    .A2(_03019_),
    .B1(_03020_),
    .C1(_04567_),
    .X(_04569_));
 sky130_fd_sc_hd__o32a_1 _32711_ (.A1(_03017_),
    .A2(_03015_),
    .A3(_03016_),
    .B1(_03019_),
    .B2(_03010_),
    .X(_04570_));
 sky130_fd_sc_hd__nor2_2 _32712_ (.A(_04570_),
    .B(_04567_),
    .Y(_04571_));
 sky130_fd_sc_hd__clkbuf_2 _32713_ (.A(_04473_),
    .X(_04572_));
 sky130_fd_sc_hd__buf_1 _32714_ (.A(_02995_),
    .X(_04573_));
 sky130_fd_sc_hd__buf_1 _32715_ (.A(_03001_),
    .X(_04574_));
 sky130_fd_sc_hd__buf_1 _32716_ (.A(_02995_),
    .X(_04575_));
 sky130_fd_sc_hd__and2b_1 _32717_ (.A_N(_04574_),
    .B(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__a21oi_1 _32718_ (.A1(_19800_),
    .A2(_19815_),
    .B1(_03005_),
    .Y(_04577_));
 sky130_fd_sc_hd__or3b_1 _32719_ (.A(_04574_),
    .B(_03008_),
    .C_N(_04575_),
    .X(_04578_));
 sky130_fd_sc_hd__o31a_1 _32720_ (.A1(_03006_),
    .A2(_04576_),
    .A3(_04577_),
    .B1(_04578_),
    .X(_04580_));
 sky130_fd_sc_hd__a21oi_1 _32721_ (.A1(_04572_),
    .A2(_04573_),
    .B1(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32722_ (.A(_01416_),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_1 _32723_ (.A(_04582_),
    .B(_04580_),
    .Y(_04583_));
 sky130_fd_sc_hd__or2b_1 _32724_ (.A(_04581_),
    .B_N(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__o21a_1 _32725_ (.A1(_04569_),
    .A2(_04571_),
    .B1(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__nor3_2 _32726_ (.A(_04571_),
    .B(_04584_),
    .C(_04569_),
    .Y(_04586_));
 sky130_fd_sc_hd__or2_2 _32727_ (.A(_04585_),
    .B(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__or3_1 _32728_ (.A(_04547_),
    .B(_04548_),
    .C(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__o21ai_1 _32729_ (.A1(_04547_),
    .A2(_04548_),
    .B1(_04587_),
    .Y(_04589_));
 sky130_fd_sc_hd__nand2_1 _32730_ (.A(_04588_),
    .B(_04589_),
    .Y(_04591_));
 sky130_fd_sc_hd__a21oi_2 _32731_ (.A1(_03608_),
    .A2(_04451_),
    .B1(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__and3_1 _32732_ (.A(_03608_),
    .B(_04450_),
    .C(_04591_),
    .X(_04593_));
 sky130_fd_sc_hd__o21ai_2 _32733_ (.A1(_03055_),
    .A2(_03028_),
    .B1(_03056_),
    .Y(_04594_));
 sky130_fd_sc_hd__o21a_1 _32734_ (.A1(_04592_),
    .A2(_04593_),
    .B1(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__nor3_2 _32735_ (.A(_04594_),
    .B(_04592_),
    .C(_04593_),
    .Y(_04596_));
 sky130_fd_sc_hd__inv_2 _32736_ (.A(_03599_),
    .Y(_04597_));
 sky130_fd_sc_hd__inv_2 _32737_ (.A(_03569_),
    .Y(_04598_));
 sky130_fd_sc_hd__and2b_1 _32738_ (.A_N(_03679_),
    .B(_03655_),
    .X(_04599_));
 sky130_fd_sc_hd__nor2_2 _32739_ (.A(_03654_),
    .B(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__o211a_1 _32740_ (.A1(_01982_),
    .A2(_01983_),
    .B1(_01987_),
    .C1(_01984_),
    .X(_04602_));
 sky130_fd_sc_hd__nand2_1 _32741_ (.A(_01979_),
    .B(_03069_),
    .Y(_04603_));
 sky130_fd_sc_hd__o21a_1 _32742_ (.A1(_04602_),
    .A2(_04603_),
    .B1(_01989_),
    .X(_04604_));
 sky130_fd_sc_hd__a2bb2oi_1 _32743_ (.A1_N(_00402_),
    .A2_N(_00404_),
    .B1(_00408_),
    .B2(_24224_),
    .Y(_04605_));
 sky130_fd_sc_hd__o22ai_1 _32744_ (.A1(_03069_),
    .A2(_03070_),
    .B1(_03532_),
    .B2(_03536_),
    .Y(_04606_));
 sky130_fd_sc_hd__a21oi_1 _32745_ (.A1(_04604_),
    .A2(_04605_),
    .B1(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__inv_2 _32746_ (.A(_03393_),
    .Y(_04608_));
 sky130_fd_sc_hd__o21ai_1 _32747_ (.A1(_01799_),
    .A2(net231),
    .B1(_03328_),
    .Y(_04609_));
 sky130_fd_sc_hd__nand2_1 _32748_ (.A(_03321_),
    .B(_03325_),
    .Y(_04610_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32749_ (.A(_21821_),
    .X(_04611_));
 sky130_fd_sc_hd__a41oi_1 _32750_ (.A1(_22448_),
    .A2(_04611_),
    .A3(_03259_),
    .A4(_03261_),
    .B1(_03264_),
    .Y(_04613_));
 sky130_fd_sc_hd__clkbuf_2 _32751_ (.A(\delay_line[9][13] ),
    .X(_04614_));
 sky130_fd_sc_hd__o21a_1 _32752_ (.A1(_03311_),
    .A2(_01682_),
    .B1(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__nor3_1 _32753_ (.A(_03311_),
    .B(_04614_),
    .C(_03265_),
    .Y(_04616_));
 sky130_fd_sc_hd__o21a_1 _32754_ (.A1(_04615_),
    .A2(_04616_),
    .B1(_22440_),
    .X(_04617_));
 sky130_fd_sc_hd__nor3_1 _32755_ (.A(_22440_),
    .B(_04615_),
    .C(_04616_),
    .Y(_04618_));
 sky130_fd_sc_hd__or3_1 _32756_ (.A(_04613_),
    .B(_04617_),
    .C(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__o21ai_1 _32757_ (.A1(_04617_),
    .A2(_04618_),
    .B1(_04613_),
    .Y(_04620_));
 sky130_fd_sc_hd__nand2_1 _32758_ (.A(_03317_),
    .B(_03319_),
    .Y(_04621_));
 sky130_fd_sc_hd__a21oi_1 _32759_ (.A1(_04619_),
    .A2(_04620_),
    .B1(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__and3_1 _32760_ (.A(_04621_),
    .B(_04619_),
    .C(_04620_),
    .X(_04624_));
 sky130_fd_sc_hd__and2b_1 _32761_ (.A_N(_03272_),
    .B(_03274_),
    .X(_04625_));
 sky130_fd_sc_hd__o21ai_1 _32762_ (.A1(_04622_),
    .A2(_04624_),
    .B1(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__or3_2 _32763_ (.A(_04625_),
    .B(_04622_),
    .C(_04624_),
    .X(_04627_));
 sky130_fd_sc_hd__nand3_1 _32764_ (.A(_04610_),
    .B(_04626_),
    .C(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__a21o_1 _32765_ (.A1(_04626_),
    .A2(_04627_),
    .B1(_04610_),
    .X(_04629_));
 sky130_fd_sc_hd__nand2_1 _32766_ (.A(_04628_),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__a21oi_1 _32767_ (.A1(_03327_),
    .A2(_04609_),
    .B1(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__and3_1 _32768_ (.A(_03327_),
    .B(_04609_),
    .C(_04630_),
    .X(_04632_));
 sky130_fd_sc_hd__a21bo_1 _32769_ (.A1(_03360_),
    .A2(_01771_),
    .B1_N(_03352_),
    .X(_04633_));
 sky130_fd_sc_hd__nand2b_1 _32770_ (.A_N(\delay_line[8][12] ),
    .B(\delay_line[8][13] ),
    .Y(_04635_));
 sky130_fd_sc_hd__nand2b_1 _32771_ (.A_N(\delay_line[8][13] ),
    .B(\delay_line[8][12] ),
    .Y(_04636_));
 sky130_fd_sc_hd__nand2_1 _32772_ (.A(_04635_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__nand2_1 _32773_ (.A(_04637_),
    .B(_03360_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand3b_1 _32774_ (.A_N(_03360_),
    .B(_04635_),
    .C(_04636_),
    .Y(_04639_));
 sky130_fd_sc_hd__nand3_2 _32775_ (.A(_04633_),
    .B(_04638_),
    .C(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__a21o_1 _32776_ (.A1(_04638_),
    .A2(_04639_),
    .B1(_04633_),
    .X(_04641_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32777_ (.A(_01739_),
    .X(_04642_));
 sky130_fd_sc_hd__a21o_1 _32778_ (.A1(_04640_),
    .A2(_04641_),
    .B1(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__nand3_2 _32779_ (.A(_04641_),
    .B(_04642_),
    .C(_04640_),
    .Y(_04644_));
 sky130_fd_sc_hd__clkbuf_2 _32780_ (.A(_03369_),
    .X(_04646_));
 sky130_fd_sc_hd__or2b_1 _32781_ (.A(_17916_),
    .B_N(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__nand3b_1 _32782_ (.A_N(_18052_),
    .B(_03347_),
    .C(_03371_),
    .Y(_04648_));
 sky130_fd_sc_hd__clkbuf_2 _32783_ (.A(net423),
    .X(_04649_));
 sky130_fd_sc_hd__xnor2_2 _32784_ (.A(_20122_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__and3_1 _32785_ (.A(_04647_),
    .B(_04648_),
    .C(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__a21oi_1 _32786_ (.A1(_04647_),
    .A2(_04648_),
    .B1(_04650_),
    .Y(_04652_));
 sky130_fd_sc_hd__a211o_1 _32787_ (.A1(_04643_),
    .A2(_04644_),
    .B1(_04651_),
    .C1(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__o211ai_2 _32788_ (.A1(_04651_),
    .A2(_04652_),
    .B1(_04643_),
    .C1(_04644_),
    .Y(_04654_));
 sky130_fd_sc_hd__nand2_1 _32789_ (.A(_04653_),
    .B(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__a31o_1 _32790_ (.A1(_25310_),
    .A2(_01772_),
    .A3(_03371_),
    .B1(_03375_),
    .X(_04657_));
 sky130_fd_sc_hd__xnor2_1 _32791_ (.A(_04655_),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32792_ (.A(\delay_line[7][14] ),
    .X(_04659_));
 sky130_fd_sc_hd__or2b_1 _32793_ (.A(_01767_),
    .B_N(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__or2b_1 _32794_ (.A(_04659_),
    .B_N(_01767_),
    .X(_04661_));
 sky130_fd_sc_hd__and3_1 _32795_ (.A(_04660_),
    .B(_04661_),
    .C(_03335_),
    .X(_04662_));
 sky130_fd_sc_hd__a21oi_1 _32796_ (.A1(_04660_),
    .A2(_04661_),
    .B1(_03336_),
    .Y(_04663_));
 sky130_fd_sc_hd__or2_1 _32797_ (.A(_04662_),
    .B(_04663_),
    .X(_04664_));
 sky130_fd_sc_hd__a21oi_1 _32798_ (.A1(_03357_),
    .A2(_03364_),
    .B1(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__and3_1 _32799_ (.A(_03357_),
    .B(_03364_),
    .C(_04664_),
    .X(_04666_));
 sky130_fd_sc_hd__or3_1 _32800_ (.A(_03336_),
    .B(_03339_),
    .C(_01748_),
    .X(_04668_));
 sky130_fd_sc_hd__o21ai_1 _32801_ (.A1(_04665_),
    .A2(_04666_),
    .B1(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__or3_1 _32802_ (.A(_04668_),
    .B(_04665_),
    .C(_04666_),
    .X(_04670_));
 sky130_fd_sc_hd__nand3_1 _32803_ (.A(_04658_),
    .B(_04669_),
    .C(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__a21o_1 _32804_ (.A1(_04670_),
    .A2(_04669_),
    .B1(_04658_),
    .X(_04672_));
 sky130_fd_sc_hd__and2_1 _32805_ (.A(_04671_),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__nor3b_2 _32806_ (.A(_04631_),
    .B(_04632_),
    .C_N(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__o21bai_1 _32807_ (.A1(_04631_),
    .A2(_04632_),
    .B1_N(_04673_),
    .Y(_04675_));
 sky130_fd_sc_hd__inv_2 _32808_ (.A(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__a21oi_2 _32809_ (.A1(_03258_),
    .A2(_03295_),
    .B1(_03302_),
    .Y(_04677_));
 sky130_fd_sc_hd__o21ai_4 _32810_ (.A1(_04674_),
    .A2(_04676_),
    .B1(_04677_),
    .Y(_04679_));
 sky130_fd_sc_hd__or3_4 _32811_ (.A(_04677_),
    .B(_04674_),
    .C(_04676_),
    .X(_04680_));
 sky130_fd_sc_hd__and4_2 _32812_ (.A(_03333_),
    .B(_03385_),
    .C(_04679_),
    .D(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__a22oi_4 _32813_ (.A1(_03333_),
    .A2(_03385_),
    .B1(_04679_),
    .B2(_04680_),
    .Y(_04682_));
 sky130_fd_sc_hd__clkbuf_2 _32814_ (.A(_00076_),
    .X(_04683_));
 sky130_fd_sc_hd__clkbuf_2 _32815_ (.A(_03145_),
    .X(_04684_));
 sky130_fd_sc_hd__and2_1 _32816_ (.A(_00059_),
    .B(net395),
    .X(_04685_));
 sky130_fd_sc_hd__nor2_1 _32817_ (.A(_00060_),
    .B(net395),
    .Y(_04686_));
 sky130_fd_sc_hd__or2_1 _32818_ (.A(_04685_),
    .B(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__a21oi_4 _32819_ (.A1(_04683_),
    .A2(_04684_),
    .B1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__and3_2 _32820_ (.A(_04687_),
    .B(_04684_),
    .C(_04683_),
    .X(_04690_));
 sky130_fd_sc_hd__inv_2 _32821_ (.A(net453),
    .Y(_04691_));
 sky130_fd_sc_hd__inv_2 _32822_ (.A(_03181_),
    .Y(_04692_));
 sky130_fd_sc_hd__a21oi_2 _32823_ (.A1(_04691_),
    .A2(_03187_),
    .B1(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__nand2b_1 _32824_ (.A_N(_25416_),
    .B(_03160_),
    .Y(_04694_));
 sky130_fd_sc_hd__xnor2_2 _32825_ (.A(\delay_line[4][9] ),
    .B(\delay_line[4][11] ),
    .Y(_04695_));
 sky130_fd_sc_hd__o211a_1 _32826_ (.A1(_01575_),
    .A2(_03163_),
    .B1(_04694_),
    .C1(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__o21a_1 _32827_ (.A1(_03163_),
    .A2(_01575_),
    .B1(_04694_),
    .X(_04697_));
 sky130_fd_sc_hd__nor2_1 _32828_ (.A(_04695_),
    .B(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__nor2_1 _32829_ (.A(_04696_),
    .B(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__clkbuf_2 _32830_ (.A(_03160_),
    .X(_04701_));
 sky130_fd_sc_hd__nand4_2 _32831_ (.A(_04701_),
    .B(_03165_),
    .C(_01576_),
    .D(_01573_),
    .Y(_04702_));
 sky130_fd_sc_hd__nand3_2 _32832_ (.A(_03185_),
    .B(_04699_),
    .C(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__and3_1 _32833_ (.A(_04701_),
    .B(_01573_),
    .C(_01579_),
    .X(_04704_));
 sky130_fd_sc_hd__o22ai_4 _32834_ (.A1(_04696_),
    .A2(_04698_),
    .B1(_04704_),
    .B2(_03173_),
    .Y(_04705_));
 sky130_fd_sc_hd__nor2b_1 _32835_ (.A(_22308_),
    .B_N(net410),
    .Y(_04706_));
 sky130_fd_sc_hd__and2b_1 _32836_ (.A_N(net410),
    .B(_22308_),
    .X(_04707_));
 sky130_fd_sc_hd__or2_2 _32837_ (.A(_04706_),
    .B(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__nand4_2 _32838_ (.A(_01560_),
    .B(_01562_),
    .C(_03155_),
    .D(_03156_),
    .Y(_04709_));
 sky130_fd_sc_hd__nor2b_2 _32839_ (.A(_23839_),
    .B_N(\delay_line[11][12] ),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2b_1 _32840_ (.A_N(\delay_line[11][12] ),
    .B(_23839_),
    .Y(_04712_));
 sky130_fd_sc_hd__nor2b_4 _32841_ (.A(_04710_),
    .B_N(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__a21oi_2 _32842_ (.A1(_01554_),
    .A2(_03153_),
    .B1(_04706_),
    .Y(_04714_));
 sky130_fd_sc_hd__xor2_4 _32843_ (.A(_04713_),
    .B(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__o221a_1 _32844_ (.A1(_01563_),
    .A2(_04708_),
    .B1(_04709_),
    .B2(_01570_),
    .C1(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__o22ai_4 _32845_ (.A1(_01563_),
    .A2(_04708_),
    .B1(_04709_),
    .B2(_01569_),
    .Y(_04717_));
 sky130_fd_sc_hd__inv_2 _32846_ (.A(_04715_),
    .Y(_04718_));
 sky130_fd_sc_hd__nand2_1 _32847_ (.A(_04717_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__inv_2 _32848_ (.A(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__o2bb2ai_2 _32849_ (.A1_N(_04703_),
    .A2_N(_04705_),
    .B1(_04716_),
    .B2(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nor2b_1 _32850_ (.A(_04716_),
    .B_N(_04719_),
    .Y(_04723_));
 sky130_fd_sc_hd__nand3_2 _32851_ (.A(_04703_),
    .B(_04705_),
    .C(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__a21o_1 _32852_ (.A1(_04721_),
    .A2(_04724_),
    .B1(net452),
    .X(_04725_));
 sky130_fd_sc_hd__nand3_1 _32853_ (.A(_04721_),
    .B(_04724_),
    .C(net452),
    .Y(_04726_));
 sky130_fd_sc_hd__nand3_1 _32854_ (.A(_04693_),
    .B(_04725_),
    .C(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__o41a_1 _32855_ (.A1(_03158_),
    .A2(_03159_),
    .A3(_03173_),
    .A4(_03180_),
    .B1(_04691_),
    .X(_04728_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32856_ (.A(net452),
    .X(_04729_));
 sky130_fd_sc_hd__a21oi_2 _32857_ (.A1(_04721_),
    .A2(_04724_),
    .B1(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__and3_1 _32858_ (.A(_04721_),
    .B(_04724_),
    .C(_04729_),
    .X(_04731_));
 sky130_fd_sc_hd__o22ai_2 _32859_ (.A1(_04692_),
    .A2(_04728_),
    .B1(_04730_),
    .B2(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__clkbuf_2 _32860_ (.A(_03198_),
    .X(_04734_));
 sky130_fd_sc_hd__a21oi_1 _32861_ (.A1(_04727_),
    .A2(_04732_),
    .B1(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__buf_4 _32862_ (.A(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__nand3_2 _32863_ (.A(_04732_),
    .B(_03198_),
    .C(_04727_),
    .Y(_04737_));
 sky130_fd_sc_hd__a2bb2o_2 _32864_ (.A1_N(_03188_),
    .A2_N(_03190_),
    .B1(_03206_),
    .B2(_03195_),
    .X(_04738_));
 sky130_fd_sc_hd__nand2_2 _32865_ (.A(_04737_),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__nor2_1 _32866_ (.A(_04736_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__nand2_1 _32867_ (.A(_04693_),
    .B(_04726_),
    .Y(_04741_));
 sky130_fd_sc_hd__nor2_1 _32868_ (.A(_04730_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__a21oi_2 _32869_ (.A1(_04725_),
    .A2(_04726_),
    .B1(_04693_),
    .Y(_04743_));
 sky130_fd_sc_hd__clkbuf_2 _32870_ (.A(_04691_),
    .X(_04745_));
 sky130_fd_sc_hd__o21ai_2 _32871_ (.A1(_04742_),
    .A2(_04743_),
    .B1(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__a21oi_4 _32872_ (.A1(_04746_),
    .A2(_04737_),
    .B1(_04738_),
    .Y(_04747_));
 sky130_fd_sc_hd__o22ai_4 _32873_ (.A1(_04688_),
    .A2(_04690_),
    .B1(_04740_),
    .B2(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__o2bb2a_1 _32874_ (.A1_N(_03211_),
    .A2_N(_03212_),
    .B1(_03208_),
    .B2(_03207_),
    .X(_04749_));
 sky130_fd_sc_hd__nor2_2 _32875_ (.A(_04688_),
    .B(_04690_),
    .Y(_04750_));
 sky130_fd_sc_hd__clkbuf_2 _32876_ (.A(_01626_),
    .X(_04751_));
 sky130_fd_sc_hd__o41a_1 _32877_ (.A1(_01590_),
    .A2(_01609_),
    .A3(_03188_),
    .A4(_03192_),
    .B1(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__o311a_1 _32878_ (.A1(_04692_),
    .A2(_04730_),
    .A3(_04731_),
    .B1(_04734_),
    .C1(_04732_),
    .X(_04753_));
 sky130_fd_sc_hd__o22ai_4 _32879_ (.A1(_03200_),
    .A2(_04752_),
    .B1(_04736_),
    .B2(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__o211ai_4 _32880_ (.A1(_04739_),
    .A2(_04736_),
    .B1(_04750_),
    .C1(_04754_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand3_2 _32881_ (.A(_04748_),
    .B(_04749_),
    .C(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__nor4_1 _32882_ (.A(_22363_),
    .B(_03144_),
    .C(_01548_),
    .D(_03149_),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_1 _32883_ (.A(_22363_),
    .B(_01547_),
    .Y(_04759_));
 sky130_fd_sc_hd__or2_1 _32884_ (.A(_22362_),
    .B(_01547_),
    .X(_04760_));
 sky130_fd_sc_hd__a21oi_1 _32885_ (.A1(_04759_),
    .A2(_04760_),
    .B1(_03147_),
    .Y(_04761_));
 sky130_fd_sc_hd__clkbuf_2 _32886_ (.A(_01549_),
    .X(_04762_));
 sky130_fd_sc_hd__and4bb_1 _32887_ (.A_N(_04758_),
    .B_N(_04761_),
    .C(_23811_),
    .D(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__o2bb2a_1 _32888_ (.A1_N(_23812_),
    .A2_N(_04762_),
    .B1(_04758_),
    .B2(_04761_),
    .X(_04764_));
 sky130_fd_sc_hd__or2_2 _32889_ (.A(_04763_),
    .B(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__inv_2 _32890_ (.A(_04765_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_1 _32891_ (.A(_04757_),
    .B(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__o211a_1 _32892_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03211_),
    .C1(_03212_),
    .X(_04769_));
 sky130_fd_sc_hd__o221ai_4 _32893_ (.A1(_04688_),
    .A2(_04690_),
    .B1(_04736_),
    .B2(_04739_),
    .C1(_04754_),
    .Y(_04770_));
 sky130_fd_sc_hd__clkbuf_2 _32894_ (.A(_04684_),
    .X(_04771_));
 sky130_fd_sc_hd__buf_1 _32895_ (.A(_04685_),
    .X(_04772_));
 sky130_fd_sc_hd__nor2_1 _32896_ (.A(_04772_),
    .B(_04686_),
    .Y(_04773_));
 sky130_fd_sc_hd__and3_1 _32897_ (.A(_04683_),
    .B(_04771_),
    .C(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__buf_2 _32898_ (.A(_04771_),
    .X(_04775_));
 sky130_fd_sc_hd__o2bb2a_1 _32899_ (.A1_N(_04683_),
    .A2_N(_04775_),
    .B1(_04772_),
    .B2(_04686_),
    .X(_04776_));
 sky130_fd_sc_hd__o22ai_2 _32900_ (.A1(_04774_),
    .A2(_04776_),
    .B1(_04740_),
    .B2(_04747_),
    .Y(_04778_));
 sky130_fd_sc_hd__o211a_2 _32901_ (.A1(_03209_),
    .A2(_04769_),
    .B1(_04770_),
    .C1(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__nor2_1 _32902_ (.A(_03231_),
    .B(_03232_),
    .Y(_04780_));
 sky130_fd_sc_hd__a32o_1 _32903_ (.A1(_03143_),
    .A2(_03210_),
    .A3(_03213_),
    .B1(_03233_),
    .B2(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__o211ai_2 _32904_ (.A1(_03209_),
    .A2(_04769_),
    .B1(_04770_),
    .C1(_04778_),
    .Y(_04782_));
 sky130_fd_sc_hd__o2bb2ai_1 _32905_ (.A1_N(_04782_),
    .A2_N(_04757_),
    .B1(_04763_),
    .B2(_04764_),
    .Y(_04783_));
 sky130_fd_sc_hd__o211ai_2 _32906_ (.A1(_04768_),
    .A2(_04779_),
    .B1(_04781_),
    .C1(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__or2_1 _32907_ (.A(net270),
    .B(_04761_),
    .X(_04785_));
 sky130_fd_sc_hd__clkbuf_2 _32908_ (.A(_04762_),
    .X(_04786_));
 sky130_fd_sc_hd__and3_1 _32909_ (.A(_04785_),
    .B(_04786_),
    .C(_23898_),
    .X(_04787_));
 sky130_fd_sc_hd__buf_2 _32910_ (.A(_04786_),
    .X(_04789_));
 sky130_fd_sc_hd__a21oi_1 _32911_ (.A1(_23898_),
    .A2(_04789_),
    .B1(_04785_),
    .Y(_04790_));
 sky130_fd_sc_hd__o2bb2ai_1 _32912_ (.A1_N(_04782_),
    .A2_N(_04757_),
    .B1(_04787_),
    .B2(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__a32oi_2 _32913_ (.A1(_03143_),
    .A2(_03210_),
    .A3(_03213_),
    .B1(_03233_),
    .B2(_04780_),
    .Y(_04792_));
 sky130_fd_sc_hd__o211ai_1 _32914_ (.A1(_04763_),
    .A2(_04764_),
    .B1(_04782_),
    .C1(_04757_),
    .Y(_04793_));
 sky130_fd_sc_hd__nand3_2 _32915_ (.A(_04791_),
    .B(_04792_),
    .C(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand2_1 _32916_ (.A(_04784_),
    .B(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__clkbuf_2 _32917_ (.A(\delay_line[12][14] ),
    .X(_04796_));
 sky130_fd_sc_hd__nor2_2 _32918_ (.A(\delay_line[12][13] ),
    .B(net400),
    .Y(_04797_));
 sky130_fd_sc_hd__inv_2 _32919_ (.A(net401),
    .Y(_04798_));
 sky130_fd_sc_hd__inv_2 _32920_ (.A(net400),
    .Y(_04800_));
 sky130_fd_sc_hd__nor2_2 _32921_ (.A(_04798_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__o21ai_1 _32922_ (.A1(_04797_),
    .A2(_04801_),
    .B1(_03126_),
    .Y(_04802_));
 sky130_fd_sc_hd__o211a_1 _32923_ (.A1(_04796_),
    .A2(_03126_),
    .B1(_25373_),
    .C1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__o21a_1 _32924_ (.A1(net400),
    .A2(_03126_),
    .B1(_04802_),
    .X(_04804_));
 sky130_fd_sc_hd__nor2_1 _32925_ (.A(_25373_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__o21bai_1 _32926_ (.A1(_04803_),
    .A2(_04805_),
    .B1_N(_03220_),
    .Y(_04806_));
 sky130_fd_sc_hd__or3b_2 _32927_ (.A(_04803_),
    .B(_04805_),
    .C_N(_18918_),
    .X(_04807_));
 sky130_fd_sc_hd__a31o_1 _32928_ (.A1(_03220_),
    .A2(_00093_),
    .A3(_03225_),
    .B1(_03223_),
    .X(_04808_));
 sky130_fd_sc_hd__and3_1 _32929_ (.A(_04806_),
    .B(_04807_),
    .C(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__a21oi_1 _32930_ (.A1(_04806_),
    .A2(_04807_),
    .B1(_04808_),
    .Y(_04811_));
 sky130_fd_sc_hd__nor2_1 _32931_ (.A(_04809_),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__and4bb_1 _32932_ (.A_N(_03133_),
    .B_N(_03134_),
    .C(_04812_),
    .D(_00099_),
    .X(_04813_));
 sky130_fd_sc_hd__nor2_1 _32933_ (.A(_03135_),
    .B(_04812_),
    .Y(_04814_));
 sky130_fd_sc_hd__nor2_1 _32934_ (.A(_04813_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_1 _32935_ (.A(_04795_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__nor2_1 _32936_ (.A(_03248_),
    .B(_03250_),
    .Y(_04817_));
 sky130_fd_sc_hd__a32oi_4 _32937_ (.A1(_03239_),
    .A2(_03240_),
    .A3(_03241_),
    .B1(_03236_),
    .B2(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__nand3b_1 _32938_ (.A_N(_04815_),
    .B(_04784_),
    .C(_04794_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand3_4 _32939_ (.A(_04816_),
    .B(_04818_),
    .C(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__clkbuf_2 _32940_ (.A(_04784_),
    .X(_04822_));
 sky130_fd_sc_hd__buf_6 _32941_ (.A(_04794_),
    .X(_04823_));
 sky130_fd_sc_hd__buf_2 _32942_ (.A(_04815_),
    .X(_04824_));
 sky130_fd_sc_hd__a31oi_1 _32943_ (.A1(_04822_),
    .A2(_04823_),
    .A3(_04824_),
    .B1(_04818_),
    .Y(_04825_));
 sky130_fd_sc_hd__a21o_1 _32944_ (.A1(_04822_),
    .A2(_04823_),
    .B1(_04824_),
    .X(_04826_));
 sky130_fd_sc_hd__nand2_1 _32945_ (.A(_04825_),
    .B(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__clkbuf_2 _32946_ (.A(\delay_line[9][14] ),
    .X(_04828_));
 sky130_fd_sc_hd__or2b_1 _32947_ (.A(_22447_),
    .B_N(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__or2b_1 _32948_ (.A(\delay_line[9][14] ),
    .B_N(_19964_),
    .X(_04830_));
 sky130_fd_sc_hd__a22o_1 _32949_ (.A1(_04611_),
    .A2(_21801_),
    .B1(_04829_),
    .B2(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__and2b_1 _32950_ (.A_N(_17921_),
    .B(_04614_),
    .X(_04833_));
 sky130_fd_sc_hd__nand4_1 _32951_ (.A(_04829_),
    .B(_04830_),
    .C(_04611_),
    .D(_22458_),
    .Y(_04834_));
 sky130_fd_sc_hd__and3_1 _32952_ (.A(_04831_),
    .B(_04833_),
    .C(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__a21oi_1 _32953_ (.A1(_04834_),
    .A2(_04831_),
    .B1(_04833_),
    .Y(_04836_));
 sky130_fd_sc_hd__nor2_1 _32954_ (.A(_22456_),
    .B(_01692_),
    .Y(_04837_));
 sky130_fd_sc_hd__and2_1 _32955_ (.A(_21800_),
    .B(_23771_),
    .X(_04838_));
 sky130_fd_sc_hd__or3b_1 _32956_ (.A(_04837_),
    .B(_04838_),
    .C_N(_25370_),
    .X(_04839_));
 sky130_fd_sc_hd__buf_1 _32957_ (.A(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__o21bai_1 _32958_ (.A1(_04837_),
    .A2(_04838_),
    .B1_N(_25376_),
    .Y(_04841_));
 sky130_fd_sc_hd__buf_1 _32959_ (.A(\delay_line[10][10] ),
    .X(_04842_));
 sky130_fd_sc_hd__clkbuf_2 _32960_ (.A(_04842_),
    .X(_04844_));
 sky130_fd_sc_hd__nor2_1 _32961_ (.A(_03267_),
    .B(_03268_),
    .Y(_04845_));
 sky130_fd_sc_hd__and4_1 _32962_ (.A(_04840_),
    .B(_04841_),
    .C(_04844_),
    .D(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__a22oi_2 _32963_ (.A1(_04844_),
    .A2(_04845_),
    .B1(_04840_),
    .B2(_04841_),
    .Y(_04847_));
 sky130_fd_sc_hd__or4_1 _32964_ (.A(_04835_),
    .B(_04836_),
    .C(_04846_),
    .D(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__o22ai_1 _32965_ (.A1(_04835_),
    .A2(_04836_),
    .B1(_04846_),
    .B2(_04847_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_1 _32966_ (.A(_04848_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand3_1 _32967_ (.A(_03277_),
    .B(_03280_),
    .C(_03284_),
    .Y(_04851_));
 sky130_fd_sc_hd__and3_1 _32968_ (.A(_04798_),
    .B(net402),
    .C(_00120_),
    .X(_04852_));
 sky130_fd_sc_hd__o211a_1 _32969_ (.A1(net402),
    .A2(net401),
    .B1(_22465_),
    .C1(_03127_),
    .X(_04853_));
 sky130_fd_sc_hd__and2_1 _32970_ (.A(_22392_),
    .B(\delay_line[10][14] ),
    .X(_04855_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _32971_ (.A(\delay_line[10][14] ),
    .X(_04856_));
 sky130_fd_sc_hd__nor2_1 _32972_ (.A(_22392_),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__or3b_1 _32973_ (.A(_04855_),
    .B(_04857_),
    .C_N(_03278_),
    .X(_04858_));
 sky130_fd_sc_hd__a2bb2o_1 _32974_ (.A1_N(_04855_),
    .A2_N(_04857_),
    .B1(_20062_),
    .B2(net411),
    .X(_04859_));
 sky130_fd_sc_hd__o211a_1 _32975_ (.A1(_04852_),
    .A2(_04853_),
    .B1(_04858_),
    .C1(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__a221oi_2 _32976_ (.A1(_25372_),
    .A2(_03129_),
    .B1(_04858_),
    .B2(_04859_),
    .C1(_04852_),
    .Y(_04861_));
 sky130_fd_sc_hd__o21a_1 _32977_ (.A1(_04860_),
    .A2(_04861_),
    .B1(_03280_),
    .X(_04862_));
 sky130_fd_sc_hd__nor3_1 _32978_ (.A(_03280_),
    .B(_04860_),
    .C(_04861_),
    .Y(_04863_));
 sky130_fd_sc_hd__a211o_1 _32979_ (.A1(_04851_),
    .A2(_03288_),
    .B1(_04862_),
    .C1(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__o221ai_1 _32980_ (.A1(_03286_),
    .A2(_01711_),
    .B1(_04863_),
    .B2(_04862_),
    .C1(_04851_),
    .Y(_04866_));
 sky130_fd_sc_hd__nand2_1 _32981_ (.A(_04864_),
    .B(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__xnor2_1 _32982_ (.A(_04850_),
    .B(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__o21ba_1 _32983_ (.A1(_03137_),
    .A2(_03248_),
    .B1_N(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__nor3b_1 _32984_ (.A(_03137_),
    .B(_03248_),
    .C_N(_04868_),
    .Y(_04870_));
 sky130_fd_sc_hd__nor2_2 _32985_ (.A(_04869_),
    .B(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__a32o_2 _32986_ (.A1(_03274_),
    .A2(_03275_),
    .A3(_03290_),
    .B1(_03287_),
    .B2(_03289_),
    .X(_04872_));
 sky130_fd_sc_hd__xor2_4 _32987_ (.A(_04871_),
    .B(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__a21oi_2 _32988_ (.A1(_04820_),
    .A2(_04827_),
    .B1(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__buf_4 _32989_ (.A(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__o21a_1 _32990_ (.A1(_03298_),
    .A2(_03299_),
    .B1(_03256_),
    .X(_04877_));
 sky130_fd_sc_hd__a21oi_4 _32991_ (.A1(_04822_),
    .A2(_04823_),
    .B1(_04824_),
    .Y(_04878_));
 sky130_fd_sc_hd__a32o_1 _32992_ (.A1(_03239_),
    .A2(_03240_),
    .A3(_03241_),
    .B1(_03236_),
    .B2(_04817_),
    .X(_04879_));
 sky130_fd_sc_hd__nand3_1 _32993_ (.A(_04822_),
    .B(_04794_),
    .C(_04815_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_2 _32994_ (.A(_04879_),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__o211ai_4 _32995_ (.A1(_04878_),
    .A2(_04881_),
    .B1(_04873_),
    .C1(_04820_),
    .Y(_04882_));
 sky130_fd_sc_hd__o21ai_4 _32996_ (.A1(_03396_),
    .A2(_04877_),
    .B1(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__o211a_1 _32997_ (.A1(_04878_),
    .A2(_04881_),
    .B1(_04873_),
    .C1(_04820_),
    .X(_04884_));
 sky130_fd_sc_hd__a21o_1 _32998_ (.A1(_03257_),
    .A2(_03394_),
    .B1(_03396_),
    .X(_04885_));
 sky130_fd_sc_hd__o21bai_4 _32999_ (.A1(_04875_),
    .A2(_04884_),
    .B1_N(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__o221ai_4 _33000_ (.A1(_04681_),
    .A2(_04682_),
    .B1(_04875_),
    .B2(_04883_),
    .C1(_04886_),
    .Y(_04888_));
 sky130_fd_sc_hd__nand2_1 _33001_ (.A(_03333_),
    .B(_03385_),
    .Y(_04889_));
 sky130_fd_sc_hd__and3_1 _33002_ (.A(_04889_),
    .B(_04679_),
    .C(_04680_),
    .X(_04890_));
 sky130_fd_sc_hd__a21oi_2 _33003_ (.A1(_04679_),
    .A2(_04680_),
    .B1(_04889_),
    .Y(_04891_));
 sky130_fd_sc_hd__nor2_1 _33004_ (.A(_04875_),
    .B(_04883_),
    .Y(_04892_));
 sky130_fd_sc_hd__inv_2 _33005_ (.A(_04873_),
    .Y(_04893_));
 sky130_fd_sc_hd__o21ai_1 _33006_ (.A1(_04878_),
    .A2(_04881_),
    .B1(_04820_),
    .Y(_04894_));
 sky130_fd_sc_hd__nand2_1 _33007_ (.A(_04893_),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__a21oi_4 _33008_ (.A1(_04895_),
    .A2(_04882_),
    .B1(_04885_),
    .Y(_04896_));
 sky130_fd_sc_hd__o22ai_2 _33009_ (.A1(_04890_),
    .A2(_04891_),
    .B1(_04892_),
    .B2(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__o211ai_4 _33010_ (.A1(_03399_),
    .A2(_04608_),
    .B1(_04888_),
    .C1(_04897_),
    .Y(_04899_));
 sky130_fd_sc_hd__o22ai_2 _33011_ (.A1(_04681_),
    .A2(_04682_),
    .B1(_04892_),
    .B2(_04896_),
    .Y(_04900_));
 sky130_fd_sc_hd__o221ai_4 _33012_ (.A1(_04890_),
    .A2(_04891_),
    .B1(_04875_),
    .B2(_04883_),
    .C1(_04886_),
    .Y(_04901_));
 sky130_fd_sc_hd__a21oi_2 _33013_ (.A1(_03307_),
    .A2(_03391_),
    .B1(_03399_),
    .Y(_04902_));
 sky130_fd_sc_hd__nand3_4 _33014_ (.A(_04900_),
    .B(_04901_),
    .C(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__o21ba_2 _33015_ (.A1(_03440_),
    .A2(_03499_),
    .B1_N(_03441_),
    .X(_04904_));
 sky130_fd_sc_hd__o21bai_4 _33016_ (.A1(_03308_),
    .A2(_03386_),
    .B1_N(_03384_),
    .Y(_04905_));
 sky130_fd_sc_hd__nor2_1 _33017_ (.A(_03490_),
    .B(_03493_),
    .Y(_04906_));
 sky130_fd_sc_hd__and4b_1 _33018_ (.A_N(_19883_),
    .B(_03485_),
    .C(_03483_),
    .D(_01861_),
    .X(_04907_));
 sky130_fd_sc_hd__buf_1 _33019_ (.A(\delay_line[2][14] ),
    .X(_04908_));
 sky130_fd_sc_hd__or2b_1 _33020_ (.A(_01861_),
    .B_N(_04908_),
    .X(_04910_));
 sky130_fd_sc_hd__or2b_1 _33021_ (.A(\delay_line[2][14] ),
    .B_N(_01861_),
    .X(_04911_));
 sky130_fd_sc_hd__a22o_1 _33022_ (.A1(_22642_),
    .A2(_03454_),
    .B1(_04910_),
    .B2(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__nand4_1 _33023_ (.A(_22642_),
    .B(_04910_),
    .C(_04911_),
    .D(_03454_),
    .Y(_04913_));
 sky130_fd_sc_hd__and3_1 _33024_ (.A(_04912_),
    .B(_03482_),
    .C(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__a21oi_1 _33025_ (.A1(_04913_),
    .A2(_04912_),
    .B1(_03482_),
    .Y(_04915_));
 sky130_fd_sc_hd__nor2_1 _33026_ (.A(_04914_),
    .B(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__xnor2_1 _33027_ (.A(_03459_),
    .B(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__or3_1 _33028_ (.A(_04907_),
    .B(_03489_),
    .C(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__o21ai_1 _33029_ (.A1(_04907_),
    .A2(_03489_),
    .B1(_04917_),
    .Y(_04919_));
 sky130_fd_sc_hd__a211oi_1 _33030_ (.A1(_04918_),
    .A2(_04919_),
    .B1(_03451_),
    .C1(_03461_),
    .Y(_04921_));
 sky130_fd_sc_hd__o211ai_2 _33031_ (.A1(_03451_),
    .A2(_03461_),
    .B1(_04918_),
    .C1(_04919_),
    .Y(_04922_));
 sky130_fd_sc_hd__and2b_1 _33032_ (.A_N(_04921_),
    .B(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__xor2_2 _33033_ (.A(_04906_),
    .B(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__a21oi_2 _33034_ (.A1(_03463_),
    .A2(_03477_),
    .B1(_03476_),
    .Y(_04925_));
 sky130_fd_sc_hd__or2_1 _33035_ (.A(_03465_),
    .B(_03472_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_2 _33036_ (.A(_01924_),
    .X(_04927_));
 sky130_fd_sc_hd__buf_2 _33037_ (.A(_03424_),
    .X(_04928_));
 sky130_fd_sc_hd__o21a_1 _33038_ (.A1(_01888_),
    .A2(_04927_),
    .B1(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__nor3_1 _33039_ (.A(_03464_),
    .B(_04927_),
    .C(_04928_),
    .Y(_04930_));
 sky130_fd_sc_hd__a211o_1 _33040_ (.A1(_03422_),
    .A2(_03426_),
    .B1(_04929_),
    .C1(_04930_),
    .X(_04932_));
 sky130_fd_sc_hd__clkbuf_2 _33041_ (.A(_04927_),
    .X(_04933_));
 sky130_fd_sc_hd__o21a_1 _33042_ (.A1(_03464_),
    .A2(_04933_),
    .B1(_01885_),
    .X(_04934_));
 sky130_fd_sc_hd__o211ai_2 _33043_ (.A1(_04929_),
    .A2(_04930_),
    .B1(_03422_),
    .C1(_03426_),
    .Y(_04935_));
 sky130_fd_sc_hd__and3_1 _33044_ (.A(_04932_),
    .B(_04934_),
    .C(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__a21oi_1 _33045_ (.A1(_04935_),
    .A2(_04932_),
    .B1(_04934_),
    .Y(_04937_));
 sky130_fd_sc_hd__a211o_1 _33046_ (.A1(_03471_),
    .A2(_04926_),
    .B1(_04936_),
    .C1(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__o221ai_2 _33047_ (.A1(_03465_),
    .A2(_03472_),
    .B1(_04936_),
    .B2(_04937_),
    .C1(_03471_),
    .Y(_04939_));
 sky130_fd_sc_hd__buf_1 _33048_ (.A(_21962_),
    .X(_04940_));
 sky130_fd_sc_hd__clkbuf_2 _33049_ (.A(net435),
    .X(_04941_));
 sky130_fd_sc_hd__nand2_1 _33050_ (.A(_04940_),
    .B(_04941_),
    .Y(_04943_));
 sky130_fd_sc_hd__or2_1 _33051_ (.A(net435),
    .B(_04940_),
    .X(_04944_));
 sky130_fd_sc_hd__clkbuf_2 _33052_ (.A(_01869_),
    .X(_04945_));
 sky130_fd_sc_hd__a21oi_1 _33053_ (.A1(_04943_),
    .A2(_04944_),
    .B1(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__and3_1 _33054_ (.A(_04944_),
    .B(_04945_),
    .C(_04943_),
    .X(_04947_));
 sky130_fd_sc_hd__nor2_1 _33055_ (.A(_04946_),
    .B(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand3_1 _33056_ (.A(_03446_),
    .B(_03444_),
    .C(_01869_),
    .Y(_04949_));
 sky130_fd_sc_hd__or2b_1 _33057_ (.A(_19904_),
    .B_N(\delay_line[5][14] ),
    .X(_04950_));
 sky130_fd_sc_hd__or2b_1 _33058_ (.A(\delay_line[5][14] ),
    .B_N(_19904_),
    .X(_04951_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33059_ (.A(\delay_line[5][13] ),
    .X(_04952_));
 sky130_fd_sc_hd__and3_1 _33060_ (.A(_04950_),
    .B(_04951_),
    .C(_04952_),
    .X(_04954_));
 sky130_fd_sc_hd__a21oi_1 _33061_ (.A1(_04950_),
    .A2(_04951_),
    .B1(_04952_),
    .Y(_04955_));
 sky130_fd_sc_hd__a211oi_2 _33062_ (.A1(_03446_),
    .A2(_04949_),
    .B1(_04954_),
    .C1(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__o211ai_1 _33063_ (.A1(_04954_),
    .A2(_04955_),
    .B1(_03446_),
    .C1(_04949_),
    .Y(_04957_));
 sky130_fd_sc_hd__nand3b_1 _33064_ (.A_N(_04956_),
    .B(_04957_),
    .C(_03449_),
    .Y(_04958_));
 sky130_fd_sc_hd__o211a_1 _33065_ (.A1(_04954_),
    .A2(_04955_),
    .B1(_03446_),
    .C1(_04949_),
    .X(_04959_));
 sky130_fd_sc_hd__o21bai_1 _33066_ (.A1(_04956_),
    .A2(_04959_),
    .B1_N(_03449_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand2_1 _33067_ (.A(_04958_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__xnor2_1 _33068_ (.A(_04948_),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__nand3_1 _33069_ (.A(_04938_),
    .B(_04939_),
    .C(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__a21o_1 _33070_ (.A1(_04938_),
    .A2(_04939_),
    .B1(_04962_),
    .X(_04965_));
 sky130_fd_sc_hd__and2_1 _33071_ (.A(_04963_),
    .B(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__xor2_2 _33072_ (.A(_04925_),
    .B(_04966_),
    .X(_04967_));
 sky130_fd_sc_hd__xnor2_2 _33073_ (.A(_04924_),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__o21a_1 _33074_ (.A1(_01929_),
    .A2(_03432_),
    .B1(_03431_),
    .X(_04969_));
 sky130_fd_sc_hd__and2_1 _33075_ (.A(_03376_),
    .B(_03350_),
    .X(_04970_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33076_ (.A(_03413_),
    .X(_04971_));
 sky130_fd_sc_hd__nor2_1 _33077_ (.A(_04971_),
    .B(_01909_),
    .Y(_04972_));
 sky130_fd_sc_hd__buf_1 _33078_ (.A(\delay_line[7][10] ),
    .X(_04973_));
 sky130_fd_sc_hd__and2_1 _33079_ (.A(_22525_),
    .B(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__o21bai_2 _33080_ (.A1(_04972_),
    .A2(_04974_),
    .B1_N(_03412_),
    .Y(_04976_));
 sky130_fd_sc_hd__or3b_2 _33081_ (.A(_04972_),
    .B(_04974_),
    .C_N(_03412_),
    .X(_04977_));
 sky130_fd_sc_hd__clkbuf_2 _33082_ (.A(\delay_line[6][14] ),
    .X(_04978_));
 sky130_fd_sc_hd__or2b_1 _33083_ (.A(_00253_),
    .B_N(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__inv_2 _33084_ (.A(\delay_line[6][14] ),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2_1 _33085_ (.A(_04980_),
    .B(_01915_),
    .Y(_04981_));
 sky130_fd_sc_hd__o21a_1 _33086_ (.A1(_22527_),
    .A2(_03413_),
    .B1(_01912_),
    .X(_04982_));
 sky130_fd_sc_hd__a221o_1 _33087_ (.A1(_03412_),
    .A2(_03413_),
    .B1(_04979_),
    .B2(_04981_),
    .C1(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__o211ai_4 _33088_ (.A1(_03416_),
    .A2(_04982_),
    .B1(_04979_),
    .C1(_04981_),
    .Y(_04984_));
 sky130_fd_sc_hd__nand3_2 _33089_ (.A(_04983_),
    .B(_04984_),
    .C(_03420_),
    .Y(_04985_));
 sky130_fd_sc_hd__a21o_1 _33090_ (.A1(_04983_),
    .A2(_04984_),
    .B1(_03420_),
    .X(_04987_));
 sky130_fd_sc_hd__nand4_4 _33091_ (.A(_04976_),
    .B(_04977_),
    .C(_04985_),
    .D(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__a22o_1 _33092_ (.A1(_04976_),
    .A2(_04977_),
    .B1(_04985_),
    .B2(_04987_),
    .X(_04989_));
 sky130_fd_sc_hd__a211oi_2 _33093_ (.A1(_04988_),
    .A2(_04989_),
    .B1(_03344_),
    .C1(_03345_),
    .Y(_04990_));
 sky130_fd_sc_hd__o211a_1 _33094_ (.A1(_03344_),
    .A2(_03345_),
    .B1(_04988_),
    .C1(_04989_),
    .X(_04991_));
 sky130_fd_sc_hd__or3_2 _33095_ (.A(_04990_),
    .B(_03428_),
    .C(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__o21ai_2 _33096_ (.A1(_04991_),
    .A2(_04990_),
    .B1(_03428_),
    .Y(_04993_));
 sky130_fd_sc_hd__o211a_1 _33097_ (.A1(_04970_),
    .A2(_03378_),
    .B1(_04992_),
    .C1(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__a221oi_4 _33098_ (.A1(_03350_),
    .A2(_03376_),
    .B1(_04992_),
    .B2(_04993_),
    .C1(_03378_),
    .Y(_04995_));
 sky130_fd_sc_hd__or3_1 _33099_ (.A(_04969_),
    .B(_04994_),
    .C(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__o21ai_2 _33100_ (.A1(_04994_),
    .A2(_04995_),
    .B1(_04969_),
    .Y(_04998_));
 sky130_fd_sc_hd__a21o_1 _33101_ (.A1(_03433_),
    .A2(_03434_),
    .B1(_03437_),
    .X(_04999_));
 sky130_fd_sc_hd__a21oi_2 _33102_ (.A1(_04996_),
    .A2(_04998_),
    .B1(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand3_2 _33103_ (.A(_04999_),
    .B(_04996_),
    .C(_04998_),
    .Y(_05001_));
 sky130_fd_sc_hd__or2b_1 _33104_ (.A(_05000_),
    .B_N(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__xor2_2 _33105_ (.A(_04968_),
    .B(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__xnor2_2 _33106_ (.A(_04905_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__xor2_2 _33107_ (.A(_04904_),
    .B(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__a21oi_2 _33108_ (.A1(_04899_),
    .A2(_04903_),
    .B1(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__a311oi_2 _33109_ (.A1(_03405_),
    .A2(_03406_),
    .A3(_03407_),
    .B1(_03508_),
    .C1(_03509_),
    .Y(_05007_));
 sky130_fd_sc_hd__nand3_1 _33110_ (.A(_04899_),
    .B(_04903_),
    .C(_05005_),
    .Y(_05009_));
 sky130_fd_sc_hd__o21ai_2 _33111_ (.A1(_03516_),
    .A2(_05007_),
    .B1(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__nor2_2 _33112_ (.A(_05006_),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__nand2_1 _33113_ (.A(_04899_),
    .B(_04903_),
    .Y(_05012_));
 sky130_fd_sc_hd__inv_2 _33114_ (.A(_05005_),
    .Y(_05013_));
 sky130_fd_sc_hd__nand2_1 _33115_ (.A(_05012_),
    .B(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__a21o_1 _33116_ (.A1(_03408_),
    .A2(_03511_),
    .B1(_03516_),
    .X(_05015_));
 sky130_fd_sc_hd__a21oi_2 _33117_ (.A1(_05014_),
    .A2(_05009_),
    .B1(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__o21ai_4 _33118_ (.A1(_03108_),
    .A2(_03109_),
    .B1(_03112_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_1 _33119_ (.A(_03099_),
    .B(_03101_),
    .Y(_05018_));
 sky130_fd_sc_hd__o21a_1 _33120_ (.A1(_00324_),
    .A2(_03090_),
    .B1(_03092_),
    .X(_05020_));
 sky130_fd_sc_hd__and2b_1 _33121_ (.A_N(_03088_),
    .B(_03096_),
    .X(_05021_));
 sky130_fd_sc_hd__inv_2 _33122_ (.A(net446),
    .Y(_05022_));
 sky130_fd_sc_hd__or2_1 _33123_ (.A(\delay_line[1][13] ),
    .B(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__buf_1 _33124_ (.A(_05022_),
    .X(_05024_));
 sky130_fd_sc_hd__buf_1 _33125_ (.A(net447),
    .X(_05025_));
 sky130_fd_sc_hd__nand2_1 _33126_ (.A(_05024_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _33127_ (.A(_05023_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__nor2_1 _33128_ (.A(_01841_),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__and2_1 _33129_ (.A(_05027_),
    .B(_01841_),
    .X(_05029_));
 sky130_fd_sc_hd__nor3_2 _33130_ (.A(_05028_),
    .B(_03085_),
    .C(_05029_),
    .Y(_05031_));
 sky130_fd_sc_hd__o21a_1 _33131_ (.A1(_05029_),
    .A2(_05028_),
    .B1(_03085_),
    .X(_05032_));
 sky130_fd_sc_hd__o21ai_1 _33132_ (.A1(_03091_),
    .A2(_05025_),
    .B1(_00319_),
    .Y(_05033_));
 sky130_fd_sc_hd__or3_1 _33133_ (.A(_03091_),
    .B(_05025_),
    .C(_00319_),
    .X(_05034_));
 sky130_fd_sc_hd__o211a_1 _33134_ (.A1(_05031_),
    .A2(_05032_),
    .B1(_05033_),
    .C1(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__a211oi_2 _33135_ (.A1(_05033_),
    .A2(_05034_),
    .B1(_05031_),
    .C1(_05032_),
    .Y(_05036_));
 sky130_fd_sc_hd__nor3_1 _33136_ (.A(_05021_),
    .B(_05035_),
    .C(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__o21a_1 _33137_ (.A1(_05035_),
    .A2(_05036_),
    .B1(_05021_),
    .X(_05038_));
 sky130_fd_sc_hd__nor2_1 _33138_ (.A(_05037_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__xnor2_1 _33139_ (.A(_05020_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a21oi_1 _33140_ (.A1(_03497_),
    .A2(_03481_),
    .B1(_03495_),
    .Y(_05042_));
 sky130_fd_sc_hd__xnor2_1 _33141_ (.A(_05040_),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__xnor2_1 _33142_ (.A(_05018_),
    .B(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__a21oi_1 _33143_ (.A1(_01896_),
    .A2(_01899_),
    .B1(_03478_),
    .Y(_05045_));
 sky130_fd_sc_hd__a211o_1 _33144_ (.A1(_03479_),
    .A2(_03498_),
    .B1(_05044_),
    .C1(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__a21o_1 _33145_ (.A1(_03479_),
    .A2(_03498_),
    .B1(_05045_),
    .X(_05047_));
 sky130_fd_sc_hd__nand2_1 _33146_ (.A(_05044_),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__o21ai_1 _33147_ (.A1(_03078_),
    .A2(_03107_),
    .B1(_03104_),
    .Y(_05049_));
 sky130_fd_sc_hd__a21oi_1 _33148_ (.A1(_05046_),
    .A2(_05048_),
    .B1(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__and3_1 _33149_ (.A(_05049_),
    .B(_05046_),
    .C(_05048_),
    .X(_05051_));
 sky130_fd_sc_hd__nor2_2 _33150_ (.A(_05050_),
    .B(_05051_),
    .Y(_05053_));
 sky130_fd_sc_hd__or2_1 _33151_ (.A(_05017_),
    .B(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__nand2_4 _33152_ (.A(_05053_),
    .B(_05017_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_1 _33153_ (.A(_05054_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_1 _33154_ (.A(_03505_),
    .B(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__o31a_1 _33155_ (.A1(_01906_),
    .A2(_01938_),
    .A3(_01939_),
    .B1(_03507_),
    .X(_05058_));
 sky130_fd_sc_hd__o21a_1 _33156_ (.A1(_05058_),
    .A2(_03504_),
    .B1(_03505_),
    .X(_05059_));
 sky130_fd_sc_hd__nor2_2 _33157_ (.A(_05059_),
    .B(_05056_),
    .Y(_05060_));
 sky130_fd_sc_hd__o21bai_2 _33158_ (.A1(_03509_),
    .A2(_05057_),
    .B1_N(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__o21a_1 _33159_ (.A1(_03077_),
    .A2(_03114_),
    .B1(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__nor3_1 _33160_ (.A(_03077_),
    .B(_03114_),
    .C(_05061_),
    .Y(_05064_));
 sky130_fd_sc_hd__nor2_1 _33161_ (.A(_05062_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__o21ai_1 _33162_ (.A1(_05011_),
    .A2(_05016_),
    .B1(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__o21a_1 _33163_ (.A1(_03522_),
    .A2(_03520_),
    .B1(_03518_),
    .X(_05067_));
 sky130_fd_sc_hd__buf_2 _33164_ (.A(_05064_),
    .X(_05068_));
 sky130_fd_sc_hd__and3_1 _33165_ (.A(_04899_),
    .B(_04903_),
    .C(_05005_),
    .X(_05069_));
 sky130_fd_sc_hd__o21bai_1 _33166_ (.A1(_05006_),
    .A2(_05069_),
    .B1_N(_05015_),
    .Y(_05070_));
 sky130_fd_sc_hd__o221ai_1 _33167_ (.A1(_05062_),
    .A2(_05068_),
    .B1(_05006_),
    .B2(_05010_),
    .C1(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand3_1 _33168_ (.A(_05066_),
    .B(_05067_),
    .C(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__buf_2 _33169_ (.A(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__o21ai_2 _33170_ (.A1(_03522_),
    .A2(_03520_),
    .B1(_03518_),
    .Y(_05075_));
 sky130_fd_sc_hd__o22ai_2 _33171_ (.A1(_05062_),
    .A2(_05068_),
    .B1(_05011_),
    .B2(_05016_),
    .Y(_05076_));
 sky130_fd_sc_hd__o211ai_2 _33172_ (.A1(_05006_),
    .A2(_05010_),
    .B1(_05065_),
    .C1(_05070_),
    .Y(_05077_));
 sky130_fd_sc_hd__nand3_4 _33173_ (.A(_05075_),
    .B(_05076_),
    .C(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__a21bo_1 _33174_ (.A1(_03075_),
    .A2(_03119_),
    .B1_N(_03120_),
    .X(_05079_));
 sky130_fd_sc_hd__buf_2 _33175_ (.A(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__a21oi_4 _33176_ (.A1(_05073_),
    .A2(_05078_),
    .B1(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__nor2_1 _33177_ (.A(_03548_),
    .B(_03539_),
    .Y(_05082_));
 sky130_fd_sc_hd__nand3_2 _33178_ (.A(_05080_),
    .B(_05073_),
    .C(_05078_),
    .Y(_05083_));
 sky130_fd_sc_hd__o21ai_2 _33179_ (.A1(_03542_),
    .A2(_05082_),
    .B1(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__and3_1 _33180_ (.A(_05080_),
    .B(_05073_),
    .C(_05078_),
    .X(_05086_));
 sky130_fd_sc_hd__a21oi_1 _33181_ (.A1(_03548_),
    .A2(_03525_),
    .B1(_03538_),
    .Y(_05087_));
 sky130_fd_sc_hd__inv_2 _33182_ (.A(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__o21ai_4 _33183_ (.A1(_05081_),
    .A2(_05086_),
    .B1(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__o21ai_1 _33184_ (.A1(_05081_),
    .A2(_05084_),
    .B1(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__o21ai_2 _33185_ (.A1(_03552_),
    .A2(_04607_),
    .B1(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__a21o_1 _33186_ (.A1(_05072_),
    .A2(_05078_),
    .B1(_05079_),
    .X(_05092_));
 sky130_fd_sc_hd__o2111ai_4 _33187_ (.A1(_03531_),
    .A2(_03542_),
    .B1(_03529_),
    .C1(_05092_),
    .D1(_05083_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand4_4 _33188_ (.A(_03544_),
    .B(_03559_),
    .C(_05093_),
    .D(_05089_),
    .Y(_05094_));
 sky130_fd_sc_hd__buf_2 _33189_ (.A(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__nand2_1 _33190_ (.A(_05091_),
    .B(_05095_),
    .Y(_05097_));
 sky130_fd_sc_hd__nor2_1 _33191_ (.A(\delay_line[23][13] ),
    .B(\delay_line[23][14] ),
    .Y(_05098_));
 sky130_fd_sc_hd__nand2_2 _33192_ (.A(\delay_line[23][13] ),
    .B(\delay_line[23][14] ),
    .Y(_05099_));
 sky130_fd_sc_hd__and2b_1 _33193_ (.A_N(_05098_),
    .B(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__buf_2 _33194_ (.A(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__nand2_1 _33195_ (.A(_05097_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__nand3b_1 _33196_ (.A_N(_05101_),
    .B(_05091_),
    .C(_05095_),
    .Y(_05103_));
 sky130_fd_sc_hd__o21a_1 _33197_ (.A1(_03552_),
    .A2(_03559_),
    .B1(_03561_),
    .X(_05104_));
 sky130_fd_sc_hd__o21ba_1 _33198_ (.A1(_03067_),
    .A2(_05104_),
    .B1_N(_03068_),
    .X(_05105_));
 sky130_fd_sc_hd__a31oi_1 _33199_ (.A1(_04600_),
    .A2(_05102_),
    .A3(_05103_),
    .B1(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__clkbuf_2 _33200_ (.A(_05106_),
    .X(_05108_));
 sky130_fd_sc_hd__a21o_1 _33201_ (.A1(_05091_),
    .A2(_05095_),
    .B1(_05100_),
    .X(_05109_));
 sky130_fd_sc_hd__nand3_1 _33202_ (.A(_05091_),
    .B(_05095_),
    .C(_05101_),
    .Y(_05110_));
 sky130_fd_sc_hd__nand3b_1 _33203_ (.A_N(_04600_),
    .B(_05109_),
    .C(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__clkbuf_2 _33204_ (.A(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__inv_2 _33205_ (.A(_03680_),
    .Y(_05113_));
 sky130_fd_sc_hd__o21a_1 _33206_ (.A1(_03729_),
    .A2(_05113_),
    .B1(_03730_),
    .X(_05114_));
 sky130_fd_sc_hd__nand3_1 _33207_ (.A(_05102_),
    .B(_05103_),
    .C(_04600_),
    .Y(_05115_));
 sky130_fd_sc_hd__a21boi_1 _33208_ (.A1(_05112_),
    .A2(_05115_),
    .B1_N(_05105_),
    .Y(_05116_));
 sky130_fd_sc_hd__a211o_2 _33209_ (.A1(_05108_),
    .A2(_05112_),
    .B1(_05114_),
    .C1(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__nand2_1 _33210_ (.A(_05108_),
    .B(_05112_),
    .Y(_05119_));
 sky130_fd_sc_hd__nand2_1 _33211_ (.A(_05112_),
    .B(_05115_),
    .Y(_05120_));
 sky130_fd_sc_hd__nand2_1 _33212_ (.A(_05120_),
    .B(_05105_),
    .Y(_05121_));
 sky130_fd_sc_hd__a21bo_1 _33213_ (.A1(_05119_),
    .A2(_05121_),
    .B1_N(_05114_),
    .X(_05122_));
 sky130_fd_sc_hd__o211ai_4 _33214_ (.A1(_03573_),
    .A2(_04598_),
    .B1(_05117_),
    .C1(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__a211oi_2 _33215_ (.A1(_05108_),
    .A2(_05112_),
    .B1(_05114_),
    .C1(_05116_),
    .Y(_05124_));
 sky130_fd_sc_hd__a21boi_2 _33216_ (.A1(_05119_),
    .A2(_05121_),
    .B1_N(_05114_),
    .Y(_05125_));
 sky130_fd_sc_hd__a21oi_2 _33217_ (.A1(_03567_),
    .A2(_03563_),
    .B1(_03573_),
    .Y(_05126_));
 sky130_fd_sc_hd__o21ai_2 _33218_ (.A1(_05124_),
    .A2(_05125_),
    .B1(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__o211a_1 _33219_ (.A1(_03600_),
    .A2(_04597_),
    .B1(_05123_),
    .C1(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__o22ai_2 _33220_ (.A1(_03573_),
    .A2(_04598_),
    .B1(_05124_),
    .B2(_05125_),
    .Y(_05130_));
 sky130_fd_sc_hd__nand3_1 _33221_ (.A(_05122_),
    .B(_05126_),
    .C(_05117_),
    .Y(_05131_));
 sky130_fd_sc_hd__a21oi_1 _33222_ (.A1(_03582_),
    .A2(_03583_),
    .B1(_03600_),
    .Y(_05132_));
 sky130_fd_sc_hd__nand2_1 _33223_ (.A(_19848_),
    .B(_17897_),
    .Y(_05133_));
 sky130_fd_sc_hd__a2bb2o_1 _33224_ (.A1_N(_17901_),
    .A2_N(_17903_),
    .B1(_19848_),
    .B2(_22781_),
    .X(_05134_));
 sky130_fd_sc_hd__o21ai_1 _33225_ (.A1(_00435_),
    .A2(_05133_),
    .B1(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__or2_1 _33226_ (.A(_24241_),
    .B(_03564_),
    .X(_05136_));
 sky130_fd_sc_hd__nand2_1 _33227_ (.A(_24252_),
    .B(_03564_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand4_4 _33228_ (.A(_05136_),
    .B(_02016_),
    .C(_24251_),
    .D(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__a22o_1 _33229_ (.A1(_24251_),
    .A2(_02016_),
    .B1(_05137_),
    .B2(_05136_),
    .X(_05139_));
 sky130_fd_sc_hd__and3_1 _33230_ (.A(_05135_),
    .B(_05138_),
    .C(_05139_),
    .X(_05141_));
 sky130_fd_sc_hd__a21oi_1 _33231_ (.A1(_05138_),
    .A2(_05139_),
    .B1(_05135_),
    .Y(_05142_));
 sky130_fd_sc_hd__nor2_1 _33232_ (.A(_05141_),
    .B(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__a31o_1 _33233_ (.A1(_05130_),
    .A2(_05131_),
    .A3(_05132_),
    .B1(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__o211ai_4 _33234_ (.A1(_03600_),
    .A2(_04597_),
    .B1(_05123_),
    .C1(_05127_),
    .Y(_05145_));
 sky130_fd_sc_hd__nand3_1 _33235_ (.A(_05130_),
    .B(_05131_),
    .C(_05132_),
    .Y(_05146_));
 sky130_fd_sc_hd__inv_2 _33236_ (.A(_05143_),
    .Y(_05147_));
 sky130_fd_sc_hd__a21o_1 _33237_ (.A1(_05145_),
    .A2(_05146_),
    .B1(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__o221ai_2 _33238_ (.A1(_03866_),
    .A2(_03868_),
    .B1(_05128_),
    .B2(_05144_),
    .C1(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__o2bb2ai_1 _33239_ (.A1_N(_05145_),
    .A2_N(_05146_),
    .B1(_05141_),
    .B2(_05142_),
    .Y(_05150_));
 sky130_fd_sc_hd__nand3_1 _33240_ (.A(_05145_),
    .B(_05146_),
    .C(_05143_),
    .Y(_05151_));
 sky130_fd_sc_hd__a21oi_2 _33241_ (.A1(_03620_),
    .A2(_03864_),
    .B1(_03866_),
    .Y(_05152_));
 sky130_fd_sc_hd__nand3_2 _33242_ (.A(_05150_),
    .B(_05151_),
    .C(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__a21oi_1 _33243_ (.A1(_03588_),
    .A2(_03597_),
    .B1(_03603_),
    .Y(_05154_));
 sky130_fd_sc_hd__a21bo_1 _33244_ (.A1(_05149_),
    .A2(_05153_),
    .B1_N(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__and2_1 _33245_ (.A(_03588_),
    .B(_03597_),
    .X(_05156_));
 sky130_fd_sc_hd__clkbuf_2 _33246_ (.A(_05149_),
    .X(_05157_));
 sky130_fd_sc_hd__o211ai_2 _33247_ (.A1(_03603_),
    .A2(_05156_),
    .B1(_05157_),
    .C1(_05153_),
    .Y(_05158_));
 sky130_fd_sc_hd__a21oi_1 _33248_ (.A1(_04433_),
    .A2(_04435_),
    .B1(_04432_),
    .Y(_05159_));
 sky130_fd_sc_hd__buf_1 _33249_ (.A(_03735_),
    .X(_05160_));
 sky130_fd_sc_hd__and3_1 _33250_ (.A(_21087_),
    .B(_02880_),
    .C(_05160_),
    .X(_05162_));
 sky130_fd_sc_hd__a21oi_1 _33251_ (.A1(_02880_),
    .A2(_05160_),
    .B1(_21087_),
    .Y(_05163_));
 sky130_fd_sc_hd__or2_1 _33252_ (.A(_03735_),
    .B(_01079_),
    .X(_05164_));
 sky130_fd_sc_hd__nand2_1 _33253_ (.A(_03735_),
    .B(_01079_),
    .Y(_05165_));
 sky130_fd_sc_hd__and2b_1 _33254_ (.A_N(net305),
    .B(net304),
    .X(_05166_));
 sky130_fd_sc_hd__and2b_1 _33255_ (.A_N(net304),
    .B(net305),
    .X(_05167_));
 sky130_fd_sc_hd__o21ai_1 _33256_ (.A1(_05166_),
    .A2(_05167_),
    .B1(_03739_),
    .Y(_05168_));
 sky130_fd_sc_hd__or3_1 _33257_ (.A(_03739_),
    .B(_05166_),
    .C(_05167_),
    .X(_05169_));
 sky130_fd_sc_hd__a22oi_1 _33258_ (.A1(_05164_),
    .A2(_05165_),
    .B1(_05168_),
    .B2(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__and4_1 _33259_ (.A(_05164_),
    .B(_05165_),
    .C(_05168_),
    .D(_05169_),
    .X(_05171_));
 sky130_fd_sc_hd__a211o_1 _33260_ (.A1(_03740_),
    .A2(_03743_),
    .B1(_05170_),
    .C1(_05171_),
    .X(_05173_));
 sky130_fd_sc_hd__inv_2 _33261_ (.A(_05173_),
    .Y(_05174_));
 sky130_fd_sc_hd__o211a_1 _33262_ (.A1(_05170_),
    .A2(_05171_),
    .B1(_03740_),
    .C1(_03743_),
    .X(_05175_));
 sky130_fd_sc_hd__or4_2 _33263_ (.A(_05162_),
    .B(_05163_),
    .C(_05174_),
    .D(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__or2_1 _33264_ (.A(_05162_),
    .B(_05163_),
    .X(_05177_));
 sky130_fd_sc_hd__o21ai_1 _33265_ (.A1(_05174_),
    .A2(_05175_),
    .B1(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__a221o_1 _33266_ (.A1(_03749_),
    .A2(_03746_),
    .B1(_05176_),
    .B2(_05178_),
    .C1(_03747_),
    .X(_05179_));
 sky130_fd_sc_hd__and3_1 _33267_ (.A(_03748_),
    .B(_03749_),
    .C(_03746_),
    .X(_05180_));
 sky130_fd_sc_hd__o211ai_2 _33268_ (.A1(_03747_),
    .A2(_05180_),
    .B1(_05176_),
    .C1(_05178_),
    .Y(_05181_));
 sky130_fd_sc_hd__or4bb_2 _33269_ (.A(_24876_),
    .B(_02882_),
    .C_N(_05179_),
    .D_N(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__a2bb2o_1 _33270_ (.A1_N(_02882_),
    .A2_N(_24876_),
    .B1(_05181_),
    .B2(_05179_),
    .X(_05184_));
 sky130_fd_sc_hd__a221o_1 _33271_ (.A1(_02879_),
    .A2(_03756_),
    .B1(_05182_),
    .B2(_05184_),
    .C1(_03754_),
    .X(_05185_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33272_ (.A(_01072_),
    .X(_05186_));
 sky130_fd_sc_hd__and4b_1 _33273_ (.A_N(_24873_),
    .B(_01075_),
    .C(_05186_),
    .D(_03756_),
    .X(_05187_));
 sky130_fd_sc_hd__o211ai_4 _33274_ (.A1(_03754_),
    .A2(_05187_),
    .B1(_05182_),
    .C1(_05184_),
    .Y(_05188_));
 sky130_fd_sc_hd__o211a_1 _33275_ (.A1(_03759_),
    .A2(_03763_),
    .B1(_05185_),
    .C1(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__a211oi_1 _33276_ (.A1(_05185_),
    .A2(_05188_),
    .B1(_03759_),
    .C1(_03763_),
    .Y(_05190_));
 sky130_fd_sc_hd__or2_1 _33277_ (.A(_05189_),
    .B(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__a31o_1 _33278_ (.A1(_02826_),
    .A2(_02817_),
    .A3(_03837_),
    .B1(_03836_),
    .X(_05192_));
 sky130_fd_sc_hd__nor2_1 _33279_ (.A(_03823_),
    .B(_03831_),
    .Y(_05193_));
 sky130_fd_sc_hd__nor2_1 _33280_ (.A(\delay_line[32][13] ),
    .B(\delay_line[32][14] ),
    .Y(_05195_));
 sky130_fd_sc_hd__buf_1 _33281_ (.A(\delay_line[32][14] ),
    .X(_05196_));
 sky130_fd_sc_hd__nand2_1 _33282_ (.A(_03811_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__nand3b_1 _33283_ (.A_N(_05195_),
    .B(_05197_),
    .C(_02793_),
    .Y(_05198_));
 sky130_fd_sc_hd__and2_1 _33284_ (.A(\delay_line[32][13] ),
    .B(\delay_line[32][14] ),
    .X(_05199_));
 sky130_fd_sc_hd__o21bai_1 _33285_ (.A1(_05195_),
    .A2(_05199_),
    .B1_N(_02793_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand2_1 _33286_ (.A(_05198_),
    .B(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__a21o_1 _33287_ (.A1(_03815_),
    .A2(_03813_),
    .B1(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__nor2_1 _33288_ (.A(_03809_),
    .B(_03812_),
    .Y(_05203_));
 sky130_fd_sc_hd__inv_2 _33289_ (.A(_01113_),
    .Y(_05204_));
 sky130_fd_sc_hd__o211ai_2 _33290_ (.A1(_05203_),
    .A2(_05204_),
    .B1(_03815_),
    .C1(_05201_),
    .Y(_05206_));
 sky130_fd_sc_hd__clkbuf_2 _33291_ (.A(_01113_),
    .X(_05207_));
 sky130_fd_sc_hd__a21oi_2 _33292_ (.A1(_05202_),
    .A2(_05206_),
    .B1(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__and3_1 _33293_ (.A(_05202_),
    .B(_05206_),
    .C(_05207_),
    .X(_05209_));
 sky130_fd_sc_hd__a211oi_4 _33294_ (.A1(_03818_),
    .A2(_03820_),
    .B1(_05208_),
    .C1(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__clkbuf_2 _33295_ (.A(_01121_),
    .X(_05211_));
 sky130_fd_sc_hd__nor2_1 _33296_ (.A(_03826_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand2_1 _33297_ (.A(_05211_),
    .B(_03826_),
    .Y(_05213_));
 sky130_fd_sc_hd__or4b_2 _33298_ (.A(_01132_),
    .B(_24969_),
    .C(_05212_),
    .D_N(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__nand2_1 _33299_ (.A(_21112_),
    .B(_21116_),
    .Y(_05215_));
 sky130_fd_sc_hd__a2bb2o_1 _33300_ (.A1_N(_01132_),
    .A2_N(_24969_),
    .B1(_05215_),
    .B2(_05213_),
    .X(_05217_));
 sky130_fd_sc_hd__nand2_1 _33301_ (.A(_05214_),
    .B(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__o211ai_1 _33302_ (.A1(_05208_),
    .A2(_05209_),
    .B1(_03818_),
    .C1(_03820_),
    .Y(_05219_));
 sky130_fd_sc_hd__inv_2 _33303_ (.A(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__nor3_1 _33304_ (.A(_05210_),
    .B(_05218_),
    .C(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__o21ai_1 _33305_ (.A1(_05220_),
    .A2(_05210_),
    .B1(_05218_),
    .Y(_05222_));
 sky130_fd_sc_hd__and2b_1 _33306_ (.A_N(_05221_),
    .B(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__xnor2_2 _33307_ (.A(_05193_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__xnor2_2 _33308_ (.A(_03827_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__nor2_1 _33309_ (.A(_05192_),
    .B(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__o21a_1 _33310_ (.A1(_03836_),
    .A2(_03839_),
    .B1(_05225_),
    .X(_05228_));
 sky130_fd_sc_hd__nor2_1 _33311_ (.A(_05226_),
    .B(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__xnor2_2 _33312_ (.A(_03844_),
    .B(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__inv_2 _33313_ (.A(_03808_),
    .Y(_05231_));
 sky130_fd_sc_hd__o21bai_1 _33314_ (.A1(_01153_),
    .A2(_01155_),
    .B1_N(_02790_),
    .Y(_05232_));
 sky130_fd_sc_hd__a21oi_2 _33315_ (.A1(_05232_),
    .A2(_02831_),
    .B1(_03806_),
    .Y(_05233_));
 sky130_fd_sc_hd__o22ai_4 _33316_ (.A1(_05231_),
    .A2(_03840_),
    .B1(_03845_),
    .B2(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__xnor2_2 _33317_ (.A(_05230_),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__a21oi_1 _33318_ (.A1(_01160_),
    .A2(_02839_),
    .B1(_03781_),
    .Y(_05236_));
 sky130_fd_sc_hd__clkbuf_2 _33319_ (.A(_02840_),
    .X(_05237_));
 sky130_fd_sc_hd__and3_1 _33320_ (.A(_01160_),
    .B(_03769_),
    .C(_05237_),
    .X(_05239_));
 sky130_fd_sc_hd__nor3_1 _33321_ (.A(_03778_),
    .B(_03784_),
    .C(_03785_),
    .Y(_05240_));
 sky130_fd_sc_hd__inv_2 _33322_ (.A(\delay_line[33][10] ),
    .Y(_05241_));
 sky130_fd_sc_hd__buf_1 _33323_ (.A(\delay_line[33][9] ),
    .X(_05242_));
 sky130_fd_sc_hd__and2_1 _33324_ (.A(_05241_),
    .B(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__nor2_1 _33325_ (.A(_05242_),
    .B(_05241_),
    .Y(_05244_));
 sky130_fd_sc_hd__nor3_1 _33326_ (.A(net310),
    .B(_05243_),
    .C(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__o21a_1 _33327_ (.A1(_05243_),
    .A2(_05244_),
    .B1(net310),
    .X(_05246_));
 sky130_fd_sc_hd__o21a_1 _33328_ (.A1(_05245_),
    .A2(_05246_),
    .B1(_03775_),
    .X(_05247_));
 sky130_fd_sc_hd__inv_2 _33329_ (.A(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__or3_1 _33330_ (.A(_03775_),
    .B(_05245_),
    .C(_05246_),
    .X(_05250_));
 sky130_fd_sc_hd__nand2_1 _33331_ (.A(_18651_),
    .B(_03769_),
    .Y(_05251_));
 sky130_fd_sc_hd__buf_1 _33332_ (.A(_05242_),
    .X(_05252_));
 sky130_fd_sc_hd__o21ai_1 _33333_ (.A1(_05252_),
    .A2(_23357_),
    .B1(_03780_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand3b_1 _33334_ (.A_N(_05252_),
    .B(_02840_),
    .C(_02836_),
    .Y(_05254_));
 sky130_fd_sc_hd__and2_1 _33335_ (.A(_05253_),
    .B(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__xnor2_1 _33336_ (.A(_05251_),
    .B(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__a21o_1 _33337_ (.A1(_05248_),
    .A2(_05250_),
    .B1(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__nand3_1 _33338_ (.A(_05256_),
    .B(_05248_),
    .C(_05250_),
    .Y(_05258_));
 sky130_fd_sc_hd__or4bb_1 _33339_ (.A(_03778_),
    .B(_05240_),
    .C_N(_05257_),
    .D_N(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__a2bb2o_1 _33340_ (.A1_N(_03778_),
    .A2_N(_05240_),
    .B1(_05257_),
    .B2(_05258_),
    .X(_05261_));
 sky130_fd_sc_hd__o211a_1 _33341_ (.A1(_05236_),
    .A2(_05239_),
    .B1(_05259_),
    .C1(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__a211oi_1 _33342_ (.A1(_05259_),
    .A2(_05261_),
    .B1(_05236_),
    .C1(_05239_),
    .Y(_05263_));
 sky130_fd_sc_hd__a211oi_1 _33343_ (.A1(_03790_),
    .A2(_03791_),
    .B1(_05262_),
    .C1(_05263_),
    .Y(_05264_));
 sky130_fd_sc_hd__o211ai_1 _33344_ (.A1(_05262_),
    .A2(_05263_),
    .B1(_03790_),
    .C1(_03791_),
    .Y(_05265_));
 sky130_fd_sc_hd__or4b_1 _33345_ (.A(_03767_),
    .B(_03793_),
    .C(_05264_),
    .D_N(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__inv_2 _33346_ (.A(_05264_),
    .Y(_05267_));
 sky130_fd_sc_hd__a2bb2o_1 _33347_ (.A1_N(_03793_),
    .A2_N(_03767_),
    .B1(_05265_),
    .B2(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__nand2_1 _33348_ (.A(_05266_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__a21oi_2 _33349_ (.A1(_03798_),
    .A2(_03797_),
    .B1(_03795_),
    .Y(_05270_));
 sky130_fd_sc_hd__xnor2_2 _33350_ (.A(_05269_),
    .B(_05270_),
    .Y(_05272_));
 sky130_fd_sc_hd__xor2_1 _33351_ (.A(_05235_),
    .B(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__xor2_1 _33352_ (.A(_05191_),
    .B(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__a21o_1 _33353_ (.A1(_04423_),
    .A2(_04427_),
    .B1(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__a21boi_1 _33354_ (.A1(_03800_),
    .A2(_03847_),
    .B1_N(_03849_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand3_1 _33355_ (.A(_04423_),
    .B(_04427_),
    .C(_05274_),
    .Y(_05277_));
 sky130_fd_sc_hd__and3_1 _33356_ (.A(_05275_),
    .B(_05276_),
    .C(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__a21oi_1 _33357_ (.A1(_05277_),
    .A2(_05275_),
    .B1(_05276_),
    .Y(_05279_));
 sky130_fd_sc_hd__o22a_1 _33358_ (.A1(_03853_),
    .A2(_03857_),
    .B1(_05278_),
    .B2(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__nor4_1 _33359_ (.A(_03853_),
    .B(_03857_),
    .C(_05278_),
    .D(_05279_),
    .Y(_05281_));
 sky130_fd_sc_hd__inv_2 _33360_ (.A(_03726_),
    .Y(_05283_));
 sky130_fd_sc_hd__buf_1 _33361_ (.A(\delay_line[37][13] ),
    .X(_05284_));
 sky130_fd_sc_hd__or2b_1 _33362_ (.A(_02732_),
    .B_N(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__or3b_1 _33363_ (.A(_01269_),
    .B(_03682_),
    .C_N(_03681_),
    .X(_05286_));
 sky130_fd_sc_hd__xnor2_1 _33364_ (.A(\delay_line[37][12] ),
    .B(\delay_line[37][14] ),
    .Y(_05287_));
 sky130_fd_sc_hd__and3_1 _33365_ (.A(_05285_),
    .B(_05286_),
    .C(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__a21oi_1 _33366_ (.A1(_05285_),
    .A2(_05286_),
    .B1(_05287_),
    .Y(_05289_));
 sky130_fd_sc_hd__nor2_1 _33367_ (.A(_05288_),
    .B(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__inv_2 _33368_ (.A(_03685_),
    .Y(_05291_));
 sky130_fd_sc_hd__o2bb2a_1 _33369_ (.A1_N(_05284_),
    .A2_N(_03683_),
    .B1(_05291_),
    .B2(_03686_),
    .X(_05292_));
 sky130_fd_sc_hd__xnor2_2 _33370_ (.A(_05290_),
    .B(_05292_),
    .Y(_05294_));
 sky130_fd_sc_hd__buf_1 _33371_ (.A(\delay_line[36][10] ),
    .X(_05295_));
 sky130_fd_sc_hd__nand2_1 _33372_ (.A(_05295_),
    .B(_03691_),
    .Y(_05296_));
 sky130_fd_sc_hd__and2b_1 _33373_ (.A_N(_02764_),
    .B(_05295_),
    .X(_05297_));
 sky130_fd_sc_hd__nor2b_1 _33374_ (.A(net296),
    .B_N(\delay_line[36][11] ),
    .Y(_05298_));
 sky130_fd_sc_hd__and2b_1 _33375_ (.A_N(\delay_line[36][11] ),
    .B(net296),
    .X(_05299_));
 sky130_fd_sc_hd__nor2_1 _33376_ (.A(_05298_),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__a211oi_1 _33377_ (.A1(_03690_),
    .A2(_03692_),
    .B1(_05297_),
    .C1(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__and3_1 _33378_ (.A(_03688_),
    .B(_03690_),
    .C(_03692_),
    .X(_05302_));
 sky130_fd_sc_hd__o21a_1 _33379_ (.A1(_05297_),
    .A2(_05302_),
    .B1(_05300_),
    .X(_05303_));
 sky130_fd_sc_hd__a211oi_2 _33380_ (.A1(_03698_),
    .A2(_05296_),
    .B1(_05301_),
    .C1(_05303_),
    .Y(_05305_));
 sky130_fd_sc_hd__nor2_1 _33381_ (.A(_03693_),
    .B(_03695_),
    .Y(_05306_));
 sky130_fd_sc_hd__nand2_1 _33382_ (.A(_01288_),
    .B(_02765_),
    .Y(_05307_));
 sky130_fd_sc_hd__nor2_1 _33383_ (.A(_02773_),
    .B(_02771_),
    .Y(_05308_));
 sky130_fd_sc_hd__a21oi_1 _33384_ (.A1(_05307_),
    .A2(_05308_),
    .B1(_03696_),
    .Y(_05309_));
 sky130_fd_sc_hd__o221a_1 _33385_ (.A1(_05306_),
    .A2(_05309_),
    .B1(_05303_),
    .B2(_05301_),
    .C1(_05296_),
    .X(_05310_));
 sky130_fd_sc_hd__nor2_1 _33386_ (.A(_05305_),
    .B(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__nor3b_1 _33387_ (.A(_03704_),
    .B(_03705_),
    .C_N(_03702_),
    .Y(_05312_));
 sky130_fd_sc_hd__nor2_1 _33388_ (.A(net300),
    .B(net299),
    .Y(_05313_));
 sky130_fd_sc_hd__and2_1 _33389_ (.A(net300),
    .B(net299),
    .X(_05314_));
 sky130_fd_sc_hd__or3b_1 _33390_ (.A(_05313_),
    .B(_05314_),
    .C_N(_03703_),
    .X(_05316_));
 sky130_fd_sc_hd__o21bai_1 _33391_ (.A1(_05313_),
    .A2(_05314_),
    .B1_N(_03703_),
    .Y(_05317_));
 sky130_fd_sc_hd__o211a_1 _33392_ (.A1(_03704_),
    .A2(_05312_),
    .B1(_05316_),
    .C1(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__buf_1 _33393_ (.A(_03703_),
    .X(_05319_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33394_ (.A(net300),
    .X(_05320_));
 sky130_fd_sc_hd__a221oi_2 _33395_ (.A1(_05319_),
    .A2(_05320_),
    .B1(_05316_),
    .B2(_05317_),
    .C1(_05312_),
    .Y(_05321_));
 sky130_fd_sc_hd__nor3_1 _33396_ (.A(_03710_),
    .B(_05318_),
    .C(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__o21ai_1 _33397_ (.A1(_05318_),
    .A2(_05321_),
    .B1(_03710_),
    .Y(_05323_));
 sky130_fd_sc_hd__inv_2 _33398_ (.A(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__nor3_1 _33399_ (.A(_23503_),
    .B(_05322_),
    .C(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__o21a_1 _33400_ (.A1(_05322_),
    .A2(_05324_),
    .B1(_23503_),
    .X(_05327_));
 sky130_fd_sc_hd__a211oi_2 _33401_ (.A1(_03712_),
    .A2(_03715_),
    .B1(net201),
    .C1(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hd__o221a_1 _33402_ (.A1(_20842_),
    .A2(_03714_),
    .B1(net201),
    .B2(_05327_),
    .C1(_03712_),
    .X(_05329_));
 sky130_fd_sc_hd__inv_2 _33403_ (.A(_03719_),
    .Y(_05330_));
 sky130_fd_sc_hd__a21oi_1 _33404_ (.A1(_03720_),
    .A2(_05330_),
    .B1(_03717_),
    .Y(_05331_));
 sky130_fd_sc_hd__o21ai_1 _33405_ (.A1(_05328_),
    .A2(_05329_),
    .B1(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__or3_1 _33406_ (.A(_05328_),
    .B(_05329_),
    .C(_05331_),
    .X(_05333_));
 sky130_fd_sc_hd__nand2_1 _33407_ (.A(_05332_),
    .B(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__xor2_2 _33408_ (.A(_05311_),
    .B(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__xnor2_2 _33409_ (.A(_05294_),
    .B(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__and3_1 _33410_ (.A(_03724_),
    .B(_05283_),
    .C(_05336_),
    .X(_05338_));
 sky130_fd_sc_hd__a21oi_4 _33411_ (.A1(_03724_),
    .A2(_05283_),
    .B1(_05336_),
    .Y(_05339_));
 sky130_fd_sc_hd__nor2_1 _33412_ (.A(_05338_),
    .B(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33413_ (.A(\delay_line[40][13] ),
    .X(_05341_));
 sky130_fd_sc_hd__buf_2 _33414_ (.A(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__nor2_1 _33415_ (.A(_05342_),
    .B(_02718_),
    .Y(_05343_));
 sky130_fd_sc_hd__and2_1 _33416_ (.A(\delay_line[40][13] ),
    .B(\delay_line[40][14] ),
    .X(_05344_));
 sky130_fd_sc_hd__nor2_1 _33417_ (.A(_05341_),
    .B(\delay_line[40][14] ),
    .Y(_05345_));
 sky130_fd_sc_hd__a2bb2o_1 _33418_ (.A1_N(_05344_),
    .A2_N(_05345_),
    .B1(_03662_),
    .B2(_05341_),
    .X(_05346_));
 sky130_fd_sc_hd__nand3b_2 _33419_ (.A_N(\delay_line[40][14] ),
    .B(_05341_),
    .C(_03662_),
    .Y(_05347_));
 sky130_fd_sc_hd__a21bo_1 _33420_ (.A1(_05346_),
    .A2(_05347_),
    .B1_N(_03658_),
    .X(_05349_));
 sky130_fd_sc_hd__nand3b_1 _33421_ (.A_N(_03658_),
    .B(_05346_),
    .C(_05347_),
    .Y(_05350_));
 sky130_fd_sc_hd__and4bb_1 _33422_ (.A_N(_05343_),
    .B_N(_03670_),
    .C(_05349_),
    .D(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__a2bb2oi_1 _33423_ (.A1_N(_05343_),
    .A2_N(_03670_),
    .B1(_05349_),
    .B2(_05350_),
    .Y(_05352_));
 sky130_fd_sc_hd__o221ai_1 _33424_ (.A1(_03660_),
    .A2(_03662_),
    .B1(_03669_),
    .B2(_03670_),
    .C1(_03671_),
    .Y(_05353_));
 sky130_fd_sc_hd__a21oi_1 _33425_ (.A1(_05353_),
    .A2(_03675_),
    .B1(_03674_),
    .Y(_05354_));
 sky130_fd_sc_hd__or3_1 _33426_ (.A(_05351_),
    .B(_05352_),
    .C(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__o21ai_1 _33427_ (.A1(_05351_),
    .A2(_05352_),
    .B1(_05354_),
    .Y(_05356_));
 sky130_fd_sc_hd__nand2_1 _33428_ (.A(_05355_),
    .B(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__buf_1 _33429_ (.A(_03624_),
    .X(_05358_));
 sky130_fd_sc_hd__buf_1 _33430_ (.A(\delay_line[39][13] ),
    .X(_05360_));
 sky130_fd_sc_hd__o21ai_1 _33431_ (.A1(_05358_),
    .A2(_05360_),
    .B1(_03622_),
    .Y(_05361_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33432_ (.A(\delay_line[39][14] ),
    .X(_05362_));
 sky130_fd_sc_hd__nand2b_1 _33433_ (.A_N(_05362_),
    .B(_05360_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2b_1 _33434_ (.A_N(_05360_),
    .B(\delay_line[39][14] ),
    .Y(_05364_));
 sky130_fd_sc_hd__and3b_1 _33435_ (.A_N(_03624_),
    .B(_05363_),
    .C(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__a21boi_1 _33436_ (.A1(_05363_),
    .A2(_05364_),
    .B1_N(_03624_),
    .Y(_05366_));
 sky130_fd_sc_hd__or2_1 _33437_ (.A(_05365_),
    .B(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__a21oi_1 _33438_ (.A1(_03627_),
    .A2(_05361_),
    .B1(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__and3_1 _33439_ (.A(_03627_),
    .B(_05361_),
    .C(_05367_),
    .X(_05369_));
 sky130_fd_sc_hd__or3b_1 _33440_ (.A(_05368_),
    .B(_05369_),
    .C_N(_03622_),
    .X(_05371_));
 sky130_fd_sc_hd__o21bai_1 _33441_ (.A1(_05368_),
    .A2(_05369_),
    .B1_N(_03622_),
    .Y(_05372_));
 sky130_fd_sc_hd__a221o_1 _33442_ (.A1(_02693_),
    .A2(_03632_),
    .B1(_05371_),
    .B2(_05372_),
    .C1(_03630_),
    .X(_05373_));
 sky130_fd_sc_hd__a21o_1 _33443_ (.A1(_03631_),
    .A2(_02693_),
    .B1(_03630_),
    .X(_05374_));
 sky130_fd_sc_hd__nand3_2 _33444_ (.A(_05374_),
    .B(_05371_),
    .C(_05372_),
    .Y(_05375_));
 sky130_fd_sc_hd__a211o_1 _33445_ (.A1(_05373_),
    .A2(_05375_),
    .B1(_03636_),
    .C1(_03639_),
    .X(_05376_));
 sky130_fd_sc_hd__o211a_1 _33446_ (.A1(_03636_),
    .A2(_03639_),
    .B1(_05373_),
    .C1(_05375_),
    .X(_05377_));
 sky130_fd_sc_hd__inv_2 _33447_ (.A(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__buf_1 _33448_ (.A(\delay_line[38][14] ),
    .X(_05379_));
 sky130_fd_sc_hd__nor2_1 _33449_ (.A(_03642_),
    .B(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__and2_1 _33450_ (.A(_03642_),
    .B(\delay_line[38][14] ),
    .X(_05382_));
 sky130_fd_sc_hd__buf_1 _33451_ (.A(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__a2111oi_1 _33452_ (.A1(_02684_),
    .A2(_03646_),
    .B1(_05380_),
    .C1(_05383_),
    .D1(_03644_),
    .Y(_05384_));
 sky130_fd_sc_hd__and3_1 _33453_ (.A(_01223_),
    .B(net285),
    .C(_03646_),
    .X(_05385_));
 sky130_fd_sc_hd__o22a_1 _33454_ (.A1(_05380_),
    .A2(_05383_),
    .B1(_05385_),
    .B2(_03644_),
    .X(_05386_));
 sky130_fd_sc_hd__a31o_1 _33455_ (.A1(_01220_),
    .A2(_03641_),
    .A3(_03646_),
    .B1(_03652_),
    .X(_05387_));
 sky130_fd_sc_hd__or3_1 _33456_ (.A(net269),
    .B(_05386_),
    .C(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__o21ai_1 _33457_ (.A1(net268),
    .A2(_05386_),
    .B1(_05387_),
    .Y(_05389_));
 sky130_fd_sc_hd__and2_1 _33458_ (.A(_05388_),
    .B(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__a21oi_2 _33459_ (.A1(_05376_),
    .A2(_05378_),
    .B1(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__and3_1 _33460_ (.A(_05378_),
    .B(_05390_),
    .C(_05376_),
    .X(_05393_));
 sky130_fd_sc_hd__or3_1 _33461_ (.A(_05357_),
    .B(_05391_),
    .C(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__o21ai_1 _33462_ (.A1(_05393_),
    .A2(_05391_),
    .B1(_05357_),
    .Y(_05395_));
 sky130_fd_sc_hd__and2_2 _33463_ (.A(_05394_),
    .B(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__and2_1 _33464_ (.A(_05340_),
    .B(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__nor2_1 _33465_ (.A(_05340_),
    .B(_05396_),
    .Y(_05398_));
 sky130_fd_sc_hd__or2_2 _33466_ (.A(_05397_),
    .B(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__o21a_1 _33467_ (.A1(_05280_),
    .A2(net83),
    .B1(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__nor3_1 _33468_ (.A(_05280_),
    .B(net83),
    .C(_05399_),
    .Y(_05401_));
 sky130_fd_sc_hd__nor2_1 _33469_ (.A(_05400_),
    .B(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__xor2_1 _33470_ (.A(_05159_),
    .B(_05402_),
    .X(_05404_));
 sky130_fd_sc_hd__o311a_1 _33471_ (.A1(_03734_),
    .A2(_03855_),
    .A3(_03857_),
    .B1(_03862_),
    .C1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__a21o_1 _33472_ (.A1(_03858_),
    .A2(_03862_),
    .B1(_05404_),
    .X(_05406_));
 sky130_fd_sc_hd__inv_2 _33473_ (.A(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__and4_1 _33474_ (.A(_06271_),
    .B(_02142_),
    .C(_02143_),
    .D(_02145_),
    .X(_05408_));
 sky130_fd_sc_hd__buf_1 _33475_ (.A(\delay_line[31][14] ),
    .X(_05409_));
 sky130_fd_sc_hd__or2b_1 _33476_ (.A(_05409_),
    .B_N(_02127_),
    .X(_05410_));
 sky130_fd_sc_hd__or2b_1 _33477_ (.A(\delay_line[31][12] ),
    .B_N(\delay_line[31][14] ),
    .X(_05411_));
 sky130_fd_sc_hd__a21o_1 _33478_ (.A1(_05410_),
    .A2(_05411_),
    .B1(\delay_line[31][13] ),
    .X(_05412_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33479_ (.A(_05411_),
    .X(_05413_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33480_ (.A(\delay_line[31][13] ),
    .X(_05415_));
 sky130_fd_sc_hd__nand3_1 _33481_ (.A(_05410_),
    .B(_05413_),
    .C(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__a21oi_1 _33482_ (.A1(_04351_),
    .A2(_05415_),
    .B1(_00885_),
    .Y(_05417_));
 sky130_fd_sc_hd__a211oi_1 _33483_ (.A1(_05412_),
    .A2(_05416_),
    .B1(_04352_),
    .C1(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__inv_2 _33484_ (.A(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__o211ai_1 _33485_ (.A1(_04352_),
    .A2(_05417_),
    .B1(_05412_),
    .C1(_05416_),
    .Y(_05420_));
 sky130_fd_sc_hd__a21boi_1 _33486_ (.A1(_05419_),
    .A2(_05420_),
    .B1_N(_04357_),
    .Y(_05421_));
 sky130_fd_sc_hd__or2_1 _33487_ (.A(_21270_),
    .B(_21262_),
    .X(_05422_));
 sky130_fd_sc_hd__buf_1 _33488_ (.A(_21262_),
    .X(_05423_));
 sky130_fd_sc_hd__nand2_1 _33489_ (.A(_05423_),
    .B(_02144_),
    .Y(_05424_));
 sky130_fd_sc_hd__and3_1 _33490_ (.A(_05422_),
    .B(_05424_),
    .C(_04346_),
    .X(_05426_));
 sky130_fd_sc_hd__o2bb2a_1 _33491_ (.A1_N(_05422_),
    .A2_N(_05424_),
    .B1(_02143_),
    .B2(_23212_),
    .X(_05427_));
 sky130_fd_sc_hd__or2_1 _33492_ (.A(_05426_),
    .B(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__nand3b_1 _33493_ (.A_N(_04357_),
    .B(_05419_),
    .C(_05420_),
    .Y(_05429_));
 sky130_fd_sc_hd__inv_2 _33494_ (.A(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__nor3_2 _33495_ (.A(_05421_),
    .B(_05428_),
    .C(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__o22a_1 _33496_ (.A1(_05426_),
    .A2(_05427_),
    .B1(_05430_),
    .B2(_05421_),
    .X(_05432_));
 sky130_fd_sc_hd__a211oi_1 _33497_ (.A1(_04359_),
    .A2(_04362_),
    .B1(_05431_),
    .C1(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__o211a_1 _33498_ (.A1(_05431_),
    .A2(_05432_),
    .B1(_04359_),
    .C1(_04362_),
    .X(_05434_));
 sky130_fd_sc_hd__or3_1 _33499_ (.A(_04348_),
    .B(_05433_),
    .C(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__o21ai_1 _33500_ (.A1(_05433_),
    .A2(_05434_),
    .B1(_04348_),
    .Y(_05437_));
 sky130_fd_sc_hd__a221o_1 _33501_ (.A1(_05408_),
    .A2(_04367_),
    .B1(_05435_),
    .B2(_05437_),
    .C1(_04365_),
    .X(_05438_));
 sky130_fd_sc_hd__o211ai_1 _33502_ (.A1(_04365_),
    .A2(_04368_),
    .B1(_05435_),
    .C1(_05437_),
    .Y(_05439_));
 sky130_fd_sc_hd__and4_1 _33503_ (.A(_04345_),
    .B(_05438_),
    .C(_05439_),
    .D(_04370_),
    .X(_05440_));
 sky130_fd_sc_hd__a22oi_1 _33504_ (.A1(_04345_),
    .A2(_04370_),
    .B1(_05438_),
    .B2(_05439_),
    .Y(_05441_));
 sky130_fd_sc_hd__or2_2 _33505_ (.A(_05440_),
    .B(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__a22oi_4 _33506_ (.A1(_04374_),
    .A2(_04372_),
    .B1(_04344_),
    .B2(_04376_),
    .Y(_05443_));
 sky130_fd_sc_hd__xnor2_2 _33507_ (.A(_05442_),
    .B(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__and2b_1 _33508_ (.A_N(net322),
    .B(\delay_line[29][12] ),
    .X(_05445_));
 sky130_fd_sc_hd__and2b_1 _33509_ (.A_N(\delay_line[29][12] ),
    .B(\delay_line[29][8] ),
    .X(_05446_));
 sky130_fd_sc_hd__nor2_1 _33510_ (.A(_05445_),
    .B(_05446_),
    .Y(_05448_));
 sky130_fd_sc_hd__a21oi_1 _33511_ (.A1(_04410_),
    .A2(_04407_),
    .B1(_04408_),
    .Y(_05449_));
 sky130_fd_sc_hd__xnor2_1 _33512_ (.A(_05448_),
    .B(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__a311oi_1 _33513_ (.A1(_00917_),
    .A2(_02078_),
    .A3(_04411_),
    .B1(_05450_),
    .C1(_04421_),
    .Y(_05451_));
 sky130_fd_sc_hd__and3_1 _33514_ (.A(_00917_),
    .B(_02078_),
    .C(_04411_),
    .X(_05452_));
 sky130_fd_sc_hd__o21ai_1 _33515_ (.A1(_04421_),
    .A2(_05452_),
    .B1(_05450_),
    .Y(_05453_));
 sky130_fd_sc_hd__or2b_1 _33516_ (.A(_05451_),
    .B_N(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__xor2_2 _33517_ (.A(_02102_),
    .B(_02099_),
    .X(_05455_));
 sky130_fd_sc_hd__or2_1 _33518_ (.A(\delay_line[30][14] ),
    .B(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_2 _33519_ (.A(\delay_line[30][13] ),
    .X(_05457_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33520_ (.A(\delay_line[30][14] ),
    .X(_05459_));
 sky130_fd_sc_hd__nand2_1 _33521_ (.A(_05459_),
    .B(_05455_),
    .Y(_05460_));
 sky130_fd_sc_hd__nand4_2 _33522_ (.A(_05456_),
    .B(_04384_),
    .C(_05457_),
    .D(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__inv_2 _33523_ (.A(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__a22oi_4 _33524_ (.A1(_05457_),
    .A2(_04384_),
    .B1(_05460_),
    .B2(_05456_),
    .Y(_05463_));
 sky130_fd_sc_hd__a211oi_1 _33525_ (.A1(_04399_),
    .A2(_04378_),
    .B1(_00933_),
    .C1(_02092_),
    .Y(_05464_));
 sky130_fd_sc_hd__a21oi_1 _33526_ (.A1(_04378_),
    .A2(_02092_),
    .B1(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__xor2_1 _33527_ (.A(_24394_),
    .B(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__nor3_1 _33528_ (.A(_05462_),
    .B(_05463_),
    .C(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__o21a_1 _33529_ (.A1(_05462_),
    .A2(_05463_),
    .B1(_05466_),
    .X(_05468_));
 sky130_fd_sc_hd__nor2_1 _33530_ (.A(_04386_),
    .B(_04392_),
    .Y(_05470_));
 sky130_fd_sc_hd__o21a_1 _33531_ (.A1(_05467_),
    .A2(_05468_),
    .B1(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__nor3_1 _33532_ (.A(_05467_),
    .B(_05468_),
    .C(_05470_),
    .Y(_05472_));
 sky130_fd_sc_hd__nor2_1 _33533_ (.A(_05471_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__o21a_1 _33534_ (.A1(_04388_),
    .A2(net252),
    .B1(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__inv_2 _33535_ (.A(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__buf_1 _33536_ (.A(_02102_),
    .X(_05476_));
 sky130_fd_sc_hd__clkbuf_2 _33537_ (.A(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__a311o_1 _33538_ (.A1(_18453_),
    .A2(_02089_),
    .A3(_05477_),
    .B1(net252),
    .C1(_05473_),
    .X(_05478_));
 sky130_fd_sc_hd__o211ai_4 _33539_ (.A1(_04395_),
    .A2(_04398_),
    .B1(_05475_),
    .C1(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__a211o_1 _33540_ (.A1(_05475_),
    .A2(_05478_),
    .B1(_04395_),
    .C1(_04398_),
    .X(_05481_));
 sky130_fd_sc_hd__nand2_1 _33541_ (.A(_05479_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__xnor2_2 _33542_ (.A(_04403_),
    .B(_05482_),
    .Y(_05483_));
 sky130_fd_sc_hd__o2bb2ai_2 _33543_ (.A1_N(_04406_),
    .A2_N(_04405_),
    .B1(_04416_),
    .B2(_04417_),
    .Y(_05484_));
 sky130_fd_sc_hd__xor2_2 _33544_ (.A(_05483_),
    .B(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__xor2_2 _33545_ (.A(_05454_),
    .B(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__nor2_4 _33546_ (.A(_05444_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__and2_1 _33547_ (.A(_05444_),
    .B(_05486_),
    .X(_05488_));
 sky130_fd_sc_hd__nor2_2 _33548_ (.A(_05487_),
    .B(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__or2b_1 _33549_ (.A(_04310_),
    .B_N(_04337_),
    .X(_05490_));
 sky130_fd_sc_hd__o31a_2 _33550_ (.A1(_04287_),
    .A2(_04288_),
    .A3(_04339_),
    .B1(_05490_),
    .X(_05492_));
 sky130_fd_sc_hd__o21ai_1 _33551_ (.A1(_02224_),
    .A2(_02226_),
    .B1(_04324_),
    .Y(_05493_));
 sky130_fd_sc_hd__or4_2 _33552_ (.A(_18493_),
    .B(_19279_),
    .C(_19275_),
    .D(_04325_),
    .X(_05494_));
 sky130_fd_sc_hd__nor2_1 _33553_ (.A(_02217_),
    .B(\delay_line[27][14] ),
    .Y(_05495_));
 sky130_fd_sc_hd__nand2_1 _33554_ (.A(_02217_),
    .B(\delay_line[27][14] ),
    .Y(_05496_));
 sky130_fd_sc_hd__and4b_1 _33555_ (.A_N(_05495_),
    .B(_04318_),
    .C(_00971_),
    .D(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__and2_1 _33556_ (.A(_02217_),
    .B(\delay_line[27][14] ),
    .X(_05498_));
 sky130_fd_sc_hd__o22a_1 _33557_ (.A1(_04314_),
    .A2(_04315_),
    .B1(_05498_),
    .B2(_05495_),
    .X(_05499_));
 sky130_fd_sc_hd__or2_1 _33558_ (.A(_05497_),
    .B(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__buf_1 _33559_ (.A(\delay_line[27][14] ),
    .X(_05501_));
 sky130_fd_sc_hd__and4b_1 _33560_ (.A_N(_05501_),
    .B(_04317_),
    .C(_02220_),
    .D(_04319_),
    .X(_05503_));
 sky130_fd_sc_hd__a21oi_1 _33561_ (.A1(_04320_),
    .A2(_05500_),
    .B1(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__buf_1 _33562_ (.A(_23151_),
    .X(_05505_));
 sky130_fd_sc_hd__nand3_1 _33563_ (.A(_05504_),
    .B(_21241_),
    .C(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__a21o_1 _33564_ (.A1(_05505_),
    .A2(_21241_),
    .B1(_05504_),
    .X(_05507_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33565_ (.A(_04318_),
    .X(_05508_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33566_ (.A(_02219_),
    .X(_05509_));
 sky130_fd_sc_hd__nor2_1 _33567_ (.A(_05508_),
    .B(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__a31o_1 _33568_ (.A1(_04323_),
    .A2(_23147_),
    .A3(_20377_),
    .B1(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__a21o_1 _33569_ (.A1(_05506_),
    .A2(_05507_),
    .B1(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__nand3_1 _33570_ (.A(_05511_),
    .B(_05506_),
    .C(_05507_),
    .Y(_05514_));
 sky130_fd_sc_hd__nand2_1 _33571_ (.A(_05512_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__xnor2_1 _33572_ (.A(_23147_),
    .B(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__and3_1 _33573_ (.A(_05493_),
    .B(_05494_),
    .C(_05516_),
    .X(_05517_));
 sky130_fd_sc_hd__a21o_1 _33574_ (.A1(_05493_),
    .A2(_05494_),
    .B1(_05516_),
    .X(_05518_));
 sky130_fd_sc_hd__inv_2 _33575_ (.A(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__a2111oi_2 _33576_ (.A1(_02236_),
    .A2(_04311_),
    .B1(_04326_),
    .C1(_05517_),
    .D1(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__inv_2 _33577_ (.A(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__o21ai_1 _33578_ (.A1(_05517_),
    .A2(_05519_),
    .B1(_04328_),
    .Y(_05522_));
 sky130_fd_sc_hd__o21bai_1 _33579_ (.A1(_04332_),
    .A2(_04336_),
    .B1_N(_04331_),
    .Y(_05523_));
 sky130_fd_sc_hd__a21o_1 _33580_ (.A1(_05521_),
    .A2(_05522_),
    .B1(_05523_),
    .X(_05525_));
 sky130_fd_sc_hd__and3_1 _33581_ (.A(_05521_),
    .B(_05522_),
    .C(_05523_),
    .X(_05526_));
 sky130_fd_sc_hd__inv_2 _33582_ (.A(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__or3_1 _33583_ (.A(_02200_),
    .B(_02190_),
    .C(_02203_),
    .X(_05528_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33584_ (.A(_04290_),
    .X(_05529_));
 sky130_fd_sc_hd__o32a_1 _33585_ (.A1(_04298_),
    .A2(_04300_),
    .A3(_05528_),
    .B1(_05529_),
    .B2(_04303_),
    .X(_05530_));
 sky130_fd_sc_hd__clkbuf_2 _33586_ (.A(net335),
    .X(_05531_));
 sky130_fd_sc_hd__or2_1 _33587_ (.A(_23140_),
    .B(net337),
    .X(_05532_));
 sky130_fd_sc_hd__nand2_1 _33588_ (.A(_23140_),
    .B(net337),
    .Y(_05533_));
 sky130_fd_sc_hd__nand3_1 _33589_ (.A(_05532_),
    .B(_05533_),
    .C(_19264_),
    .Y(_05534_));
 sky130_fd_sc_hd__a21o_1 _33590_ (.A1(_05532_),
    .A2(_05533_),
    .B1(_19264_),
    .X(_05536_));
 sky130_fd_sc_hd__nand2_1 _33591_ (.A(_05534_),
    .B(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__a21oi_1 _33592_ (.A1(_04292_),
    .A2(_04299_),
    .B1(_05537_),
    .Y(_05538_));
 sky130_fd_sc_hd__and3_1 _33593_ (.A(_04292_),
    .B(_04299_),
    .C(_05537_),
    .X(_05539_));
 sky130_fd_sc_hd__nor2_1 _33594_ (.A(_05538_),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__a32o_1 _33595_ (.A1(_04299_),
    .A2(_04296_),
    .A3(_04297_),
    .B1(_04301_),
    .B2(_02203_),
    .X(_05541_));
 sky130_fd_sc_hd__xor2_1 _33596_ (.A(_05540_),
    .B(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__xor2_1 _33597_ (.A(_05531_),
    .B(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__and2b_1 _33598_ (.A_N(_05530_),
    .B(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__or2b_1 _33599_ (.A(_05543_),
    .B_N(_05530_),
    .X(_05545_));
 sky130_fd_sc_hd__inv_2 _33600_ (.A(_05545_),
    .Y(_05547_));
 sky130_fd_sc_hd__nor2_1 _33601_ (.A(_05544_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__and2b_1 _33602_ (.A_N(_04306_),
    .B(_04304_),
    .X(_05549_));
 sky130_fd_sc_hd__a21oi_1 _33603_ (.A1(_04309_),
    .A2(_04307_),
    .B1(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__xnor2_1 _33604_ (.A(_05548_),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__nand3_1 _33605_ (.A(_05525_),
    .B(_05527_),
    .C(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__a21oi_1 _33606_ (.A1(_05525_),
    .A2(_05527_),
    .B1(_05551_),
    .Y(_05553_));
 sky130_fd_sc_hd__inv_2 _33607_ (.A(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2_2 _33608_ (.A(_05552_),
    .B(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__o211a_1 _33609_ (.A1(_01038_),
    .A2(_01041_),
    .B1(_02180_),
    .C1(_04284_),
    .X(_05556_));
 sky130_fd_sc_hd__nand2_1 _33610_ (.A(_04269_),
    .B(_04273_),
    .Y(_05558_));
 sky130_fd_sc_hd__buf_1 _33611_ (.A(_04270_),
    .X(_05559_));
 sky130_fd_sc_hd__buf_1 _33612_ (.A(\delay_line[28][14] ),
    .X(_05560_));
 sky130_fd_sc_hd__buf_1 _33613_ (.A(net324),
    .X(_05561_));
 sky130_fd_sc_hd__or3b_1 _33614_ (.A(_05559_),
    .B(_05560_),
    .C_N(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__nand3_1 _33615_ (.A(_05559_),
    .B(\delay_line[28][13] ),
    .C(\delay_line[28][14] ),
    .Y(_05563_));
 sky130_fd_sc_hd__o21a_1 _33616_ (.A1(_05561_),
    .A2(_05560_),
    .B1(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_2 _33617_ (.A(_23178_),
    .X(_05565_));
 sky130_fd_sc_hd__and3_1 _33618_ (.A(_05562_),
    .B(_05564_),
    .C(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__a21oi_2 _33619_ (.A1(_05562_),
    .A2(_05564_),
    .B1(_05565_),
    .Y(_05567_));
 sky130_fd_sc_hd__a211oi_4 _33620_ (.A1(_04274_),
    .A2(_05558_),
    .B1(_05566_),
    .C1(_05567_),
    .Y(_05569_));
 sky130_fd_sc_hd__o211a_1 _33621_ (.A1(_05566_),
    .A2(_05567_),
    .B1(_04274_),
    .C1(_05558_),
    .X(_05570_));
 sky130_fd_sc_hd__nor3b_2 _33622_ (.A(_05569_),
    .B(_05570_),
    .C_N(_04269_),
    .Y(_05571_));
 sky130_fd_sc_hd__o21bai_1 _33623_ (.A1(_05569_),
    .A2(_05570_),
    .B1_N(_04269_),
    .Y(_05572_));
 sky130_fd_sc_hd__nand2b_1 _33624_ (.A_N(_05571_),
    .B(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__nor2b_1 _33625_ (.A(_04277_),
    .B_N(_04280_),
    .Y(_05574_));
 sky130_fd_sc_hd__xor2_1 _33626_ (.A(_05573_),
    .B(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__o2111a_1 _33627_ (.A1(_02176_),
    .A2(net230),
    .B1(_04279_),
    .C1(_04280_),
    .D1(_05575_),
    .X(_05576_));
 sky130_fd_sc_hd__nor2_1 _33628_ (.A(_04281_),
    .B(_05575_),
    .Y(_05577_));
 sky130_fd_sc_hd__or2_1 _33629_ (.A(_05576_),
    .B(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__nor3b_1 _33630_ (.A(_05556_),
    .B(_04287_),
    .C_N(_05578_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21ba_1 _33631_ (.A1(_05556_),
    .A2(_04287_),
    .B1_N(_05578_),
    .X(_05581_));
 sky130_fd_sc_hd__or2_2 _33632_ (.A(_05580_),
    .B(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__xnor2_4 _33633_ (.A(_05555_),
    .B(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__xnor2_4 _33634_ (.A(_05492_),
    .B(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__xnor2_4 _33635_ (.A(_05489_),
    .B(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__o21a_1 _33636_ (.A1(_04254_),
    .A2(_04256_),
    .B1(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__nor3_1 _33637_ (.A(_04254_),
    .B(_04256_),
    .C(_05585_),
    .Y(_05587_));
 sky130_fd_sc_hd__or2_1 _33638_ (.A(_05586_),
    .B(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__a21o_2 _33639_ (.A1(_04343_),
    .A2(_04430_),
    .B1(_04342_),
    .X(_05589_));
 sky130_fd_sc_hd__xnor2_1 _33640_ (.A(_05588_),
    .B(_05589_),
    .Y(_05591_));
 sky130_fd_sc_hd__o21a_1 _33641_ (.A1(_04258_),
    .A2(_04136_),
    .B1(_04133_),
    .X(_05592_));
 sky130_fd_sc_hd__inv_2 _33642_ (.A(_04120_),
    .Y(_05593_));
 sky130_fd_sc_hd__a21oi_1 _33643_ (.A1(_18362_),
    .A2(_04119_),
    .B1(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_2 _33644_ (.A(_18361_),
    .B(_04086_),
    .Y(_05595_));
 sky130_fd_sc_hd__o22a_1 _33645_ (.A1(_18361_),
    .A2(_04090_),
    .B1(_20513_),
    .B2(_20515_),
    .X(_05596_));
 sky130_fd_sc_hd__buf_1 _33646_ (.A(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33647_ (.A(_04090_),
    .X(_05598_));
 sky130_fd_sc_hd__a21oi_1 _33648_ (.A1(_18361_),
    .A2(_05598_),
    .B1(_18350_),
    .Y(_05599_));
 sky130_fd_sc_hd__buf_1 _33649_ (.A(\delay_line[21][13] ),
    .X(_05600_));
 sky130_fd_sc_hd__nor2_1 _33650_ (.A(_04103_),
    .B(_05600_),
    .Y(_05602_));
 sky130_fd_sc_hd__and2_1 _33651_ (.A(\delay_line[21][12] ),
    .B(_05600_),
    .X(_05603_));
 sky130_fd_sc_hd__a2bb2o_1 _33652_ (.A1_N(_05602_),
    .A2_N(_05603_),
    .B1(_04106_),
    .B2(_04094_),
    .X(_05604_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33653_ (.A(\delay_line[21][13] ),
    .X(_05605_));
 sky130_fd_sc_hd__nand2_2 _33654_ (.A(_04095_),
    .B(_04103_),
    .Y(_05606_));
 sky130_fd_sc_hd__or2_1 _33655_ (.A(_05605_),
    .B(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__and3_1 _33656_ (.A(_05604_),
    .B(_05607_),
    .C(_22992_),
    .X(_05608_));
 sky130_fd_sc_hd__clkbuf_2 _33657_ (.A(_22992_),
    .X(_05609_));
 sky130_fd_sc_hd__a21oi_2 _33658_ (.A1(_05604_),
    .A2(_05607_),
    .B1(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__a211o_1 _33659_ (.A1(_04104_),
    .A2(_04102_),
    .B1(_05608_),
    .C1(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__o221ai_4 _33660_ (.A1(_04097_),
    .A2(_04094_),
    .B1(_05610_),
    .B2(_05608_),
    .C1(_04102_),
    .Y(_05613_));
 sky130_fd_sc_hd__buf_1 _33661_ (.A(_21411_),
    .X(_05614_));
 sky130_fd_sc_hd__or3b_1 _33662_ (.A(_21410_),
    .B(_05614_),
    .C_N(_21412_),
    .X(_05615_));
 sky130_fd_sc_hd__nor2_1 _33663_ (.A(_21410_),
    .B(_05614_),
    .Y(_05616_));
 sky130_fd_sc_hd__or2_1 _33664_ (.A(_04090_),
    .B(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__nor2_1 _33665_ (.A(_20513_),
    .B(_20515_),
    .Y(_05618_));
 sky130_fd_sc_hd__a21oi_2 _33666_ (.A1(_18348_),
    .A2(_05618_),
    .B1(_20513_),
    .Y(_05619_));
 sky130_fd_sc_hd__a21oi_1 _33667_ (.A1(_05615_),
    .A2(_05617_),
    .B1(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__and3_1 _33668_ (.A(_05619_),
    .B(_05615_),
    .C(_05617_),
    .X(_05621_));
 sky130_fd_sc_hd__nor2_1 _33669_ (.A(_05620_),
    .B(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__a21o_1 _33670_ (.A1(_05611_),
    .A2(_05613_),
    .B1(_05622_),
    .X(_05624_));
 sky130_fd_sc_hd__nand2_1 _33671_ (.A(_04092_),
    .B(_04093_),
    .Y(_05625_));
 sky130_fd_sc_hd__a32oi_2 _33672_ (.A1(_04102_),
    .A2(_04105_),
    .A3(_04108_),
    .B1(_04110_),
    .B2(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__nand3_1 _33673_ (.A(_05611_),
    .B(_05613_),
    .C(_05622_),
    .Y(_05627_));
 sky130_fd_sc_hd__nand3_1 _33674_ (.A(_05624_),
    .B(_05626_),
    .C(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__a21o_1 _33675_ (.A1(_05627_),
    .A2(_05624_),
    .B1(_05626_),
    .X(_05629_));
 sky130_fd_sc_hd__o211a_1 _33676_ (.A1(_05597_),
    .A2(_05599_),
    .B1(_05628_),
    .C1(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__or2_1 _33677_ (.A(_05596_),
    .B(_05599_),
    .X(_05631_));
 sky130_fd_sc_hd__a21oi_1 _33678_ (.A1(_05628_),
    .A2(_05629_),
    .B1(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__nor2_1 _33679_ (.A(_05630_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__a41o_1 _33680_ (.A1(_02549_),
    .A2(_04088_),
    .A3(_04111_),
    .A4(_04112_),
    .B1(_04087_),
    .X(_05635_));
 sky130_fd_sc_hd__nand3_1 _33681_ (.A(_05633_),
    .B(_05635_),
    .C(_04114_),
    .Y(_05636_));
 sky130_fd_sc_hd__o2bb2ai_1 _33682_ (.A1_N(_04114_),
    .A2_N(_05635_),
    .B1(_05630_),
    .B2(_05632_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_1 _33683_ (.A(_05636_),
    .B(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__xor2_2 _33684_ (.A(_05595_),
    .B(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__xnor2_2 _33685_ (.A(_05594_),
    .B(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__o21bai_2 _33686_ (.A1(_04124_),
    .A2(_04126_),
    .B1_N(_04123_),
    .Y(_05641_));
 sky130_fd_sc_hd__xnor2_1 _33687_ (.A(_05640_),
    .B(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__and3_1 _33688_ (.A(_04027_),
    .B(_04028_),
    .C(_04029_),
    .X(_05643_));
 sky130_fd_sc_hd__nand2_1 _33689_ (.A(_04016_),
    .B(_04020_),
    .Y(_05644_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33690_ (.A(\delay_line[18][13] ),
    .X(_05646_));
 sky130_fd_sc_hd__nor2_1 _33691_ (.A(_24694_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand2_1 _33692_ (.A(_24694_),
    .B(\delay_line[18][13] ),
    .Y(_05648_));
 sky130_fd_sc_hd__nor3b_1 _33693_ (.A(_05647_),
    .B(_04015_),
    .C_N(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__or2_1 _33694_ (.A(_24694_),
    .B(_05646_),
    .X(_05650_));
 sky130_fd_sc_hd__a22o_1 _33695_ (.A1(_22931_),
    .A2(_04013_),
    .B1(_05648_),
    .B2(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__a21oi_1 _33696_ (.A1(_18388_),
    .A2(_19391_),
    .B1(_20542_),
    .Y(_05652_));
 sky130_fd_sc_hd__and3_1 _33697_ (.A(_18387_),
    .B(_19391_),
    .C(_21362_),
    .X(_05653_));
 sky130_fd_sc_hd__nor2_1 _33698_ (.A(_05652_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand3b_1 _33699_ (.A_N(net277),
    .B(_05651_),
    .C(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__a21oi_1 _33700_ (.A1(_05648_),
    .A2(_05650_),
    .B1(_04017_),
    .Y(_05657_));
 sky130_fd_sc_hd__o22ai_2 _33701_ (.A1(_05652_),
    .A2(_05653_),
    .B1(net277),
    .B2(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand3_2 _33702_ (.A(_05644_),
    .B(_05655_),
    .C(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2_1 _33703_ (.A(_05655_),
    .B(_05658_),
    .Y(_05660_));
 sky130_fd_sc_hd__nand3_2 _33704_ (.A(_04016_),
    .B(_04020_),
    .C(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__o2111ai_4 _33705_ (.A1(_16338_),
    .A2(_21354_),
    .B1(_18385_),
    .C1(_05659_),
    .D1(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__and3_1 _33706_ (.A(_19395_),
    .B(_18384_),
    .C(_24704_),
    .X(_05663_));
 sky130_fd_sc_hd__o2bb2ai_1 _33707_ (.A1_N(_05661_),
    .A2_N(_05659_),
    .B1(_18389_),
    .B2(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__a211o_1 _33708_ (.A1(_05662_),
    .A2(_05664_),
    .B1(_04024_),
    .C1(_04025_),
    .X(_05665_));
 sky130_fd_sc_hd__o211ai_1 _33709_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_05662_),
    .C1(_05664_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_1 _33710_ (.A(_05665_),
    .B(_05666_),
    .Y(_05668_));
 sky130_fd_sc_hd__xor2_1 _33711_ (.A(_04010_),
    .B(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__nand2_1 _33712_ (.A(_04027_),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__a21o_1 _33713_ (.A1(_04027_),
    .A2(_04031_),
    .B1(_05669_),
    .X(_05671_));
 sky130_fd_sc_hd__o21a_1 _33714_ (.A1(_05643_),
    .A2(_05670_),
    .B1(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__a21boi_1 _33715_ (.A1(_02632_),
    .A2(_02659_),
    .B1_N(_02662_),
    .Y(_05673_));
 sky130_fd_sc_hd__o21bai_1 _33716_ (.A1(_04034_),
    .A2(_05673_),
    .B1_N(_04035_),
    .Y(_05674_));
 sky130_fd_sc_hd__nor2_1 _33717_ (.A(_05672_),
    .B(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__or2_1 _33718_ (.A(_04071_),
    .B(_04072_),
    .X(_05676_));
 sky130_fd_sc_hd__o22a_1 _33719_ (.A1(_18380_),
    .A2(_00668_),
    .B1(_20548_),
    .B2(_20549_),
    .X(_05677_));
 sky130_fd_sc_hd__a21o_1 _33720_ (.A1(_19400_),
    .A2(_04039_),
    .B1(_05677_),
    .X(_05679_));
 sky130_fd_sc_hd__buf_1 _33721_ (.A(_21374_),
    .X(_05680_));
 sky130_fd_sc_hd__or3_1 _33722_ (.A(_19405_),
    .B(_05680_),
    .C(_22953_),
    .X(_05681_));
 sky130_fd_sc_hd__o21ai_1 _33723_ (.A1(_05680_),
    .A2(_22953_),
    .B1(_19405_),
    .Y(_05682_));
 sky130_fd_sc_hd__o21a_1 _33724_ (.A1(_18370_),
    .A2(_20549_),
    .B1(_21376_),
    .X(_05683_));
 sky130_fd_sc_hd__a21oi_1 _33725_ (.A1(_05681_),
    .A2(_05682_),
    .B1(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__and3_1 _33726_ (.A(_05681_),
    .B(_05682_),
    .C(_05683_),
    .X(_05685_));
 sky130_fd_sc_hd__nor2_1 _33727_ (.A(_05684_),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__nor2_1 _33728_ (.A(_04045_),
    .B(net369),
    .Y(_05687_));
 sky130_fd_sc_hd__and2_2 _33729_ (.A(\delay_line[19][12] ),
    .B(net369),
    .X(_05688_));
 sky130_fd_sc_hd__o21bai_2 _33730_ (.A1(_05687_),
    .A2(_05688_),
    .B1_N(_04048_),
    .Y(_05690_));
 sky130_fd_sc_hd__clkbuf_2 _33731_ (.A(_04048_),
    .X(_05691_));
 sky130_fd_sc_hd__inv_2 _33732_ (.A(net369),
    .Y(_05692_));
 sky130_fd_sc_hd__nand2_1 _33733_ (.A(_05691_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__and3_1 _33734_ (.A(_05690_),
    .B(_05693_),
    .C(_22946_),
    .X(_05694_));
 sky130_fd_sc_hd__a21oi_2 _33735_ (.A1(_05690_),
    .A2(_05693_),
    .B1(_22946_),
    .Y(_05695_));
 sky130_fd_sc_hd__a211o_1 _33736_ (.A1(_04051_),
    .A2(_04050_),
    .B1(_05694_),
    .C1(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__clkbuf_2 _33737_ (.A(_04046_),
    .X(_05697_));
 sky130_fd_sc_hd__clkbuf_2 _33738_ (.A(_04045_),
    .X(_05698_));
 sky130_fd_sc_hd__o221ai_4 _33739_ (.A1(_05697_),
    .A2(_05698_),
    .B1(_05695_),
    .B2(_05694_),
    .C1(_04050_),
    .Y(_05699_));
 sky130_fd_sc_hd__and3_1 _33740_ (.A(_05686_),
    .B(_05696_),
    .C(_05699_),
    .X(_05701_));
 sky130_fd_sc_hd__a21oi_1 _33741_ (.A1(_05696_),
    .A2(_05699_),
    .B1(_05686_),
    .Y(_05702_));
 sky130_fd_sc_hd__nor2_1 _33742_ (.A(_05701_),
    .B(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__a21bo_1 _33743_ (.A1(_04040_),
    .A2(_04042_),
    .B1_N(_04058_),
    .X(_05704_));
 sky130_fd_sc_hd__nand3_1 _33744_ (.A(_05703_),
    .B(_05704_),
    .C(_04054_),
    .Y(_05705_));
 sky130_fd_sc_hd__o2bb2ai_1 _33745_ (.A1_N(_04054_),
    .A2_N(_05704_),
    .B1(_05701_),
    .B2(_05702_),
    .Y(_05706_));
 sky130_fd_sc_hd__and3_1 _33746_ (.A(_05679_),
    .B(_05705_),
    .C(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__a21oi_1 _33747_ (.A1(_05705_),
    .A2(_05706_),
    .B1(_05679_),
    .Y(_05708_));
 sky130_fd_sc_hd__nor2_1 _33748_ (.A(_05707_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__a41o_1 _33749_ (.A1(_02596_),
    .A2(_02610_),
    .A3(_04059_),
    .A4(_04060_),
    .B1(_04066_),
    .X(_05710_));
 sky130_fd_sc_hd__nand3_1 _33750_ (.A(_05709_),
    .B(_05710_),
    .C(_04062_),
    .Y(_05712_));
 sky130_fd_sc_hd__o2bb2ai_2 _33751_ (.A1_N(_04062_),
    .A2_N(_05710_),
    .B1(_05707_),
    .B2(_05708_),
    .Y(_05713_));
 sky130_fd_sc_hd__o221a_1 _33752_ (.A1(_07470_),
    .A2(_20574_),
    .B1(_19401_),
    .B2(_19403_),
    .C1(_18380_),
    .X(_05714_));
 sky130_fd_sc_hd__and3_1 _33753_ (.A(_05712_),
    .B(_05713_),
    .C(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__a21oi_1 _33754_ (.A1(_05712_),
    .A2(_05713_),
    .B1(_05714_),
    .Y(_05716_));
 sky130_fd_sc_hd__nor2_1 _33755_ (.A(_05715_),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__xnor2_1 _33756_ (.A(_05676_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__o21ai_1 _33757_ (.A1(_04073_),
    .A2(_04080_),
    .B1(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__o211ai_1 _33758_ (.A1(_04080_),
    .A2(_04073_),
    .B1(_04076_),
    .C1(_04078_),
    .Y(_05720_));
 sky130_fd_sc_hd__a21oi_1 _33759_ (.A1(_04077_),
    .A2(_05720_),
    .B1(_05718_),
    .Y(_05721_));
 sky130_fd_sc_hd__o21bai_2 _33760_ (.A1(_04079_),
    .A2(_05719_),
    .B1_N(_05721_),
    .Y(_05723_));
 sky130_fd_sc_hd__o21ai_1 _33761_ (.A1(_04035_),
    .A2(_04036_),
    .B1(_05672_),
    .Y(_05724_));
 sky130_fd_sc_hd__or3b_4 _33762_ (.A(_05675_),
    .B(_05723_),
    .C_N(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__or2b_1 _33763_ (.A(_05675_),
    .B_N(_05724_),
    .X(_05726_));
 sky130_fd_sc_hd__nand2_1 _33764_ (.A(_05726_),
    .B(_05723_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand2_1 _33765_ (.A(_05725_),
    .B(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__or2_4 _33766_ (.A(_05642_),
    .B(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__nand2_1 _33767_ (.A(_05642_),
    .B(_05728_),
    .Y(_05730_));
 sky130_fd_sc_hd__o21ai_1 _33768_ (.A1(_02528_),
    .A2(_03873_),
    .B1(_03919_),
    .Y(_05731_));
 sky130_fd_sc_hd__and3_1 _33769_ (.A(_03915_),
    .B(_03912_),
    .C(_03914_),
    .X(_05732_));
 sky130_fd_sc_hd__and2_1 _33770_ (.A(_03911_),
    .B(_03912_),
    .X(_05734_));
 sky130_fd_sc_hd__nand2_1 _33771_ (.A(_03913_),
    .B(_03875_),
    .Y(_05735_));
 sky130_fd_sc_hd__or2_1 _33772_ (.A(_03913_),
    .B(_03875_),
    .X(_05736_));
 sky130_fd_sc_hd__nand2_1 _33773_ (.A(_03894_),
    .B(_03896_),
    .Y(_05737_));
 sky130_fd_sc_hd__and2_1 _33774_ (.A(_24819_),
    .B(net382),
    .X(_05738_));
 sky130_fd_sc_hd__inv_2 _33775_ (.A(\delay_line[16][9] ),
    .Y(_05739_));
 sky130_fd_sc_hd__nand2_1 _33776_ (.A(_05739_),
    .B(_02497_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand3b_1 _33777_ (.A_N(_05738_),
    .B(_23023_),
    .C(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__nor2_1 _33778_ (.A(_24819_),
    .B(net382),
    .Y(_05742_));
 sky130_fd_sc_hd__o21bai_2 _33779_ (.A1(_05742_),
    .A2(_05738_),
    .B1_N(_23023_),
    .Y(_05743_));
 sky130_fd_sc_hd__buf_1 _33780_ (.A(\delay_line[16][13] ),
    .X(_05745_));
 sky130_fd_sc_hd__and3_1 _33781_ (.A(_05741_),
    .B(_05743_),
    .C(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33782_ (.A(_05745_),
    .X(_05747_));
 sky130_fd_sc_hd__a21o_1 _33783_ (.A1(_05741_),
    .A2(_05743_),
    .B1(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__nand3b_2 _33784_ (.A_N(_05746_),
    .B(_05748_),
    .C(_03883_),
    .Y(_05749_));
 sky130_fd_sc_hd__a21oi_1 _33785_ (.A1(_05741_),
    .A2(_05743_),
    .B1(_05747_),
    .Y(_05750_));
 sky130_fd_sc_hd__o21ai_2 _33786_ (.A1(_05746_),
    .A2(_05750_),
    .B1(_03890_),
    .Y(_05751_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33787_ (.A(_23026_),
    .X(_05752_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33788_ (.A(_24821_),
    .X(_05753_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33789_ (.A(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__clkbuf_2 _33790_ (.A(_21518_),
    .X(_05756_));
 sky130_fd_sc_hd__a21oi_1 _33791_ (.A1(_05752_),
    .A2(_05754_),
    .B1(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__o21a_1 _33792_ (.A1(_23026_),
    .A2(_05753_),
    .B1(_21518_),
    .X(_05758_));
 sky130_fd_sc_hd__o2bb2ai_1 _33793_ (.A1_N(_05749_),
    .A2_N(_05751_),
    .B1(_05757_),
    .B2(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__o2111ai_4 _33794_ (.A1(_05756_),
    .A2(_03878_),
    .B1(_03879_),
    .C1(_05749_),
    .D1(_05751_),
    .Y(_05760_));
 sky130_fd_sc_hd__nand3_1 _33795_ (.A(_05737_),
    .B(_05759_),
    .C(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__a21o_1 _33796_ (.A1(_05759_),
    .A2(_05760_),
    .B1(_05737_),
    .X(_05762_));
 sky130_fd_sc_hd__nand4_2 _33797_ (.A(_05735_),
    .B(_05736_),
    .C(_05761_),
    .D(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__a22o_1 _33798_ (.A1(_05735_),
    .A2(_05736_),
    .B1(_05761_),
    .B2(_05762_),
    .X(_05764_));
 sky130_fd_sc_hd__nand2_1 _33799_ (.A(_03905_),
    .B(_03906_),
    .Y(_05765_));
 sky130_fd_sc_hd__a21o_1 _33800_ (.A1(_05763_),
    .A2(_05764_),
    .B1(_05765_),
    .X(_05767_));
 sky130_fd_sc_hd__nand3_1 _33801_ (.A(_05765_),
    .B(_05763_),
    .C(_05764_),
    .Y(_05768_));
 sky130_fd_sc_hd__and3_1 _33802_ (.A(_05767_),
    .B(_05768_),
    .C(_03902_),
    .X(_05769_));
 sky130_fd_sc_hd__a21oi_1 _33803_ (.A1(_05767_),
    .A2(_05768_),
    .B1(_03902_),
    .Y(_05770_));
 sky130_fd_sc_hd__nor2_1 _33804_ (.A(_05769_),
    .B(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__xnor2_2 _33805_ (.A(_05734_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__nor2_1 _33806_ (.A(_05732_),
    .B(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__o21a_1 _33807_ (.A1(_05732_),
    .A2(_03918_),
    .B1(_05772_),
    .X(_05774_));
 sky130_fd_sc_hd__nand2_1 _33808_ (.A(_18408_),
    .B(_02410_),
    .Y(_05775_));
 sky130_fd_sc_hd__a21oi_1 _33809_ (.A1(_03923_),
    .A2(_23054_),
    .B1(_19452_),
    .Y(_05776_));
 sky130_fd_sc_hd__and3_1 _33810_ (.A(_19451_),
    .B(_21497_),
    .C(_23054_),
    .X(_05778_));
 sky130_fd_sc_hd__nor2_1 _33811_ (.A(net390),
    .B(_24783_),
    .Y(_05779_));
 sky130_fd_sc_hd__and2_1 _33812_ (.A(\delay_line[14][8] ),
    .B(\delay_line[14][9] ),
    .X(_05780_));
 sky130_fd_sc_hd__or3b_1 _33813_ (.A(_05779_),
    .B(_05780_),
    .C_N(\delay_line[14][13] ),
    .X(_05781_));
 sky130_fd_sc_hd__o21bai_1 _33814_ (.A1(_05779_),
    .A2(_05780_),
    .B1_N(\delay_line[14][13] ),
    .Y(_05782_));
 sky130_fd_sc_hd__nand3b_1 _33815_ (.A_N(_03929_),
    .B(_05781_),
    .C(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__a21boi_1 _33816_ (.A1(_05781_),
    .A2(_05782_),
    .B1_N(_03929_),
    .Y(_05784_));
 sky130_fd_sc_hd__inv_2 _33817_ (.A(_05784_),
    .Y(_05785_));
 sky130_fd_sc_hd__or4bb_1 _33818_ (.A(_05776_),
    .B(_05778_),
    .C_N(_05783_),
    .D_N(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__buf_1 _33819_ (.A(_05778_),
    .X(_05787_));
 sky130_fd_sc_hd__a2bb2o_1 _33820_ (.A1_N(_05776_),
    .A2_N(_05787_),
    .B1(_05783_),
    .B2(_05785_),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_1 _33821_ (.A(_05786_),
    .B(_05789_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand3_1 _33822_ (.A(_03932_),
    .B(_03935_),
    .C(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__a21o_1 _33823_ (.A1(_03932_),
    .A2(_03935_),
    .B1(_05790_),
    .X(_05792_));
 sky130_fd_sc_hd__nand2_1 _33824_ (.A(_05791_),
    .B(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__xor2_1 _33825_ (.A(_05775_),
    .B(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__nor2_1 _33826_ (.A(_03940_),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__a21boi_2 _33827_ (.A1(_03939_),
    .A2(_03941_),
    .B1_N(_05794_),
    .Y(_05796_));
 sky130_fd_sc_hd__a21oi_4 _33828_ (.A1(_03941_),
    .A2(_05795_),
    .B1(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__o21bai_4 _33829_ (.A1(_03945_),
    .A2(_03950_),
    .B1_N(_03946_),
    .Y(_05798_));
 sky130_fd_sc_hd__xor2_4 _33830_ (.A(_05797_),
    .B(_05798_),
    .X(_05800_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33831_ (.A(_03971_),
    .X(_05801_));
 sky130_fd_sc_hd__or3_2 _33832_ (.A(_05801_),
    .B(_21454_),
    .C(_18429_),
    .X(_05802_));
 sky130_fd_sc_hd__nand2_1 _33833_ (.A(_03967_),
    .B(_03976_),
    .Y(_05803_));
 sky130_fd_sc_hd__nor3_1 _33834_ (.A(_03958_),
    .B(_03955_),
    .C(_03956_),
    .Y(_05804_));
 sky130_fd_sc_hd__buf_1 _33835_ (.A(\delay_line[15][14] ),
    .X(_05805_));
 sky130_fd_sc_hd__nor2_1 _33836_ (.A(_03957_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__nand2_1 _33837_ (.A(_03957_),
    .B(_05805_),
    .Y(_05807_));
 sky130_fd_sc_hd__nand3b_1 _33838_ (.A_N(_05806_),
    .B(_03956_),
    .C(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__and2_2 _33839_ (.A(_02431_),
    .B(\delay_line[15][14] ),
    .X(_05809_));
 sky130_fd_sc_hd__o21ai_1 _33840_ (.A1(_05809_),
    .A2(_05806_),
    .B1(_03961_),
    .Y(_05811_));
 sky130_fd_sc_hd__a21o_1 _33841_ (.A1(_05808_),
    .A2(_05811_),
    .B1(_23076_),
    .X(_05812_));
 sky130_fd_sc_hd__buf_1 _33842_ (.A(_23076_),
    .X(_05813_));
 sky130_fd_sc_hd__nand3_1 _33843_ (.A(_05811_),
    .B(_05813_),
    .C(_05808_),
    .Y(_05814_));
 sky130_fd_sc_hd__o211ai_1 _33844_ (.A1(_05804_),
    .A2(_03968_),
    .B1(_05812_),
    .C1(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__a21o_1 _33845_ (.A1(_03959_),
    .A2(_03960_),
    .B1(_05804_),
    .X(_05816_));
 sky130_fd_sc_hd__a21o_1 _33846_ (.A1(_05812_),
    .A2(_05814_),
    .B1(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__o21a_1 _33847_ (.A1(_20603_),
    .A2(_20604_),
    .B1(_03971_),
    .X(_05818_));
 sky130_fd_sc_hd__clkbuf_2 _33848_ (.A(_02433_),
    .X(_05819_));
 sky130_fd_sc_hd__nor2_1 _33849_ (.A(_05801_),
    .B(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__o2bb2ai_1 _33850_ (.A1_N(_05815_),
    .A2_N(_05817_),
    .B1(_05818_),
    .B2(_05820_),
    .Y(_05822_));
 sky130_fd_sc_hd__clkbuf_2 _33851_ (.A(_20596_),
    .X(_05823_));
 sky130_fd_sc_hd__nor2_1 _33852_ (.A(_05801_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__and3_1 _33853_ (.A(_20597_),
    .B(_20601_),
    .C(_03971_),
    .X(_05825_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33854_ (.A(_05815_),
    .X(_05826_));
 sky130_fd_sc_hd__o211ai_1 _33855_ (.A1(_05824_),
    .A2(_05825_),
    .B1(_05826_),
    .C1(_05817_),
    .Y(_05827_));
 sky130_fd_sc_hd__nand3_1 _33856_ (.A(_05803_),
    .B(_05822_),
    .C(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__o2bb2ai_1 _33857_ (.A1_N(_05826_),
    .A2_N(_05817_),
    .B1(_05824_),
    .B2(_05825_),
    .Y(_05829_));
 sky130_fd_sc_hd__a21boi_1 _33858_ (.A1(_03970_),
    .A2(_03974_),
    .B1_N(_03967_),
    .Y(_05830_));
 sky130_fd_sc_hd__o211ai_1 _33859_ (.A1(_05818_),
    .A2(_05820_),
    .B1(_05826_),
    .C1(_05817_),
    .Y(_05831_));
 sky130_fd_sc_hd__nand3_1 _33860_ (.A(_05829_),
    .B(_05830_),
    .C(_05831_),
    .Y(_05833_));
 sky130_fd_sc_hd__a22oi_2 _33861_ (.A1(_05802_),
    .A2(_19467_),
    .B1(_05828_),
    .B2(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__and4_1 _33862_ (.A(_05802_),
    .B(_05833_),
    .C(_05828_),
    .D(_19467_),
    .X(_05835_));
 sky130_fd_sc_hd__o221a_1 _33863_ (.A1(_03987_),
    .A2(_03985_),
    .B1(_05834_),
    .B2(_05835_),
    .C1(_03983_),
    .X(_05836_));
 sky130_fd_sc_hd__a211o_1 _33864_ (.A1(_03982_),
    .A2(_03983_),
    .B1(_05835_),
    .C1(_05834_),
    .X(_05837_));
 sky130_fd_sc_hd__and2b_1 _33865_ (.A_N(_05836_),
    .B(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__xor2_2 _33866_ (.A(_03981_),
    .B(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__o21ai_2 _33867_ (.A1(_02467_),
    .A2(_03993_),
    .B1(_03992_),
    .Y(_05840_));
 sky130_fd_sc_hd__xor2_2 _33868_ (.A(_05839_),
    .B(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__a21boi_2 _33869_ (.A1(_03952_),
    .A2(_03998_),
    .B1_N(_03995_),
    .Y(_05842_));
 sky130_fd_sc_hd__xor2_2 _33870_ (.A(_05841_),
    .B(_05842_),
    .X(_05844_));
 sky130_fd_sc_hd__xnor2_1 _33871_ (.A(_05800_),
    .B(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__a211oi_1 _33872_ (.A1(_05731_),
    .A2(_05773_),
    .B1(_05774_),
    .C1(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_1 _33873_ (.A(_03916_),
    .B(_03917_),
    .Y(_05847_));
 sky130_fd_sc_hd__a31oi_2 _33874_ (.A1(_03872_),
    .A2(_02529_),
    .A3(_00863_),
    .B1(_02527_),
    .Y(_05848_));
 sky130_fd_sc_hd__o21a_1 _33875_ (.A1(_05847_),
    .A2(_05848_),
    .B1(_05773_),
    .X(_05849_));
 sky130_fd_sc_hd__o21a_1 _33876_ (.A1(_05849_),
    .A2(_05774_),
    .B1(_05845_),
    .X(_05850_));
 sky130_fd_sc_hd__nor2_1 _33877_ (.A(_05846_),
    .B(_05850_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21ai_2 _33878_ (.A1(_03951_),
    .A2(_03999_),
    .B1(_04002_),
    .Y(_05852_));
 sky130_fd_sc_hd__and2_1 _33879_ (.A(_05851_),
    .B(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__or2_1 _33880_ (.A(_05852_),
    .B(_05851_),
    .X(_05855_));
 sky130_fd_sc_hd__and2b_1 _33881_ (.A_N(_05853_),
    .B(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__a21oi_1 _33882_ (.A1(_05729_),
    .A2(_05730_),
    .B1(_05856_),
    .Y(_05857_));
 sky130_fd_sc_hd__and3_2 _33883_ (.A(_05856_),
    .B(_05729_),
    .C(_05730_),
    .X(_05858_));
 sky130_fd_sc_hd__o211a_2 _33884_ (.A1(_05857_),
    .A2(_05858_),
    .B1(_04005_),
    .C1(_04131_),
    .X(_05859_));
 sky130_fd_sc_hd__a21o_1 _33885_ (.A1(_04172_),
    .A2(_04251_),
    .B1(_04248_),
    .X(_05860_));
 sky130_fd_sc_hd__nor2_1 _33886_ (.A(_02275_),
    .B(net340),
    .Y(_05861_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33887_ (.A(_02275_),
    .X(_05862_));
 sky130_fd_sc_hd__buf_1 _33888_ (.A(net340),
    .X(_05863_));
 sky130_fd_sc_hd__nand2_1 _33889_ (.A(_05862_),
    .B(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__nand3b_1 _33890_ (.A_N(_05861_),
    .B(_05864_),
    .C(_04143_),
    .Y(_05866_));
 sky130_fd_sc_hd__buf_2 _33891_ (.A(_00474_),
    .X(_05867_));
 sky130_fd_sc_hd__clkbuf_2 _33892_ (.A(\delay_line[25][13] ),
    .X(_05868_));
 sky130_fd_sc_hd__and2_1 _33893_ (.A(_02275_),
    .B(net340),
    .X(_05869_));
 sky130_fd_sc_hd__o2bb2ai_2 _33894_ (.A1_N(_05867_),
    .A2_N(_05868_),
    .B1(_05861_),
    .B2(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__clkbuf_2 _33895_ (.A(_22819_),
    .X(_05871_));
 sky130_fd_sc_hd__a21o_1 _33896_ (.A1(_05866_),
    .A2(_05870_),
    .B1(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__nand3_2 _33897_ (.A(_05870_),
    .B(_05871_),
    .C(_05866_),
    .Y(_05873_));
 sky130_fd_sc_hd__and3_1 _33898_ (.A(_24511_),
    .B(_05862_),
    .C(_04144_),
    .X(_05874_));
 sky130_fd_sc_hd__a21o_1 _33899_ (.A1(_21570_),
    .A2(_04146_),
    .B1(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__nand3_1 _33900_ (.A(_05872_),
    .B(_05873_),
    .C(_05875_),
    .Y(_05877_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33901_ (.A(_21570_),
    .X(_05878_));
 sky130_fd_sc_hd__a221o_2 _33902_ (.A1(_05878_),
    .A2(_04146_),
    .B1(_05872_),
    .B2(_05873_),
    .C1(_05874_),
    .X(_05879_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33903_ (.A(_21565_),
    .X(_05880_));
 sky130_fd_sc_hd__and2b_1 _33904_ (.A_N(_00484_),
    .B(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__a31o_1 _33905_ (.A1(_20484_),
    .A2(_20485_),
    .A3(_00484_),
    .B1(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__a21o_1 _33906_ (.A1(_05877_),
    .A2(_05879_),
    .B1(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__nand3_1 _33907_ (.A(_05877_),
    .B(_05879_),
    .C(_05882_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand2_1 _33908_ (.A(_04150_),
    .B(_04154_),
    .Y(_05885_));
 sky130_fd_sc_hd__a21oi_1 _33909_ (.A1(_05883_),
    .A2(_05884_),
    .B1(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33910_ (.A(_00484_),
    .X(_05888_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _33911_ (.A(_24507_),
    .X(_05889_));
 sky130_fd_sc_hd__nand3b_2 _33912_ (.A_N(_05888_),
    .B(_05889_),
    .C(_17215_),
    .Y(_05890_));
 sky130_fd_sc_hd__nand2_1 _33913_ (.A(_05890_),
    .B(_05889_),
    .Y(_05891_));
 sky130_fd_sc_hd__and3_1 _33914_ (.A(_05885_),
    .B(_05883_),
    .C(_05884_),
    .X(_05892_));
 sky130_fd_sc_hd__nor3_1 _33915_ (.A(_05886_),
    .B(_05891_),
    .C(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__o2bb2a_1 _33916_ (.A1_N(_05890_),
    .A2_N(_05889_),
    .B1(_05886_),
    .B2(_05892_),
    .X(_05894_));
 sky130_fd_sc_hd__o211a_1 _33917_ (.A1(_05893_),
    .A2(_05894_),
    .B1(_04159_),
    .C1(_04160_),
    .X(_05895_));
 sky130_fd_sc_hd__a211o_1 _33918_ (.A1(_04159_),
    .A2(_04160_),
    .B1(_05893_),
    .C1(_05894_),
    .X(_05896_));
 sky130_fd_sc_hd__and2b_1 _33919_ (.A_N(_05895_),
    .B(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__xnor2_1 _33920_ (.A(_04158_),
    .B(_05897_),
    .Y(_05899_));
 sky130_fd_sc_hd__nor3_1 _33921_ (.A(_04164_),
    .B(_04166_),
    .C(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__o211ai_1 _33922_ (.A1(_04166_),
    .A2(_04167_),
    .B1(_02305_),
    .C1(_04168_),
    .Y(_05901_));
 sky130_fd_sc_hd__a21oi_1 _33923_ (.A1(_04141_),
    .A2(_05901_),
    .B1(_04170_),
    .Y(_05902_));
 sky130_fd_sc_hd__o21a_1 _33924_ (.A1(_04164_),
    .A2(_04166_),
    .B1(_05899_),
    .X(_05903_));
 sky130_fd_sc_hd__o21ai_1 _33925_ (.A1(_05900_),
    .A2(_05903_),
    .B1(_05902_),
    .Y(_05904_));
 sky130_fd_sc_hd__o21a_2 _33926_ (.A1(_05900_),
    .A2(_05902_),
    .B1(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__inv_2 _33927_ (.A(_04198_),
    .Y(_05906_));
 sky130_fd_sc_hd__nor2_1 _33928_ (.A(_05906_),
    .B(_04197_),
    .Y(_05907_));
 sky130_fd_sc_hd__a21o_1 _33929_ (.A1(_04174_),
    .A2(_06876_),
    .B1(_17095_),
    .X(_05908_));
 sky130_fd_sc_hd__a21oi_1 _33930_ (.A1(_04174_),
    .A2(_00512_),
    .B1(_20450_),
    .Y(_05910_));
 sky130_fd_sc_hd__and3_1 _33931_ (.A(_02371_),
    .B(_19501_),
    .C(_20449_),
    .X(_05911_));
 sky130_fd_sc_hd__nor2_1 _33932_ (.A(_05910_),
    .B(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__nor2_1 _33933_ (.A(_24555_),
    .B(\delay_line[22][13] ),
    .Y(_05913_));
 sky130_fd_sc_hd__nand2_1 _33934_ (.A(_24555_),
    .B(\delay_line[22][13] ),
    .Y(_05914_));
 sky130_fd_sc_hd__nand3b_1 _33935_ (.A_N(_05913_),
    .B(_04182_),
    .C(_05914_),
    .Y(_05915_));
 sky130_fd_sc_hd__and2_1 _33936_ (.A(_24555_),
    .B(\delay_line[22][13] ),
    .X(_05916_));
 sky130_fd_sc_hd__o21ai_1 _33937_ (.A1(_05916_),
    .A2(_05913_),
    .B1(_04180_),
    .Y(_05917_));
 sky130_fd_sc_hd__nand3_2 _33938_ (.A(_05912_),
    .B(_05915_),
    .C(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__a2bb2o_1 _33939_ (.A1_N(_05910_),
    .A2_N(_05911_),
    .B1(_05915_),
    .B2(_05917_),
    .X(_05919_));
 sky130_fd_sc_hd__nand2_1 _33940_ (.A(_04181_),
    .B(_04185_),
    .Y(_05921_));
 sky130_fd_sc_hd__a21o_1 _33941_ (.A1(_05918_),
    .A2(_05919_),
    .B1(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__or3_1 _33942_ (.A(_19502_),
    .B(_04174_),
    .C(_17084_),
    .X(_05923_));
 sky130_fd_sc_hd__nand3_2 _33943_ (.A(_05921_),
    .B(_05918_),
    .C(_05919_),
    .Y(_05924_));
 sky130_fd_sc_hd__and4_1 _33944_ (.A(_05922_),
    .B(_18317_),
    .C(_05923_),
    .D(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__a22oi_1 _33945_ (.A1(_18317_),
    .A2(_05923_),
    .B1(_05922_),
    .B2(_05924_),
    .Y(_05926_));
 sky130_fd_sc_hd__o221ai_1 _33946_ (.A1(_05908_),
    .A2(_04190_),
    .B1(_05925_),
    .B2(_05926_),
    .C1(_04189_),
    .Y(_05927_));
 sky130_fd_sc_hd__o21ai_1 _33947_ (.A1(_05908_),
    .A2(_04190_),
    .B1(_04189_),
    .Y(_05928_));
 sky130_fd_sc_hd__nor2_1 _33948_ (.A(_05925_),
    .B(_05926_),
    .Y(_05929_));
 sky130_fd_sc_hd__nand2_1 _33949_ (.A(_05928_),
    .B(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__nand2_1 _33950_ (.A(_05927_),
    .B(_05930_),
    .Y(_05932_));
 sky130_fd_sc_hd__xor2_1 _33951_ (.A(_04192_),
    .B(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__xor2_1 _33952_ (.A(_05907_),
    .B(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__a21boi_1 _33953_ (.A1(_04202_),
    .A2(_04200_),
    .B1_N(_04201_),
    .Y(_05935_));
 sky130_fd_sc_hd__xor2_1 _33954_ (.A(_05934_),
    .B(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__nand2_1 _33955_ (.A(_04237_),
    .B(_04238_),
    .Y(_05937_));
 sky130_fd_sc_hd__or3_1 _33956_ (.A(_22876_),
    .B(_22871_),
    .C(_02318_),
    .X(_05938_));
 sky130_fd_sc_hd__o21ai_1 _33957_ (.A1(_22871_),
    .A2(_02318_),
    .B1(_22876_),
    .Y(_05939_));
 sky130_fd_sc_hd__inv_2 _33958_ (.A(_04218_),
    .Y(_05940_));
 sky130_fd_sc_hd__o21ai_2 _33959_ (.A1(_24579_),
    .A2(_00559_),
    .B1(_22883_),
    .Y(_05941_));
 sky130_fd_sc_hd__a21o_1 _33960_ (.A1(_24583_),
    .A2(_00551_),
    .B1(_05941_),
    .X(_05943_));
 sky130_fd_sc_hd__and2_1 _33961_ (.A(\delay_line[24][9] ),
    .B(\delay_line[24][10] ),
    .X(_05944_));
 sky130_fd_sc_hd__nor2_1 _33962_ (.A(_24579_),
    .B(_00559_),
    .Y(_05945_));
 sky130_fd_sc_hd__o21bai_2 _33963_ (.A1(_05944_),
    .A2(_05945_),
    .B1_N(_22884_),
    .Y(_05946_));
 sky130_fd_sc_hd__buf_1 _33964_ (.A(\delay_line[24][13] ),
    .X(_05947_));
 sky130_fd_sc_hd__clkbuf_2 _33965_ (.A(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__a21o_1 _33966_ (.A1(_05943_),
    .A2(_05946_),
    .B1(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__and3_1 _33967_ (.A(_04212_),
    .B(_04214_),
    .C(_04209_),
    .X(_05950_));
 sky130_fd_sc_hd__o211ai_1 _33968_ (.A1(_05944_),
    .A2(_05941_),
    .B1(_05948_),
    .C1(_05946_),
    .Y(_05951_));
 sky130_fd_sc_hd__nand3_2 _33969_ (.A(_05949_),
    .B(_05950_),
    .C(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__o211a_1 _33970_ (.A1(_05944_),
    .A2(_05941_),
    .B1(_05948_),
    .C1(_05946_),
    .X(_05954_));
 sky130_fd_sc_hd__a21oi_1 _33971_ (.A1(_05943_),
    .A2(_05946_),
    .B1(_05948_),
    .Y(_05955_));
 sky130_fd_sc_hd__o21ai_2 _33972_ (.A1(_05954_),
    .A2(_05955_),
    .B1(_04216_),
    .Y(_05956_));
 sky130_fd_sc_hd__clkbuf_2 _33973_ (.A(_24583_),
    .X(_05957_));
 sky130_fd_sc_hd__o21ai_2 _33974_ (.A1(_22891_),
    .A2(_05957_),
    .B1(_21628_),
    .Y(_05958_));
 sky130_fd_sc_hd__o21a_1 _33975_ (.A1(_21628_),
    .A2(_04210_),
    .B1(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__a21o_1 _33976_ (.A1(_05952_),
    .A2(_05956_),
    .B1(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__clkbuf_2 _33977_ (.A(_21628_),
    .X(_05961_));
 sky130_fd_sc_hd__o2111ai_4 _33978_ (.A1(_05961_),
    .A2(_04210_),
    .B1(_05952_),
    .C1(_05956_),
    .D1(_05958_),
    .Y(_05962_));
 sky130_fd_sc_hd__o211ai_4 _33979_ (.A1(_05940_),
    .A2(_04222_),
    .B1(_05960_),
    .C1(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__a211o_1 _33980_ (.A1(_05960_),
    .A2(_05962_),
    .B1(_05940_),
    .C1(_04222_),
    .X(_05965_));
 sky130_fd_sc_hd__nand4_2 _33981_ (.A(_05938_),
    .B(_05939_),
    .C(_05963_),
    .D(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__a22o_1 _33982_ (.A1(_05938_),
    .A2(_05939_),
    .B1(_05963_),
    .B2(_05965_),
    .X(_05967_));
 sky130_fd_sc_hd__nand2_1 _33983_ (.A(_04232_),
    .B(_04233_),
    .Y(_05968_));
 sky130_fd_sc_hd__a21oi_1 _33984_ (.A1(_05966_),
    .A2(_05967_),
    .B1(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand3_1 _33985_ (.A(_05968_),
    .B(_05966_),
    .C(_05967_),
    .Y(_05970_));
 sky130_fd_sc_hd__nand3b_1 _33986_ (.A_N(_05969_),
    .B(_05970_),
    .C(_04226_),
    .Y(_05971_));
 sky130_fd_sc_hd__and3_1 _33987_ (.A(_05968_),
    .B(_05966_),
    .C(_05967_),
    .X(_05972_));
 sky130_fd_sc_hd__o21bai_1 _33988_ (.A1(_05969_),
    .A2(_05972_),
    .B1_N(_04226_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand2_1 _33989_ (.A(_05971_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__xnor2_1 _33990_ (.A(_05937_),
    .B(_05974_),
    .Y(_05976_));
 sky130_fd_sc_hd__o21bai_2 _33991_ (.A1(_04242_),
    .A2(_04205_),
    .B1_N(_04243_),
    .Y(_05977_));
 sky130_fd_sc_hd__xor2_1 _33992_ (.A(_05976_),
    .B(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__nand2_1 _33993_ (.A(_05936_),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__or2_1 _33994_ (.A(_05936_),
    .B(_05978_),
    .X(_05980_));
 sky130_fd_sc_hd__nand2_1 _33995_ (.A(_05979_),
    .B(_05980_),
    .Y(_05981_));
 sky130_fd_sc_hd__xor2_2 _33996_ (.A(_05905_),
    .B(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__and3_1 _33997_ (.A(_05982_),
    .B(_04130_),
    .C(_04084_),
    .X(_05983_));
 sky130_fd_sc_hd__a21oi_1 _33998_ (.A1(_04084_),
    .A2(_04130_),
    .B1(_05982_),
    .Y(_05984_));
 sky130_fd_sc_hd__nor2_1 _33999_ (.A(_05983_),
    .B(_05984_),
    .Y(_05985_));
 sky130_fd_sc_hd__xnor2_2 _34000_ (.A(_05860_),
    .B(_05985_),
    .Y(_05987_));
 sky130_fd_sc_hd__a211o_2 _34001_ (.A1(_04005_),
    .A2(_04131_),
    .B1(_05857_),
    .C1(_05858_),
    .X(_05988_));
 sky130_fd_sc_hd__o21ai_2 _34002_ (.A1(_05987_),
    .A2(_05859_),
    .B1(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__nor2_1 _34003_ (.A(_05987_),
    .B(_05859_),
    .Y(_05990_));
 sky130_fd_sc_hd__a21o_1 _34004_ (.A1(_05990_),
    .A2(_05988_),
    .B1(_05987_),
    .X(_05991_));
 sky130_fd_sc_hd__o21a_1 _34005_ (.A1(_05859_),
    .A2(_05989_),
    .B1(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__xor2_1 _34006_ (.A(_05592_),
    .B(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__nand2_1 _34007_ (.A(_05591_),
    .B(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__or2_1 _34008_ (.A(_05591_),
    .B(_05993_),
    .X(_05995_));
 sky130_fd_sc_hd__nand2_1 _34009_ (.A(_05994_),
    .B(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__a21o_1 _34010_ (.A1(_04263_),
    .A2(_04439_),
    .B1(_05996_),
    .X(_05998_));
 sky130_fd_sc_hd__o211ai_1 _34011_ (.A1(_04260_),
    .A2(_04259_),
    .B1(_04439_),
    .C1(_05996_),
    .Y(_05999_));
 sky130_fd_sc_hd__nand2_1 _34012_ (.A(_05998_),
    .B(_05999_),
    .Y(_06000_));
 sky130_fd_sc_hd__or3_2 _34013_ (.A(_05405_),
    .B(_05407_),
    .C(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__o21ai_1 _34014_ (.A1(_05405_),
    .A2(_05407_),
    .B1(_06000_),
    .Y(_06002_));
 sky130_fd_sc_hd__o32ai_2 _34015_ (.A1(_03868_),
    .A2(_03869_),
    .A3(_04441_),
    .B1(_04440_),
    .B2(_03871_),
    .Y(_06003_));
 sky130_fd_sc_hd__a21oi_1 _34016_ (.A1(_06001_),
    .A2(_06002_),
    .B1(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__and3_2 _34017_ (.A(_06003_),
    .B(_06001_),
    .C(_06002_),
    .X(_06005_));
 sky130_fd_sc_hd__nor2_1 _34018_ (.A(_06004_),
    .B(_06005_),
    .Y(_06006_));
 sky130_fd_sc_hd__nand3_2 _34019_ (.A(_05155_),
    .B(_05158_),
    .C(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__inv_2 _34020_ (.A(_06007_),
    .Y(_06009_));
 sky130_fd_sc_hd__o31a_1 _34021_ (.A1(_03868_),
    .A2(_03869_),
    .A3(_04441_),
    .B1(_04442_),
    .X(_06010_));
 sky130_fd_sc_hd__a2bb2o_1 _34022_ (.A1_N(_03617_),
    .A2_N(_04456_),
    .B1(_03619_),
    .B2(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__a21boi_1 _34023_ (.A1(_05157_),
    .A2(_05153_),
    .B1_N(_05154_),
    .Y(_06012_));
 sky130_fd_sc_hd__o211a_1 _34024_ (.A1(_03603_),
    .A2(_05156_),
    .B1(_05157_),
    .C1(_05153_),
    .X(_06013_));
 sky130_fd_sc_hd__o21bai_2 _34025_ (.A1(_06012_),
    .A2(_06013_),
    .B1_N(_06006_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_1 _34026_ (.A(_06011_),
    .B(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__a21o_1 _34027_ (.A1(_06014_),
    .A2(_06007_),
    .B1(_06011_),
    .X(_06016_));
 sky130_fd_sc_hd__o221ai_4 _34028_ (.A1(_04595_),
    .A2(_04596_),
    .B1(_06009_),
    .B2(_06015_),
    .C1(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__a21oi_1 _34029_ (.A1(_06014_),
    .A2(_06007_),
    .B1(_06011_),
    .Y(_06018_));
 sky130_fd_sc_hd__and3_1 _34030_ (.A(_06011_),
    .B(_06014_),
    .C(_06007_),
    .X(_06020_));
 sky130_fd_sc_hd__nor2_1 _34031_ (.A(_04595_),
    .B(_04596_),
    .Y(_06021_));
 sky130_fd_sc_hd__o21ai_1 _34032_ (.A1(_06018_),
    .A2(_06020_),
    .B1(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__nand3_1 _34033_ (.A(_04522_),
    .B(_06017_),
    .C(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__a21o_1 _34034_ (.A1(_06017_),
    .A2(_06022_),
    .B1(_04522_),
    .X(_06024_));
 sky130_fd_sc_hd__nand2_1 _34035_ (.A(_11328_),
    .B(_25159_),
    .Y(_06025_));
 sky130_fd_sc_hd__xor2_2 _34036_ (.A(_25238_),
    .B(_18727_),
    .X(_06026_));
 sky130_fd_sc_hd__nand3_4 _34037_ (.A(_18824_),
    .B(_06025_),
    .C(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__a21o_2 _34038_ (.A1(_18824_),
    .A2(_06025_),
    .B1(_06026_),
    .X(_06028_));
 sky130_fd_sc_hd__and3_2 _34039_ (.A(_02998_),
    .B(_04473_),
    .C(_25240_),
    .X(_06029_));
 sky130_fd_sc_hd__a21oi_2 _34040_ (.A1(_18799_),
    .A2(_19813_),
    .B1(_02997_),
    .Y(_06031_));
 sky130_fd_sc_hd__a211oi_4 _34041_ (.A1(_06027_),
    .A2(_06028_),
    .B1(_06029_),
    .C1(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__o211ai_4 _34042_ (.A1(_06031_),
    .A2(_06029_),
    .B1(_06028_),
    .C1(_06027_),
    .Y(_06033_));
 sky130_fd_sc_hd__inv_2 _34043_ (.A(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__o21ai_2 _34044_ (.A1(_06032_),
    .A2(_06034_),
    .B1(_04477_),
    .Y(_06035_));
 sky130_fd_sc_hd__or3_2 _34045_ (.A(_04477_),
    .B(_06032_),
    .C(_06034_),
    .X(_06036_));
 sky130_fd_sc_hd__a221oi_4 _34046_ (.A1(_06035_),
    .A2(_06036_),
    .B1(_03025_),
    .B2(_03000_),
    .C1(_03024_),
    .Y(_06037_));
 sky130_fd_sc_hd__o211a_2 _34047_ (.A1(_03024_),
    .A2(_03027_),
    .B1(_06035_),
    .C1(_06036_),
    .X(_06038_));
 sky130_fd_sc_hd__or3b_4 _34048_ (.A(_04480_),
    .B(_04475_),
    .C_N(_02954_),
    .X(_06039_));
 sky130_fd_sc_hd__o211ai_2 _34049_ (.A1(_06037_),
    .A2(_06038_),
    .B1(_04478_),
    .C1(_06039_),
    .Y(_06040_));
 sky130_fd_sc_hd__inv_2 _34050_ (.A(_06040_),
    .Y(_06042_));
 sky130_fd_sc_hd__a211oi_4 _34051_ (.A1(_04478_),
    .A2(_06039_),
    .B1(_06037_),
    .C1(_06038_),
    .Y(_06043_));
 sky130_fd_sc_hd__a21oi_4 _34052_ (.A1(_04467_),
    .A2(_04483_),
    .B1(_04486_),
    .Y(_06044_));
 sky130_fd_sc_hd__o21a_1 _34053_ (.A1(_06042_),
    .A2(_06043_),
    .B1(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__nor3_1 _34054_ (.A(_06044_),
    .B(_06042_),
    .C(_06043_),
    .Y(_06046_));
 sky130_fd_sc_hd__nor2_1 _34055_ (.A(_06045_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__o21a_1 _34056_ (.A1(_02933_),
    .A2(_02994_),
    .B1(_03058_),
    .X(_06048_));
 sky130_fd_sc_hd__a211oi_1 _34057_ (.A1(_03060_),
    .A2(_03063_),
    .B1(_06047_),
    .C1(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__o21ai_2 _34058_ (.A1(_06048_),
    .A2(_03065_),
    .B1(_06047_),
    .Y(_06050_));
 sky130_fd_sc_hd__or2b_1 _34059_ (.A(_06049_),
    .B_N(_06050_),
    .X(_06051_));
 sky130_fd_sc_hd__xor2_2 _34060_ (.A(_04489_),
    .B(_06051_),
    .X(_06053_));
 sky130_fd_sc_hd__a21bo_1 _34061_ (.A1(_06023_),
    .A2(_06024_),
    .B1_N(_06053_),
    .X(_06054_));
 sky130_fd_sc_hd__nand3b_1 _34062_ (.A_N(_06053_),
    .B(_06023_),
    .C(_06024_),
    .Y(_06055_));
 sky130_fd_sc_hd__a31o_1 _34063_ (.A1(_02993_),
    .A2(_04458_),
    .A3(_04464_),
    .B1(_04499_),
    .X(_06056_));
 sky130_fd_sc_hd__a21oi_1 _34064_ (.A1(_06054_),
    .A2(_06055_),
    .B1(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__nand3_1 _34065_ (.A(_06056_),
    .B(_06054_),
    .C(_06055_),
    .Y(_06058_));
 sky130_fd_sc_hd__o21a_1 _34066_ (.A1(_02970_),
    .A2(_04491_),
    .B1(_04493_),
    .X(_06059_));
 sky130_fd_sc_hd__nand3b_1 _34067_ (.A_N(_06057_),
    .B(_06058_),
    .C(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__inv_2 _34068_ (.A(_06058_),
    .Y(_06061_));
 sky130_fd_sc_hd__o21ai_1 _34069_ (.A1(_02970_),
    .A2(_04491_),
    .B1(_04493_),
    .Y(_06062_));
 sky130_fd_sc_hd__o21ai_1 _34070_ (.A1(_06057_),
    .A2(_06061_),
    .B1(_06062_),
    .Y(_06064_));
 sky130_fd_sc_hd__o21ai_1 _34071_ (.A1(_04507_),
    .A2(_04504_),
    .B1(_04510_),
    .Y(_06065_));
 sky130_fd_sc_hd__a21o_1 _34072_ (.A1(_06060_),
    .A2(_06064_),
    .B1(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__nand3_2 _34073_ (.A(_06065_),
    .B(_06060_),
    .C(_06064_),
    .Y(_06067_));
 sky130_fd_sc_hd__a21o_1 _34074_ (.A1(_02982_),
    .A2(_04513_),
    .B1(_04508_),
    .X(_06068_));
 sky130_fd_sc_hd__o22ai_1 _34075_ (.A1(_04512_),
    .A2(_06068_),
    .B1(_04519_),
    .B2(_04521_),
    .Y(_06069_));
 sky130_fd_sc_hd__a21boi_1 _34076_ (.A1(_06066_),
    .A2(_06067_),
    .B1_N(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__o2111ai_1 _34077_ (.A1(_04521_),
    .A2(_04519_),
    .B1(_04518_),
    .C1(_06067_),
    .D1(_06066_),
    .Y(_06071_));
 sky130_fd_sc_hd__or2b_2 _34078_ (.A(_06070_),
    .B_N(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__clkbuf_1 _34079_ (.A(_06072_),
    .X(_00008_));
 sky130_fd_sc_hd__a211o_1 _34080_ (.A1(_02965_),
    .A2(_02967_),
    .B1(_04487_),
    .C1(_06051_),
    .X(_06074_));
 sky130_fd_sc_hd__a21oi_1 _34081_ (.A1(_06017_),
    .A2(_06022_),
    .B1(_04522_),
    .Y(_06075_));
 sky130_fd_sc_hd__o22ai_2 _34082_ (.A1(_06015_),
    .A2(_06009_),
    .B1(_06018_),
    .B2(_06021_),
    .Y(_06076_));
 sky130_fd_sc_hd__o31a_4 _34083_ (.A1(_05159_),
    .A2(_05400_),
    .A3(_05401_),
    .B1(_05406_),
    .X(_06077_));
 sky130_fd_sc_hd__inv_2 _34084_ (.A(_05111_),
    .Y(_06078_));
 sky130_fd_sc_hd__xor2_1 _34085_ (.A(_03115_),
    .B(_05061_),
    .X(_06079_));
 sky130_fd_sc_hd__nor2_1 _34086_ (.A(_06079_),
    .B(_05016_),
    .Y(_06080_));
 sky130_fd_sc_hd__o21ai_4 _34087_ (.A1(_05000_),
    .A2(_04968_),
    .B1(_05001_),
    .Y(_06081_));
 sky130_fd_sc_hd__nand2_1 _34088_ (.A(_04889_),
    .B(_04679_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand2_2 _34089_ (.A(_04680_),
    .B(_06082_),
    .Y(_06083_));
 sky130_fd_sc_hd__nand3_1 _34090_ (.A(_04653_),
    .B(_04654_),
    .C(_04657_),
    .Y(_06085_));
 sky130_fd_sc_hd__nand2_1 _34091_ (.A(_06085_),
    .B(_04671_),
    .Y(_06086_));
 sky130_fd_sc_hd__o21ba_1 _34092_ (.A1(_04668_),
    .A2(_04666_),
    .B1_N(_04665_),
    .X(_06087_));
 sky130_fd_sc_hd__buf_1 _34093_ (.A(\delay_line[6][15] ),
    .X(_06088_));
 sky130_fd_sc_hd__or2b_2 _34094_ (.A(_00261_),
    .B_N(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__inv_2 _34095_ (.A(\delay_line[6][15] ),
    .Y(_06090_));
 sky130_fd_sc_hd__clkbuf_2 _34096_ (.A(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__nand2_1 _34097_ (.A(_06091_),
    .B(_00265_),
    .Y(_06092_));
 sky130_fd_sc_hd__o21a_1 _34098_ (.A1(_22525_),
    .A2(_24091_),
    .B1(_21862_),
    .X(_06093_));
 sky130_fd_sc_hd__a221o_1 _34099_ (.A1(_03413_),
    .A2(_24091_),
    .B1(_06089_),
    .B2(_06092_),
    .C1(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__o211ai_4 _34100_ (.A1(_04974_),
    .A2(_06093_),
    .B1(_06089_),
    .C1(_06092_),
    .Y(_06096_));
 sky130_fd_sc_hd__clkbuf_2 _34101_ (.A(_04978_),
    .X(_06097_));
 sky130_fd_sc_hd__and4b_1 _34102_ (.A_N(_01915_),
    .B(_06094_),
    .C(_06096_),
    .D(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__o2bb2a_1 _34103_ (.A1_N(_06094_),
    .A2_N(_06096_),
    .B1(_01915_),
    .B2(_04980_),
    .X(_06099_));
 sky130_fd_sc_hd__nor2_1 _34104_ (.A(_01909_),
    .B(_01747_),
    .Y(_06100_));
 sky130_fd_sc_hd__and2_1 _34105_ (.A(_04973_),
    .B(\delay_line[7][11] ),
    .X(_06101_));
 sky130_fd_sc_hd__o21bai_1 _34106_ (.A1(_06100_),
    .A2(_06101_),
    .B1_N(_04971_),
    .Y(_06102_));
 sky130_fd_sc_hd__or3b_1 _34107_ (.A(_06100_),
    .B(_06101_),
    .C_N(_04971_),
    .X(_06103_));
 sky130_fd_sc_hd__nand2_1 _34108_ (.A(_06102_),
    .B(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__o21a_1 _34109_ (.A1(_06098_),
    .A2(_06099_),
    .B1(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__nor2_1 _34110_ (.A(_06087_),
    .B(_06105_),
    .Y(_06107_));
 sky130_fd_sc_hd__or3_1 _34111_ (.A(_06104_),
    .B(_06099_),
    .C(_06098_),
    .X(_06108_));
 sky130_fd_sc_hd__and4bb_1 _34112_ (.A_N(_06098_),
    .B_N(_06099_),
    .C(_06102_),
    .D(_06103_),
    .X(_06109_));
 sky130_fd_sc_hd__o21a_1 _34113_ (.A1(_06105_),
    .A2(_06109_),
    .B1(_06087_),
    .X(_06110_));
 sky130_fd_sc_hd__a21oi_1 _34114_ (.A1(_06107_),
    .A2(_06108_),
    .B1(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__xor2_1 _34115_ (.A(_04988_),
    .B(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__xnor2_1 _34116_ (.A(_06086_),
    .B(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__o21ba_1 _34117_ (.A1(_03428_),
    .A2(_04990_),
    .B1_N(_04991_),
    .X(_06114_));
 sky130_fd_sc_hd__or2b_1 _34118_ (.A(_06113_),
    .B_N(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__or2b_2 _34119_ (.A(_06114_),
    .B_N(_06113_),
    .X(_06116_));
 sky130_fd_sc_hd__o21bai_2 _34120_ (.A1(_04969_),
    .A2(_04995_),
    .B1_N(_04994_),
    .Y(_06118_));
 sky130_fd_sc_hd__a21oi_1 _34121_ (.A1(_06115_),
    .A2(_06116_),
    .B1(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__inv_2 _34122_ (.A(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__nand3_4 _34123_ (.A(_06118_),
    .B(_06115_),
    .C(_06116_),
    .Y(_06121_));
 sky130_fd_sc_hd__and4bb_1 _34124_ (.A_N(_03455_),
    .B_N(_03456_),
    .C(_04916_),
    .D(_03457_),
    .X(_06122_));
 sky130_fd_sc_hd__o21a_1 _34125_ (.A1(_04907_),
    .A2(_03489_),
    .B1(_04917_),
    .X(_06123_));
 sky130_fd_sc_hd__and3_1 _34126_ (.A(_03455_),
    .B(_04910_),
    .C(_04911_),
    .X(_06124_));
 sky130_fd_sc_hd__buf_1 _34127_ (.A(net438),
    .X(_06125_));
 sky130_fd_sc_hd__or2b_1 _34128_ (.A(\delay_line[3][13] ),
    .B_N(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__or2b_1 _34129_ (.A(net438),
    .B_N(_03454_),
    .X(_06127_));
 sky130_fd_sc_hd__nand4_2 _34130_ (.A(_04940_),
    .B(_06126_),
    .C(_06127_),
    .D(_04941_),
    .Y(_06129_));
 sky130_fd_sc_hd__a22o_1 _34131_ (.A1(_04940_),
    .A2(net435),
    .B1(_06126_),
    .B2(_06127_),
    .X(_06130_));
 sky130_fd_sc_hd__and2b_1 _34132_ (.A_N(_01861_),
    .B(_04908_),
    .X(_06131_));
 sky130_fd_sc_hd__a21o_1 _34133_ (.A1(_06129_),
    .A2(_06130_),
    .B1(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__nand3_2 _34134_ (.A(_06130_),
    .B(_06131_),
    .C(_06129_),
    .Y(_06133_));
 sky130_fd_sc_hd__nand3_1 _34135_ (.A(_06132_),
    .B(_04947_),
    .C(_06133_),
    .Y(_06134_));
 sky130_fd_sc_hd__a32o_1 _34136_ (.A1(_04945_),
    .A2(_04943_),
    .A3(_04944_),
    .B1(_06133_),
    .B2(_06132_),
    .X(_06135_));
 sky130_fd_sc_hd__o211ai_2 _34137_ (.A1(_06124_),
    .A2(_04914_),
    .B1(_06134_),
    .C1(_06135_),
    .Y(_06136_));
 sky130_fd_sc_hd__a211o_1 _34138_ (.A1(_06134_),
    .A2(_06135_),
    .B1(_06124_),
    .C1(_04914_),
    .X(_06137_));
 sky130_fd_sc_hd__o31ai_1 _34139_ (.A1(_04946_),
    .A2(_04947_),
    .A3(_04961_),
    .B1(_04958_),
    .Y(_06138_));
 sky130_fd_sc_hd__a21oi_1 _34140_ (.A1(_06136_),
    .A2(_06137_),
    .B1(_06138_),
    .Y(_06140_));
 sky130_fd_sc_hd__and3_1 _34141_ (.A(_06138_),
    .B(_06136_),
    .C(_06137_),
    .X(_06141_));
 sky130_fd_sc_hd__nor2_1 _34142_ (.A(_06140_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__or3_1 _34143_ (.A(_06122_),
    .B(_06123_),
    .C(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__inv_2 _34144_ (.A(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__o21a_1 _34145_ (.A1(_06122_),
    .A2(_06123_),
    .B1(_06142_),
    .X(_06145_));
 sky130_fd_sc_hd__or2b_1 _34146_ (.A(\delay_line[5][9] ),
    .B_N(\delay_line[3][15] ),
    .X(_06146_));
 sky130_fd_sc_hd__inv_2 _34147_ (.A(\delay_line[3][15] ),
    .Y(_06147_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34148_ (.A(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__nand2_1 _34149_ (.A(_06148_),
    .B(_24040_),
    .Y(_06149_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34150_ (.A(_04952_),
    .X(_06151_));
 sky130_fd_sc_hd__a21o_1 _34151_ (.A1(_06146_),
    .A2(_06149_),
    .B1(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__nand3_2 _34152_ (.A(_06149_),
    .B(_04952_),
    .C(_06146_),
    .Y(_06153_));
 sky130_fd_sc_hd__or2b_1 _34153_ (.A(_22606_),
    .B_N(\delay_line[5][15] ),
    .X(_06154_));
 sky130_fd_sc_hd__or2b_1 _34154_ (.A(\delay_line[5][15] ),
    .B_N(_22606_),
    .X(_06155_));
 sky130_fd_sc_hd__nand3_2 _34155_ (.A(_06154_),
    .B(_06155_),
    .C(\delay_line[5][14] ),
    .Y(_06156_));
 sky130_fd_sc_hd__clkbuf_2 _34156_ (.A(\delay_line[5][14] ),
    .X(_06157_));
 sky130_fd_sc_hd__a21o_1 _34157_ (.A1(_06154_),
    .A2(_06155_),
    .B1(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__a21bo_1 _34158_ (.A1(_04952_),
    .A2(_04951_),
    .B1_N(_04950_),
    .X(_06159_));
 sky130_fd_sc_hd__a21oi_1 _34159_ (.A1(_06156_),
    .A2(_06158_),
    .B1(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__inv_2 _34160_ (.A(_06160_),
    .Y(_06162_));
 sky130_fd_sc_hd__nand3_2 _34161_ (.A(_06156_),
    .B(_06158_),
    .C(_06159_),
    .Y(_06163_));
 sky130_fd_sc_hd__nand3_1 _34162_ (.A(_06162_),
    .B(_04956_),
    .C(_06163_),
    .Y(_06164_));
 sky130_fd_sc_hd__a21o_1 _34163_ (.A1(_06163_),
    .A2(_06162_),
    .B1(_04956_),
    .X(_06165_));
 sky130_fd_sc_hd__and4_1 _34164_ (.A(_06152_),
    .B(_06153_),
    .C(_06164_),
    .D(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__a22oi_2 _34165_ (.A1(_06152_),
    .A2(_06153_),
    .B1(_06164_),
    .B2(_06165_),
    .Y(_06167_));
 sky130_fd_sc_hd__buf_1 _34166_ (.A(net426),
    .X(_06168_));
 sky130_fd_sc_hd__o21ba_1 _34167_ (.A1(_01924_),
    .A2(_01920_),
    .B1_N(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__nor3b_1 _34168_ (.A(_01924_),
    .B(_03424_),
    .C_N(_06168_),
    .Y(_06170_));
 sky130_fd_sc_hd__nor2_1 _34169_ (.A(_06169_),
    .B(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__nand3_1 _34170_ (.A(_04984_),
    .B(_04985_),
    .C(_06171_),
    .Y(_06173_));
 sky130_fd_sc_hd__o2bb2ai_1 _34171_ (.A1_N(_04984_),
    .A2_N(_04985_),
    .B1(_06169_),
    .B2(_06170_),
    .Y(_06174_));
 sky130_fd_sc_hd__nand2_1 _34172_ (.A(_06173_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__o21ai_1 _34173_ (.A1(_04933_),
    .A2(_04928_),
    .B1(_03464_),
    .Y(_06176_));
 sky130_fd_sc_hd__xnor2_1 _34174_ (.A(_06175_),
    .B(_06176_),
    .Y(_06177_));
 sky130_fd_sc_hd__a21boi_1 _34175_ (.A1(_04934_),
    .A2(_04935_),
    .B1_N(_04932_),
    .Y(_06178_));
 sky130_fd_sc_hd__xnor2_1 _34176_ (.A(_06177_),
    .B(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__o21a_1 _34177_ (.A1(_06166_),
    .A2(_06167_),
    .B1(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__nor3_1 _34178_ (.A(_06166_),
    .B(_06167_),
    .C(_06179_),
    .Y(_06181_));
 sky130_fd_sc_hd__a211o_1 _34179_ (.A1(_04938_),
    .A2(_04963_),
    .B1(_06180_),
    .C1(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__o211ai_1 _34180_ (.A1(_06180_),
    .A2(_06181_),
    .B1(_04938_),
    .C1(_04963_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand2_1 _34181_ (.A(_06182_),
    .B(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__or3_1 _34182_ (.A(_06144_),
    .B(_06145_),
    .C(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__o21ai_1 _34183_ (.A1(_06144_),
    .A2(_06145_),
    .B1(_06185_),
    .Y(_06187_));
 sky130_fd_sc_hd__and2_1 _34184_ (.A(_06186_),
    .B(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__nand3_2 _34185_ (.A(_06120_),
    .B(_06121_),
    .C(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__a21o_1 _34186_ (.A1(_06120_),
    .A2(_06121_),
    .B1(_06188_),
    .X(_06190_));
 sky130_fd_sc_hd__and3_1 _34187_ (.A(_06083_),
    .B(_06189_),
    .C(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__a21oi_1 _34188_ (.A1(_06189_),
    .A2(_06190_),
    .B1(_06083_),
    .Y(_06192_));
 sky130_fd_sc_hd__nor2_2 _34189_ (.A(_06191_),
    .B(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__xor2_4 _34190_ (.A(_06081_),
    .B(_06193_),
    .X(_06195_));
 sky130_fd_sc_hd__inv_2 _34191_ (.A(_06195_),
    .Y(_06196_));
 sky130_fd_sc_hd__a21bo_1 _34192_ (.A1(_04824_),
    .A2(_04823_),
    .B1_N(_04822_),
    .X(_06197_));
 sky130_fd_sc_hd__xor2_2 _34193_ (.A(_04796_),
    .B(net399),
    .X(_06198_));
 sky130_fd_sc_hd__a21o_1 _34194_ (.A1(_03125_),
    .A2(_04796_),
    .B1(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__clkbuf_2 _34195_ (.A(_04798_),
    .X(_06200_));
 sky130_fd_sc_hd__or3_2 _34196_ (.A(net399),
    .B(_04800_),
    .C(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__clkbuf_2 _34197_ (.A(_23795_),
    .X(_06202_));
 sky130_fd_sc_hd__a21o_2 _34198_ (.A1(_06199_),
    .A2(_06201_),
    .B1(_06202_),
    .X(_06203_));
 sky130_fd_sc_hd__o211ai_4 _34199_ (.A1(_04801_),
    .A2(_06198_),
    .B1(_06202_),
    .C1(_06201_),
    .Y(_06204_));
 sky130_fd_sc_hd__nand3_2 _34200_ (.A(_06203_),
    .B(_23812_),
    .C(_06204_),
    .Y(_06206_));
 sky130_fd_sc_hd__a21o_1 _34201_ (.A1(_06204_),
    .A2(_06203_),
    .B1(_23812_),
    .X(_06207_));
 sky130_fd_sc_hd__o211a_1 _34202_ (.A1(net270),
    .A2(_04763_),
    .B1(_06206_),
    .C1(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__a211oi_1 _34203_ (.A1(_06206_),
    .A2(_06207_),
    .B1(net270),
    .C1(_04763_),
    .Y(_06209_));
 sky130_fd_sc_hd__nor3_1 _34204_ (.A(_04807_),
    .B(_06208_),
    .C(_06209_),
    .Y(_06210_));
 sky130_fd_sc_hd__o21a_1 _34205_ (.A1(_06208_),
    .A2(_06209_),
    .B1(_04807_),
    .X(_06211_));
 sky130_fd_sc_hd__o22a_2 _34206_ (.A1(_04735_),
    .A2(_04739_),
    .B1(_04750_),
    .B2(_04747_),
    .X(_06212_));
 sky130_fd_sc_hd__o21a_1 _34207_ (.A1(_04730_),
    .A2(_04741_),
    .B1(_04745_),
    .X(_06213_));
 sky130_fd_sc_hd__o2bb2a_1 _34208_ (.A1_N(_04703_),
    .A2_N(_04705_),
    .B1(_04716_),
    .B2(_04720_),
    .X(_06214_));
 sky130_fd_sc_hd__a31oi_2 _34209_ (.A1(_04723_),
    .A2(_04705_),
    .A3(_04703_),
    .B1(net452),
    .Y(_06215_));
 sky130_fd_sc_hd__or2b_1 _34210_ (.A(_03169_),
    .B_N(\delay_line[4][11] ),
    .X(_06217_));
 sky130_fd_sc_hd__nand2_1 _34211_ (.A(_03162_),
    .B(_04695_),
    .Y(_06218_));
 sky130_fd_sc_hd__xnor2_2 _34212_ (.A(_03160_),
    .B(net433),
    .Y(_06219_));
 sky130_fd_sc_hd__and3_1 _34213_ (.A(_06217_),
    .B(_06218_),
    .C(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__a21oi_2 _34214_ (.A1(_06217_),
    .A2(_06218_),
    .B1(_06219_),
    .Y(_06221_));
 sky130_fd_sc_hd__or2_1 _34215_ (.A(_06220_),
    .B(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__a21o_1 _34216_ (.A1(_03166_),
    .A2(_03168_),
    .B1(_04699_),
    .X(_06223_));
 sky130_fd_sc_hd__o21bai_4 _34217_ (.A1(_03178_),
    .A2(_03179_),
    .B1_N(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__clkbuf_2 _34218_ (.A(\delay_line[4][11] ),
    .X(_06225_));
 sky130_fd_sc_hd__and4bb_1 _34219_ (.A_N(_23827_),
    .B_N(_03163_),
    .C(_03169_),
    .D(_04694_),
    .X(_06226_));
 sky130_fd_sc_hd__o2bb2a_1 _34220_ (.A1_N(_06225_),
    .A2_N(_06226_),
    .B1(_04702_),
    .B2(_04699_),
    .X(_06228_));
 sky130_fd_sc_hd__nand3b_2 _34221_ (.A_N(_06222_),
    .B(_06224_),
    .C(_06228_),
    .Y(_06229_));
 sky130_fd_sc_hd__a2bb2o_1 _34222_ (.A1_N(_04702_),
    .A2_N(_04699_),
    .B1(_06226_),
    .B2(_06225_),
    .X(_06230_));
 sky130_fd_sc_hd__a21oi_2 _34223_ (.A1(_01604_),
    .A2(_03171_),
    .B1(_06223_),
    .Y(_06231_));
 sky130_fd_sc_hd__o22ai_1 _34224_ (.A1(_06220_),
    .A2(_06221_),
    .B1(_06230_),
    .B2(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__buf_2 _34225_ (.A(_01555_),
    .X(_06233_));
 sky130_fd_sc_hd__nand4_4 _34226_ (.A(_06233_),
    .B(_03153_),
    .C(_04713_),
    .D(_21728_),
    .Y(_06234_));
 sky130_fd_sc_hd__xnor2_1 _34227_ (.A(_25433_),
    .B(\delay_line[11][13] ),
    .Y(_06235_));
 sky130_fd_sc_hd__a21oi_1 _34228_ (.A1(_04712_),
    .A2(_04706_),
    .B1(_04710_),
    .Y(_06236_));
 sky130_fd_sc_hd__xor2_1 _34229_ (.A(_06235_),
    .B(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34230_ (.A(_06237_),
    .X(_06239_));
 sky130_fd_sc_hd__a21oi_1 _34231_ (.A1(_04719_),
    .A2(_06234_),
    .B1(_06239_),
    .Y(_06240_));
 sky130_fd_sc_hd__and3_1 _34232_ (.A(_04719_),
    .B(_06234_),
    .C(_06239_),
    .X(_06241_));
 sky130_fd_sc_hd__o2bb2ai_1 _34233_ (.A1_N(_06229_),
    .A2_N(_06232_),
    .B1(_06240_),
    .B2(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__clkbuf_2 _34234_ (.A(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_2 _34235_ (.A(_06232_),
    .X(_06244_));
 sky130_fd_sc_hd__and4_1 _34236_ (.A(_01560_),
    .B(_01562_),
    .C(_03155_),
    .D(_03156_),
    .X(_06245_));
 sky130_fd_sc_hd__a2bb2oi_2 _34237_ (.A1_N(_01563_),
    .A2_N(_04708_),
    .B1(_06245_),
    .B2(_01597_),
    .Y(_06246_));
 sky130_fd_sc_hd__o21ai_1 _34238_ (.A1(_04715_),
    .A2(_06246_),
    .B1(_06234_),
    .Y(_06247_));
 sky130_fd_sc_hd__inv_2 _34239_ (.A(_06239_),
    .Y(_06248_));
 sky130_fd_sc_hd__nand2_1 _34240_ (.A(_06247_),
    .B(_06248_),
    .Y(_06250_));
 sky130_fd_sc_hd__o211ai_2 _34241_ (.A1(_04715_),
    .A2(_06246_),
    .B1(_06234_),
    .C1(_06239_),
    .Y(_06251_));
 sky130_fd_sc_hd__nand4_2 _34242_ (.A(_06229_),
    .B(_06244_),
    .C(_06250_),
    .D(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__clkbuf_2 _34243_ (.A(\delay_line[0][15] ),
    .X(_06253_));
 sky130_fd_sc_hd__a21oi_1 _34244_ (.A1(_06243_),
    .A2(_06252_),
    .B1(_06253_),
    .Y(_06254_));
 sky130_fd_sc_hd__a2bb2oi_4 _34245_ (.A1_N(_06220_),
    .A2_N(_06221_),
    .B1(_06228_),
    .B2(_06224_),
    .Y(_06255_));
 sky130_fd_sc_hd__nand3_1 _34246_ (.A(_06229_),
    .B(_06250_),
    .C(_06251_),
    .Y(_06256_));
 sky130_fd_sc_hd__o211a_1 _34247_ (.A1(_06255_),
    .A2(_06256_),
    .B1(\delay_line[0][15] ),
    .C1(_06242_),
    .X(_06257_));
 sky130_fd_sc_hd__o22ai_2 _34248_ (.A1(_06214_),
    .A2(_06215_),
    .B1(_06254_),
    .B2(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__buf_6 _34249_ (.A(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__inv_2 _34250_ (.A(net452),
    .Y(_06261_));
 sky130_fd_sc_hd__a21oi_1 _34251_ (.A1(_06261_),
    .A2(_04724_),
    .B1(_06214_),
    .Y(_06262_));
 sky130_fd_sc_hd__a21o_1 _34252_ (.A1(_06243_),
    .A2(_06252_),
    .B1(_06253_),
    .X(_06263_));
 sky130_fd_sc_hd__o211ai_2 _34253_ (.A1(_06255_),
    .A2(_06256_),
    .B1(_06253_),
    .C1(_06243_),
    .Y(_06264_));
 sky130_fd_sc_hd__nand3_2 _34254_ (.A(_06262_),
    .B(_06263_),
    .C(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__clkbuf_2 _34255_ (.A(_04729_),
    .X(_06266_));
 sky130_fd_sc_hd__a21oi_1 _34256_ (.A1(_06259_),
    .A2(_06265_),
    .B1(_06266_),
    .Y(_06267_));
 sky130_fd_sc_hd__o311a_2 _34257_ (.A1(_06214_),
    .A2(_06254_),
    .A3(_06257_),
    .B1(_06266_),
    .C1(_06259_),
    .X(_06268_));
 sky130_fd_sc_hd__o22ai_4 _34258_ (.A1(_04743_),
    .A2(_06213_),
    .B1(_06267_),
    .B2(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__a21o_1 _34259_ (.A1(_06258_),
    .A2(_06265_),
    .B1(_04729_),
    .X(_06270_));
 sky130_fd_sc_hd__clkbuf_2 _34260_ (.A(_06261_),
    .X(_06272_));
 sky130_fd_sc_hd__a31oi_2 _34261_ (.A1(_06262_),
    .A2(_06263_),
    .A3(_06264_),
    .B1(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nand2_1 _34262_ (.A(_06273_),
    .B(_06259_),
    .Y(_06274_));
 sky130_fd_sc_hd__o21ai_1 _34263_ (.A1(_04691_),
    .A2(_04743_),
    .B1(_04727_),
    .Y(_06275_));
 sky130_fd_sc_hd__nand3_1 _34264_ (.A(_06270_),
    .B(_06274_),
    .C(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__buf_4 _34265_ (.A(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__or2_1 _34266_ (.A(_01617_),
    .B(\delay_line[13][15] ),
    .X(_06278_));
 sky130_fd_sc_hd__nand2_1 _34267_ (.A(_01617_),
    .B(\delay_line[13][15] ),
    .Y(_06279_));
 sky130_fd_sc_hd__clkbuf_2 _34268_ (.A(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__and3b_1 _34269_ (.A_N(_04772_),
    .B(_06278_),
    .C(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__and2_1 _34270_ (.A(_06278_),
    .B(_06279_),
    .X(_06283_));
 sky130_fd_sc_hd__and3b_1 _34271_ (.A_N(_06283_),
    .B(net395),
    .C(_00077_),
    .X(_06284_));
 sky130_fd_sc_hd__o2bb2ai_4 _34272_ (.A1_N(_06269_),
    .A2_N(_06277_),
    .B1(_06281_),
    .B2(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__nand2_1 _34273_ (.A(_04772_),
    .B(_06283_),
    .Y(_06286_));
 sky130_fd_sc_hd__clkbuf_2 _34274_ (.A(net395),
    .X(_06287_));
 sky130_fd_sc_hd__a22o_1 _34275_ (.A1(_00077_),
    .A2(_06287_),
    .B1(_06278_),
    .B2(_06280_),
    .X(_06288_));
 sky130_fd_sc_hd__nand2_2 _34276_ (.A(_06286_),
    .B(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__nand3_4 _34277_ (.A(_06269_),
    .B(_06277_),
    .C(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__nand3_4 _34278_ (.A(_06212_),
    .B(_06285_),
    .C(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__o22ai_1 _34279_ (.A1(_04736_),
    .A2(_04739_),
    .B1(_04750_),
    .B2(_04747_),
    .Y(_06292_));
 sky130_fd_sc_hd__or2_1 _34280_ (.A(_06281_),
    .B(_06284_),
    .X(_06294_));
 sky130_fd_sc_hd__a21o_1 _34281_ (.A1(_06269_),
    .A2(_06277_),
    .B1(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__nand4_1 _34282_ (.A(_06269_),
    .B(_06277_),
    .C(_06286_),
    .D(_06288_),
    .Y(_06296_));
 sky130_fd_sc_hd__nand3_2 _34283_ (.A(_06292_),
    .B(_06295_),
    .C(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__and4b_2 _34284_ (.A_N(_23884_),
    .B(_04684_),
    .C(_04773_),
    .D(_00076_),
    .X(_06298_));
 sky130_fd_sc_hd__clkbuf_2 _34285_ (.A(_22363_),
    .X(_06299_));
 sky130_fd_sc_hd__nand2_1 _34286_ (.A(_23884_),
    .B(_03145_),
    .Y(_06300_));
 sky130_fd_sc_hd__or2_1 _34287_ (.A(_23884_),
    .B(_03145_),
    .X(_06301_));
 sky130_fd_sc_hd__a32o_1 _34288_ (.A1(_04683_),
    .A2(_04684_),
    .A3(_04773_),
    .B1(_06300_),
    .B2(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__and4b_2 _34289_ (.A_N(_06298_),
    .B(_06299_),
    .C(_06302_),
    .D(_03148_),
    .X(_06303_));
 sky130_fd_sc_hd__o31ai_1 _34290_ (.A1(_00108_),
    .A2(_03146_),
    .A3(_04687_),
    .B1(_06302_),
    .Y(_06305_));
 sky130_fd_sc_hd__and2_1 _34291_ (.A(_04759_),
    .B(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__o2bb2ai_2 _34292_ (.A1_N(_06291_),
    .A2_N(_06297_),
    .B1(_06303_),
    .B2(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__nor2_2 _34293_ (.A(_06303_),
    .B(_06306_),
    .Y(_06308_));
 sky130_fd_sc_hd__nand3_4 _34294_ (.A(_06291_),
    .B(_06297_),
    .C(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__nand2_1 _34295_ (.A(_04782_),
    .B(_04768_),
    .Y(_06310_));
 sky130_fd_sc_hd__a21oi_2 _34296_ (.A1(_06307_),
    .A2(_06309_),
    .B1(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__a21oi_2 _34297_ (.A1(_06291_),
    .A2(_06297_),
    .B1(_06308_),
    .Y(_06312_));
 sky130_fd_sc_hd__a31oi_4 _34298_ (.A1(_04748_),
    .A2(_04749_),
    .A3(_04756_),
    .B1(_04765_),
    .Y(_06313_));
 sky130_fd_sc_hd__o21ai_2 _34299_ (.A1(_04779_),
    .A2(_06313_),
    .B1(_06309_),
    .Y(_06314_));
 sky130_fd_sc_hd__nor2_1 _34300_ (.A(_06312_),
    .B(_06314_),
    .Y(_06316_));
 sky130_fd_sc_hd__o22ai_2 _34301_ (.A1(_06210_),
    .A2(_06211_),
    .B1(_06311_),
    .B2(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__or2_2 _34302_ (.A(_06210_),
    .B(_06211_),
    .X(_06318_));
 sky130_fd_sc_hd__inv_2 _34303_ (.A(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__a21o_2 _34304_ (.A1(_06307_),
    .A2(_06309_),
    .B1(_06310_),
    .X(_06320_));
 sky130_fd_sc_hd__o211ai_2 _34305_ (.A1(_06312_),
    .A2(_06314_),
    .B1(_06319_),
    .C1(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__nand3_4 _34306_ (.A(_06197_),
    .B(_06317_),
    .C(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__o21ai_4 _34307_ (.A1(_06311_),
    .A2(_06316_),
    .B1(_06319_),
    .Y(_06323_));
 sky130_fd_sc_hd__o211ai_4 _34308_ (.A1(_06314_),
    .A2(_06312_),
    .B1(_06318_),
    .C1(_06320_),
    .Y(_06324_));
 sky130_fd_sc_hd__a21boi_4 _34309_ (.A1(_04824_),
    .A2(_04823_),
    .B1_N(_04784_),
    .Y(_06325_));
 sky130_fd_sc_hd__nand3_4 _34310_ (.A(_06323_),
    .B(_06324_),
    .C(_06325_),
    .Y(_06327_));
 sky130_fd_sc_hd__o221a_1 _34311_ (.A1(_03286_),
    .A2(_01711_),
    .B1(_04863_),
    .B2(_04862_),
    .C1(_04851_),
    .X(_06328_));
 sky130_fd_sc_hd__or3b_1 _34312_ (.A(_06328_),
    .B(_04850_),
    .C_N(_04864_),
    .X(_06329_));
 sky130_fd_sc_hd__inv_2 _34313_ (.A(\delay_line[9][15] ),
    .Y(_06330_));
 sky130_fd_sc_hd__buf_1 _34314_ (.A(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__or2_1 _34315_ (.A(_25392_),
    .B(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__nand2_1 _34316_ (.A(_06331_),
    .B(_21821_),
    .Y(_06333_));
 sky130_fd_sc_hd__a22o_1 _34317_ (.A1(_21801_),
    .A2(_01692_),
    .B1(_06332_),
    .B2(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__clkbuf_2 _34318_ (.A(\delay_line[9][14] ),
    .X(_06335_));
 sky130_fd_sc_hd__and2b_1 _34319_ (.A_N(_22448_),
    .B(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__nand4_1 _34320_ (.A(_06332_),
    .B(_06333_),
    .C(_22458_),
    .D(_01694_),
    .Y(_06338_));
 sky130_fd_sc_hd__and3_1 _34321_ (.A(_06334_),
    .B(_06336_),
    .C(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__a21oi_1 _34322_ (.A1(_06338_),
    .A2(_06334_),
    .B1(_06336_),
    .Y(_06340_));
 sky130_fd_sc_hd__inv_2 _34323_ (.A(_23771_),
    .Y(_06341_));
 sky130_fd_sc_hd__nand2_1 _34324_ (.A(_06341_),
    .B(_23762_),
    .Y(_06342_));
 sky130_fd_sc_hd__nand2_1 _34325_ (.A(_01692_),
    .B(_04842_),
    .Y(_06343_));
 sky130_fd_sc_hd__nand3_1 _34326_ (.A(_06342_),
    .B(_06343_),
    .C(_03283_),
    .Y(_06344_));
 sky130_fd_sc_hd__a21o_1 _34327_ (.A1(_06342_),
    .A2(_06343_),
    .B1(_03281_),
    .X(_06345_));
 sky130_fd_sc_hd__and3b_1 _34328_ (.A_N(_04839_),
    .B(_06344_),
    .C(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__a21boi_1 _34329_ (.A1(_06344_),
    .A2(_06345_),
    .B1_N(_04840_),
    .Y(_06347_));
 sky130_fd_sc_hd__or4_2 _34330_ (.A(_06339_),
    .B(_06340_),
    .C(_06346_),
    .D(_06347_),
    .X(_06349_));
 sky130_fd_sc_hd__o22ai_1 _34331_ (.A1(_06339_),
    .A2(_06340_),
    .B1(_06346_),
    .B2(_06347_),
    .Y(_06350_));
 sky130_fd_sc_hd__nand2_2 _34332_ (.A(_06349_),
    .B(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__or2_1 _34333_ (.A(_04860_),
    .B(_04863_),
    .X(_06352_));
 sky130_fd_sc_hd__buf_1 _34334_ (.A(\delay_line[10][15] ),
    .X(_06353_));
 sky130_fd_sc_hd__nor2_1 _34335_ (.A(_23799_),
    .B(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand2_1 _34336_ (.A(_23799_),
    .B(_06353_),
    .Y(_06355_));
 sky130_fd_sc_hd__and4b_1 _34337_ (.A_N(_06354_),
    .B(_06355_),
    .C(_22465_),
    .D(_04856_),
    .X(_06356_));
 sky130_fd_sc_hd__and2_1 _34338_ (.A(_23798_),
    .B(\delay_line[10][15] ),
    .X(_06357_));
 sky130_fd_sc_hd__o2bb2a_1 _34339_ (.A1_N(_22465_),
    .A2_N(_04856_),
    .B1(_06354_),
    .B2(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__o2bb2a_1 _34340_ (.A1_N(_23799_),
    .A2_N(_04802_),
    .B1(_03126_),
    .B2(net400),
    .X(_06360_));
 sky130_fd_sc_hd__or3_1 _34341_ (.A(_06356_),
    .B(_06358_),
    .C(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__o21ai_1 _34342_ (.A1(_06356_),
    .A2(_06358_),
    .B1(_06360_),
    .Y(_06362_));
 sky130_fd_sc_hd__buf_1 _34343_ (.A(net411),
    .X(_06363_));
 sky130_fd_sc_hd__clkbuf_2 _34344_ (.A(_04856_),
    .X(_06364_));
 sky130_fd_sc_hd__nand2_1 _34345_ (.A(_25372_),
    .B(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__and4b_1 _34346_ (.A_N(_04857_),
    .B(_06363_),
    .C(_21805_),
    .D(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__a21o_1 _34347_ (.A1(_06361_),
    .A2(_06362_),
    .B1(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nand3_1 _34348_ (.A(_06361_),
    .B(_06362_),
    .C(_06366_),
    .Y(_06368_));
 sky130_fd_sc_hd__a21oi_1 _34349_ (.A1(_06368_),
    .A2(_06367_),
    .B1(_06352_),
    .Y(_06369_));
 sky130_fd_sc_hd__a21o_1 _34350_ (.A1(_06352_),
    .A2(_06367_),
    .B1(_06369_),
    .X(_06371_));
 sky130_fd_sc_hd__xor2_4 _34351_ (.A(_06351_),
    .B(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__o21a_1 _34352_ (.A1(_04809_),
    .A2(_04813_),
    .B1(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__a31o_1 _34353_ (.A1(_04806_),
    .A2(_04807_),
    .A3(_04808_),
    .B1(_04813_),
    .X(_06374_));
 sky130_fd_sc_hd__nor2_1 _34354_ (.A(_06374_),
    .B(_06372_),
    .Y(_06375_));
 sky130_fd_sc_hd__or2_1 _34355_ (.A(_06373_),
    .B(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__a21oi_4 _34356_ (.A1(_04864_),
    .A2(_06329_),
    .B1(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__o211a_1 _34357_ (.A1(_06328_),
    .A2(_04850_),
    .B1(_04864_),
    .C1(_06376_),
    .X(_06378_));
 sky130_fd_sc_hd__nor2_1 _34358_ (.A(_06377_),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__clkbuf_2 _34359_ (.A(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__a21oi_4 _34360_ (.A1(_06322_),
    .A2(_06327_),
    .B1(_06380_),
    .Y(_06382_));
 sky130_fd_sc_hd__o211ai_4 _34361_ (.A1(_04779_),
    .A2(_06313_),
    .B1(_06307_),
    .C1(_06309_),
    .Y(_06383_));
 sky130_fd_sc_hd__a21oi_2 _34362_ (.A1(_06320_),
    .A2(_06383_),
    .B1(_06318_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand2_1 _34363_ (.A(_06324_),
    .B(_06325_),
    .Y(_06385_));
 sky130_fd_sc_hd__o211a_1 _34364_ (.A1(_06384_),
    .A2(_06385_),
    .B1(_06380_),
    .C1(_06322_),
    .X(_06386_));
 sky130_fd_sc_hd__o2bb2ai_2 _34365_ (.A1_N(_04873_),
    .A2_N(_04820_),
    .B1(_04881_),
    .B2(_04878_),
    .Y(_06387_));
 sky130_fd_sc_hd__o21bai_4 _34366_ (.A1(_06382_),
    .A2(_06386_),
    .B1_N(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__nand2_2 _34367_ (.A(_06327_),
    .B(_06380_),
    .Y(_06389_));
 sky130_fd_sc_hd__a21oi_2 _34368_ (.A1(_06323_),
    .A2(_06324_),
    .B1(_06325_),
    .Y(_06390_));
 sky130_fd_sc_hd__buf_4 _34369_ (.A(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__buf_2 _34370_ (.A(_06387_),
    .X(_06393_));
 sky130_fd_sc_hd__o2bb2ai_4 _34371_ (.A1_N(_06322_),
    .A2_N(_06327_),
    .B1(_06377_),
    .B2(_06378_),
    .Y(_06394_));
 sky130_fd_sc_hd__o211ai_4 _34372_ (.A1(_06389_),
    .A2(_06391_),
    .B1(_06393_),
    .C1(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__or2_1 _34373_ (.A(_04631_),
    .B(_04674_),
    .X(_06396_));
 sky130_fd_sc_hd__nand3b_1 _34374_ (.A_N(_03365_),
    .B(_03371_),
    .C(_04650_),
    .Y(_06397_));
 sky130_fd_sc_hd__o21ai_2 _34375_ (.A1(_03367_),
    .A2(net423),
    .B1(\delay_line[8][12] ),
    .Y(_06398_));
 sky130_fd_sc_hd__and2_1 _34376_ (.A(\delay_line[8][13] ),
    .B(\delay_line[8][14] ),
    .X(_06399_));
 sky130_fd_sc_hd__buf_2 _34377_ (.A(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__and2_1 _34378_ (.A(_01770_),
    .B(_03367_),
    .X(_06401_));
 sky130_fd_sc_hd__a21boi_1 _34379_ (.A1(_04635_),
    .A2(_04636_),
    .B1_N(\delay_line[8][11] ),
    .Y(_06402_));
 sky130_fd_sc_hd__nor2_1 _34380_ (.A(_03367_),
    .B(_04649_),
    .Y(_06404_));
 sky130_fd_sc_hd__o21bai_2 _34381_ (.A1(_06399_),
    .A2(_06404_),
    .B1_N(_01770_),
    .Y(_06405_));
 sky130_fd_sc_hd__o221ai_4 _34382_ (.A1(_06398_),
    .A2(_06400_),
    .B1(_06401_),
    .B2(_06402_),
    .C1(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__o21ai_1 _34383_ (.A1(_06400_),
    .A2(_06398_),
    .B1(_06405_),
    .Y(_06407_));
 sky130_fd_sc_hd__a21oi_1 _34384_ (.A1(_04637_),
    .A2(_25308_),
    .B1(_06401_),
    .Y(_06408_));
 sky130_fd_sc_hd__nand2_1 _34385_ (.A(_06407_),
    .B(_06408_),
    .Y(_06409_));
 sky130_fd_sc_hd__a21o_1 _34386_ (.A1(_06406_),
    .A2(_06409_),
    .B1(_01740_),
    .X(_06410_));
 sky130_fd_sc_hd__nand3_1 _34387_ (.A(_06406_),
    .B(_06409_),
    .C(_25313_),
    .Y(_06411_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34388_ (.A(_04649_),
    .X(_06412_));
 sky130_fd_sc_hd__nand2_1 _34389_ (.A(_22543_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__nand3b_1 _34390_ (.A_N(_17915_),
    .B(_03369_),
    .C(_04650_),
    .Y(_06415_));
 sky130_fd_sc_hd__clkbuf_2 _34391_ (.A(\delay_line[8][15] ),
    .X(_06416_));
 sky130_fd_sc_hd__and2b_1 _34392_ (.A_N(_20125_),
    .B(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__and2b_1 _34393_ (.A_N(_06416_),
    .B(_20125_),
    .X(_06418_));
 sky130_fd_sc_hd__nor2_1 _34394_ (.A(_06417_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__and3_1 _34395_ (.A(_06413_),
    .B(_06415_),
    .C(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__a21oi_1 _34396_ (.A1(_06413_),
    .A2(_06415_),
    .B1(_06419_),
    .Y(_06421_));
 sky130_fd_sc_hd__a211oi_1 _34397_ (.A1(_06410_),
    .A2(_06411_),
    .B1(_06420_),
    .C1(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__o211a_1 _34398_ (.A1(_06420_),
    .A2(_06421_),
    .B1(_06410_),
    .C1(_06411_),
    .X(_06423_));
 sky130_fd_sc_hd__a211oi_1 _34399_ (.A1(_04654_),
    .A2(_06397_),
    .B1(_06422_),
    .C1(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__o211ai_1 _34400_ (.A1(_06422_),
    .A2(_06423_),
    .B1(_04654_),
    .C1(_06397_),
    .Y(_06426_));
 sky130_fd_sc_hd__and2b_1 _34401_ (.A_N(_06424_),
    .B(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__buf_1 _34402_ (.A(\delay_line[7][15] ),
    .X(_06428_));
 sky130_fd_sc_hd__and2_1 _34403_ (.A(_23953_),
    .B(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__buf_1 _34404_ (.A(_06428_),
    .X(_06430_));
 sky130_fd_sc_hd__nor2_1 _34405_ (.A(_23953_),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__clkbuf_2 _34406_ (.A(_04659_),
    .X(_06432_));
 sky130_fd_sc_hd__and2b_1 _34407_ (.A_N(_01767_),
    .B(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__o21a_1 _34408_ (.A1(_06429_),
    .A2(_06431_),
    .B1(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__nor3_1 _34409_ (.A(_06433_),
    .B(_06429_),
    .C(_06431_),
    .Y(_06435_));
 sky130_fd_sc_hd__a211oi_2 _34410_ (.A1(_04640_),
    .A2(_04644_),
    .B1(_06434_),
    .C1(net251),
    .Y(_06437_));
 sky130_fd_sc_hd__inv_2 _34411_ (.A(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__o211ai_2 _34412_ (.A1(_06434_),
    .A2(net251),
    .B1(_04640_),
    .C1(_04644_),
    .Y(_06439_));
 sky130_fd_sc_hd__a32o_1 _34413_ (.A1(_03336_),
    .A2(_04660_),
    .A3(_04661_),
    .B1(_06438_),
    .B2(_06439_),
    .X(_06440_));
 sky130_fd_sc_hd__nand3_1 _34414_ (.A(_06438_),
    .B(_06439_),
    .C(_04662_),
    .Y(_06441_));
 sky130_fd_sc_hd__nand3_1 _34415_ (.A(_06427_),
    .B(_06440_),
    .C(_06441_),
    .Y(_06442_));
 sky130_fd_sc_hd__a21o_1 _34416_ (.A1(_06441_),
    .A2(_06440_),
    .B1(_06427_),
    .X(_06443_));
 sky130_fd_sc_hd__nand4_1 _34417_ (.A(_04840_),
    .B(_04841_),
    .C(_04844_),
    .D(_04845_),
    .Y(_06444_));
 sky130_fd_sc_hd__clkbuf_2 _34418_ (.A(_04614_),
    .X(_06445_));
 sky130_fd_sc_hd__o21ba_1 _34419_ (.A1(_06445_),
    .A2(_03314_),
    .B1_N(_04617_),
    .X(_06446_));
 sky130_fd_sc_hd__a21boi_1 _34420_ (.A1(_04831_),
    .A2(_04833_),
    .B1_N(_04834_),
    .Y(_06448_));
 sky130_fd_sc_hd__a21oi_1 _34421_ (.A1(_01682_),
    .A2(net416),
    .B1(_04828_),
    .Y(_06449_));
 sky130_fd_sc_hd__and3_1 _34422_ (.A(_01681_),
    .B(net416),
    .C(\delay_line[9][14] ),
    .X(_06450_));
 sky130_fd_sc_hd__o21a_1 _34423_ (.A1(_06449_),
    .A2(_06450_),
    .B1(_23755_),
    .X(_06451_));
 sky130_fd_sc_hd__inv_2 _34424_ (.A(_06451_),
    .Y(_06452_));
 sky130_fd_sc_hd__or3_2 _34425_ (.A(_23755_),
    .B(_06449_),
    .C(_06450_),
    .X(_06453_));
 sky130_fd_sc_hd__and3b_1 _34426_ (.A_N(_06448_),
    .B(_06452_),
    .C(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__a21boi_1 _34427_ (.A1(_06452_),
    .A2(_06453_),
    .B1_N(_06448_),
    .Y(_06455_));
 sky130_fd_sc_hd__nor2_1 _34428_ (.A(_06454_),
    .B(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__xor2_1 _34429_ (.A(_06446_),
    .B(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__o311a_1 _34430_ (.A1(_04835_),
    .A2(_04836_),
    .A3(_04847_),
    .B1(_06444_),
    .C1(_06457_),
    .X(_06459_));
 sky130_fd_sc_hd__a21oi_1 _34431_ (.A1(_06444_),
    .A2(_04848_),
    .B1(_06457_),
    .Y(_06460_));
 sky130_fd_sc_hd__a21boi_1 _34432_ (.A1(_04621_),
    .A2(_04620_),
    .B1_N(_04619_),
    .Y(_06461_));
 sky130_fd_sc_hd__o21a_1 _34433_ (.A1(_06459_),
    .A2(_06460_),
    .B1(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__nor3_1 _34434_ (.A(_06461_),
    .B(_06459_),
    .C(_06460_),
    .Y(_06463_));
 sky130_fd_sc_hd__o211ai_1 _34435_ (.A1(_06462_),
    .A2(_06463_),
    .B1(_04627_),
    .C1(_04628_),
    .Y(_06464_));
 sky130_fd_sc_hd__a211o_1 _34436_ (.A1(_04627_),
    .A2(_04628_),
    .B1(_06462_),
    .C1(_06463_),
    .X(_06465_));
 sky130_fd_sc_hd__and4_1 _34437_ (.A(_06442_),
    .B(_06443_),
    .C(_06464_),
    .D(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34438_ (.A(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__a22oi_1 _34439_ (.A1(_06442_),
    .A2(_06443_),
    .B1(_06464_),
    .B2(_06465_),
    .Y(_06468_));
 sky130_fd_sc_hd__a21oi_2 _34440_ (.A1(_04871_),
    .A2(_04872_),
    .B1(_04869_),
    .Y(_06470_));
 sky130_fd_sc_hd__o21ai_1 _34441_ (.A1(_06467_),
    .A2(_06468_),
    .B1(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__or3_1 _34442_ (.A(_06470_),
    .B(_06466_),
    .C(_06468_),
    .X(_06472_));
 sky130_fd_sc_hd__and3_1 _34443_ (.A(_06396_),
    .B(_06471_),
    .C(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__a21oi_1 _34444_ (.A1(_06471_),
    .A2(_06472_),
    .B1(_06396_),
    .Y(_06474_));
 sky130_fd_sc_hd__or2_4 _34445_ (.A(_06473_),
    .B(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__inv_2 _34446_ (.A(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__a21oi_4 _34447_ (.A1(_06388_),
    .A2(_06395_),
    .B1(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__nor2_1 _34448_ (.A(_04681_),
    .B(_04682_),
    .Y(_06478_));
 sky130_fd_sc_hd__o22ai_4 _34449_ (.A1(_04883_),
    .A2(_04875_),
    .B1(_06478_),
    .B2(_04896_),
    .Y(_06479_));
 sky130_fd_sc_hd__nand3_2 _34450_ (.A(_06388_),
    .B(_06395_),
    .C(_06476_),
    .Y(_06481_));
 sky130_fd_sc_hd__nand2_4 _34451_ (.A(_06479_),
    .B(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__o211ai_2 _34452_ (.A1(_06384_),
    .A2(_06385_),
    .B1(_06380_),
    .C1(_06322_),
    .Y(_06483_));
 sky130_fd_sc_hd__a21oi_4 _34453_ (.A1(_06394_),
    .A2(_06483_),
    .B1(_06393_),
    .Y(_06484_));
 sky130_fd_sc_hd__o211a_1 _34454_ (.A1(_06389_),
    .A2(_06390_),
    .B1(_06393_),
    .C1(_06394_),
    .X(_06485_));
 sky130_fd_sc_hd__o21bai_4 _34455_ (.A1(_06484_),
    .A2(_06485_),
    .B1_N(_06475_),
    .Y(_06486_));
 sky130_fd_sc_hd__o22a_2 _34456_ (.A1(_04883_),
    .A2(_04874_),
    .B1(_06478_),
    .B2(_04896_),
    .X(_06487_));
 sky130_fd_sc_hd__o21ai_4 _34457_ (.A1(_06390_),
    .A2(_06389_),
    .B1(_06393_),
    .Y(_06488_));
 sky130_fd_sc_hd__o211ai_4 _34458_ (.A1(_06488_),
    .A2(_06382_),
    .B1(_06475_),
    .C1(_06388_),
    .Y(_06489_));
 sky130_fd_sc_hd__nand3_1 _34459_ (.A(_06486_),
    .B(_06487_),
    .C(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__o21ai_1 _34460_ (.A1(_06477_),
    .A2(_06482_),
    .B1(_06490_),
    .Y(_06492_));
 sky130_fd_sc_hd__nand2_1 _34461_ (.A(_06196_),
    .B(_06492_),
    .Y(_06493_));
 sky130_fd_sc_hd__buf_6 _34462_ (.A(_06490_),
    .X(_06494_));
 sky130_fd_sc_hd__o211ai_4 _34463_ (.A1(_06477_),
    .A2(_06482_),
    .B1(_06195_),
    .C1(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__a31o_1 _34464_ (.A1(_04900_),
    .A2(_04901_),
    .A3(_04902_),
    .B1(_05013_),
    .X(_06496_));
 sky130_fd_sc_hd__nand2_2 _34465_ (.A(_04899_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__a21oi_2 _34466_ (.A1(_06493_),
    .A2(_06495_),
    .B1(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand2_2 _34467_ (.A(_06497_),
    .B(_06495_),
    .Y(_06499_));
 sky130_fd_sc_hd__a21oi_1 _34468_ (.A1(_06196_),
    .A2(_06492_),
    .B1(_06499_),
    .Y(_06500_));
 sky130_fd_sc_hd__nand2_1 _34469_ (.A(_05003_),
    .B(_04905_),
    .Y(_06501_));
 sky130_fd_sc_hd__or2_1 _34470_ (.A(_04904_),
    .B(_05004_),
    .X(_06503_));
 sky130_fd_sc_hd__a21boi_1 _34471_ (.A1(_05049_),
    .A2(_05046_),
    .B1_N(_05048_),
    .Y(_06504_));
 sky130_fd_sc_hd__a21oi_1 _34472_ (.A1(_03099_),
    .A2(_03101_),
    .B1(_05043_),
    .Y(_06505_));
 sky130_fd_sc_hd__o21ba_1 _34473_ (.A1(_05040_),
    .A2(_05042_),
    .B1_N(_06505_),
    .X(_06506_));
 sky130_fd_sc_hd__o21ai_1 _34474_ (.A1(_03490_),
    .A2(_03493_),
    .B1(_04923_),
    .Y(_06507_));
 sky130_fd_sc_hd__a21oi_1 _34475_ (.A1(_03090_),
    .A2(_03091_),
    .B1(_03086_),
    .Y(_06508_));
 sky130_fd_sc_hd__xnor2_1 _34476_ (.A(_01493_),
    .B(_05026_),
    .Y(_06509_));
 sky130_fd_sc_hd__inv_2 _34477_ (.A(net445),
    .Y(_06510_));
 sky130_fd_sc_hd__nand2_1 _34478_ (.A(_05024_),
    .B(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__nand2_1 _34479_ (.A(net446),
    .B(net445),
    .Y(_06512_));
 sky130_fd_sc_hd__a21o_1 _34480_ (.A1(_06511_),
    .A2(_06512_),
    .B1(_03488_),
    .X(_06514_));
 sky130_fd_sc_hd__nand3_1 _34481_ (.A(_06511_),
    .B(_06512_),
    .C(_03488_),
    .Y(_06515_));
 sky130_fd_sc_hd__and3_1 _34482_ (.A(_05029_),
    .B(_06514_),
    .C(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__a21oi_1 _34483_ (.A1(_06514_),
    .A2(_06515_),
    .B1(_05029_),
    .Y(_06517_));
 sky130_fd_sc_hd__nor3_1 _34484_ (.A(_06509_),
    .B(_06516_),
    .C(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__o21a_1 _34485_ (.A1(_06516_),
    .A2(_06517_),
    .B1(_06509_),
    .X(_06519_));
 sky130_fd_sc_hd__nor4_1 _34486_ (.A(_05031_),
    .B(_05036_),
    .C(_06518_),
    .D(_06519_),
    .Y(_06520_));
 sky130_fd_sc_hd__o22a_1 _34487_ (.A1(_05031_),
    .A2(_05036_),
    .B1(_06518_),
    .B2(_06519_),
    .X(_06521_));
 sky130_fd_sc_hd__nor4_1 _34488_ (.A(_00319_),
    .B(_06508_),
    .C(_06520_),
    .D(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__o22a_1 _34489_ (.A1(_00319_),
    .A2(_06508_),
    .B1(_06520_),
    .B2(_06521_),
    .X(_06523_));
 sky130_fd_sc_hd__or2_1 _34490_ (.A(_06522_),
    .B(_06523_),
    .X(_06525_));
 sky130_fd_sc_hd__a21o_1 _34491_ (.A1(_04922_),
    .A2(_06507_),
    .B1(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__o211ai_1 _34492_ (.A1(_04906_),
    .A2(_04921_),
    .B1(_04922_),
    .C1(_06525_),
    .Y(_06527_));
 sky130_fd_sc_hd__nand2_1 _34493_ (.A(_06526_),
    .B(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__a21o_1 _34494_ (.A1(_05020_),
    .A2(_05039_),
    .B1(_05037_),
    .X(_06529_));
 sky130_fd_sc_hd__nand2_1 _34495_ (.A(_06528_),
    .B(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__a211o_1 _34496_ (.A1(_05020_),
    .A2(_05039_),
    .B1(_05037_),
    .C1(_06528_),
    .X(_06531_));
 sky130_fd_sc_hd__nand3b_1 _34497_ (.A_N(_04925_),
    .B(_04963_),
    .C(_04965_),
    .Y(_06532_));
 sky130_fd_sc_hd__o2111ai_1 _34498_ (.A1(_04924_),
    .A2(_04967_),
    .B1(_06530_),
    .C1(_06531_),
    .D1(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__o21ai_1 _34499_ (.A1(_04924_),
    .A2(_04967_),
    .B1(_06532_),
    .Y(_06534_));
 sky130_fd_sc_hd__a21bo_1 _34500_ (.A1(_06530_),
    .A2(_06531_),
    .B1_N(_06534_),
    .X(_06536_));
 sky130_fd_sc_hd__nand2_1 _34501_ (.A(_06533_),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__nor2_1 _34502_ (.A(_06506_),
    .B(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__and2_1 _34503_ (.A(_06537_),
    .B(_06506_),
    .X(_06539_));
 sky130_fd_sc_hd__or3_1 _34504_ (.A(_06504_),
    .B(_06538_),
    .C(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__o21ai_1 _34505_ (.A1(_06538_),
    .A2(_06539_),
    .B1(_06504_),
    .Y(_06541_));
 sky130_fd_sc_hd__nand2_1 _34506_ (.A(_06540_),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__a21oi_2 _34507_ (.A1(_06501_),
    .A2(_06503_),
    .B1(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__o211ai_2 _34508_ (.A1(_05004_),
    .A2(_04904_),
    .B1(_06501_),
    .C1(_06542_),
    .Y(_06544_));
 sky130_fd_sc_hd__or2b_2 _34509_ (.A(_06543_),
    .B_N(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__xnor2_2 _34510_ (.A(_05055_),
    .B(_06545_),
    .Y(_06547_));
 sky130_fd_sc_hd__o21ai_2 _34511_ (.A1(_06498_),
    .A2(_06500_),
    .B1(_06547_),
    .Y(_06548_));
 sky130_fd_sc_hd__or2_1 _34512_ (.A(_06081_),
    .B(_06193_),
    .X(_06549_));
 sky130_fd_sc_hd__nand2_2 _34513_ (.A(_06193_),
    .B(_06081_),
    .Y(_06550_));
 sky130_fd_sc_hd__o21ai_1 _34514_ (.A1(_06484_),
    .A2(_06485_),
    .B1(_06475_),
    .Y(_06551_));
 sky130_fd_sc_hd__nand3_2 _34515_ (.A(_06479_),
    .B(_06551_),
    .C(_06481_),
    .Y(_06552_));
 sky130_fd_sc_hd__a22oi_4 _34516_ (.A1(_06549_),
    .A2(_06550_),
    .B1(_06552_),
    .B2(_06494_),
    .Y(_06553_));
 sky130_fd_sc_hd__xor2_4 _34517_ (.A(_05055_),
    .B(_06545_),
    .X(_06554_));
 sky130_fd_sc_hd__o211a_1 _34518_ (.A1(_06477_),
    .A2(_06482_),
    .B1(_06195_),
    .C1(_06494_),
    .X(_06555_));
 sky130_fd_sc_hd__o21bai_4 _34519_ (.A1(_06553_),
    .A2(_06555_),
    .B1_N(_06497_),
    .Y(_06556_));
 sky130_fd_sc_hd__o211ai_4 _34520_ (.A1(_06499_),
    .A2(_06553_),
    .B1(_06554_),
    .C1(_06556_),
    .Y(_06558_));
 sky130_fd_sc_hd__o211ai_2 _34521_ (.A1(_05011_),
    .A2(_06080_),
    .B1(_06548_),
    .C1(_06558_),
    .Y(_06559_));
 sky130_fd_sc_hd__nand3_1 _34522_ (.A(_06497_),
    .B(_06493_),
    .C(_06495_),
    .Y(_06560_));
 sky130_fd_sc_hd__a21oi_2 _34523_ (.A1(_06556_),
    .A2(_06560_),
    .B1(_06554_),
    .Y(_06561_));
 sky130_fd_sc_hd__o211a_1 _34524_ (.A1(_06499_),
    .A2(_06553_),
    .B1(_06554_),
    .C1(_06556_),
    .X(_06562_));
 sky130_fd_sc_hd__a2bb2o_1 _34525_ (.A1_N(_05006_),
    .A2_N(_05010_),
    .B1(_05065_),
    .B2(_05070_),
    .X(_06563_));
 sky130_fd_sc_hd__o21bai_4 _34526_ (.A1(_06561_),
    .A2(_06562_),
    .B1_N(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__or2_2 _34527_ (.A(_05060_),
    .B(_05068_),
    .X(_06565_));
 sky130_fd_sc_hd__a21oi_2 _34528_ (.A1(_06559_),
    .A2(_06564_),
    .B1(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__and3_1 _34529_ (.A(_05075_),
    .B(_05076_),
    .C(_05077_),
    .X(_06567_));
 sky130_fd_sc_hd__a21o_1 _34530_ (.A1(_05080_),
    .A2(_05073_),
    .B1(_06567_),
    .X(_06569_));
 sky130_fd_sc_hd__buf_2 _34531_ (.A(_06561_),
    .X(_06570_));
 sky130_fd_sc_hd__o21ai_4 _34532_ (.A1(_05011_),
    .A2(_06080_),
    .B1(_06558_),
    .Y(_06571_));
 sky130_fd_sc_hd__o221ai_4 _34533_ (.A1(_05060_),
    .A2(_05068_),
    .B1(_06570_),
    .B2(_06571_),
    .C1(_06564_),
    .Y(_06572_));
 sky130_fd_sc_hd__nand2_1 _34534_ (.A(_06569_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__nor2_1 _34535_ (.A(_06570_),
    .B(_06571_),
    .Y(_06574_));
 sky130_fd_sc_hd__a21oi_4 _34536_ (.A1(_06548_),
    .A2(_06558_),
    .B1(_06563_),
    .Y(_06575_));
 sky130_fd_sc_hd__o22ai_4 _34537_ (.A1(_05060_),
    .A2(_05068_),
    .B1(_06574_),
    .B2(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__a21boi_4 _34538_ (.A1(_05080_),
    .A2(_05073_),
    .B1_N(_05078_),
    .Y(_06577_));
 sky130_fd_sc_hd__inv_2 _34539_ (.A(_06565_),
    .Y(_06578_));
 sky130_fd_sc_hd__o211ai_4 _34540_ (.A1(_06570_),
    .A2(_06571_),
    .B1(_06578_),
    .C1(_06564_),
    .Y(_06580_));
 sky130_fd_sc_hd__nand3_4 _34541_ (.A(_06576_),
    .B(_06577_),
    .C(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__o21ai_4 _34542_ (.A1(_06566_),
    .A2(_06573_),
    .B1(_06581_),
    .Y(_06582_));
 sky130_fd_sc_hd__a21oi_4 _34543_ (.A1(_05093_),
    .A2(_05095_),
    .B1(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__nand2_1 _34544_ (.A(_05092_),
    .B(_05083_),
    .Y(_06584_));
 sky130_fd_sc_hd__o211ai_4 _34545_ (.A1(_06584_),
    .A2(_05088_),
    .B1(_06582_),
    .C1(_05094_),
    .Y(_06585_));
 sky130_fd_sc_hd__clkbuf_4 _34546_ (.A(\delay_line[23][15] ),
    .X(_06586_));
 sky130_fd_sc_hd__nand2_2 _34547_ (.A(_06585_),
    .B(_06586_),
    .Y(_06587_));
 sky130_fd_sc_hd__clkbuf_2 _34548_ (.A(\delay_line[23][14] ),
    .X(_06588_));
 sky130_fd_sc_hd__a21oi_1 _34549_ (.A1(_05092_),
    .A2(_05083_),
    .B1(_05087_),
    .Y(_06589_));
 sky130_fd_sc_hd__a31o_1 _34550_ (.A1(_01975_),
    .A2(_01973_),
    .A3(_01962_),
    .B1(_03533_),
    .X(_06591_));
 sky130_fd_sc_hd__a2bb2o_1 _34551_ (.A1_N(_03539_),
    .A2_N(_03540_),
    .B1(_03534_),
    .B2(_03531_),
    .X(_06592_));
 sky130_fd_sc_hd__o2bb2ai_4 _34552_ (.A1_N(_03558_),
    .A2_N(_01999_),
    .B1(_06591_),
    .B2(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__o21ai_1 _34553_ (.A1(_06589_),
    .A2(_06593_),
    .B1(_05093_),
    .Y(_06594_));
 sky130_fd_sc_hd__a31oi_2 _34554_ (.A1(_06559_),
    .A2(_06564_),
    .A3(_06565_),
    .B1(_06577_),
    .Y(_06595_));
 sky130_fd_sc_hd__o21ai_2 _34555_ (.A1(_06574_),
    .A2(_06575_),
    .B1(_06578_),
    .Y(_06596_));
 sky130_fd_sc_hd__a32oi_4 _34556_ (.A1(_06576_),
    .A2(_06577_),
    .A3(_06580_),
    .B1(_06595_),
    .B2(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__nand2_1 _34557_ (.A(_06594_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__a21o_1 _34558_ (.A1(_06598_),
    .A2(_06585_),
    .B1(_06586_),
    .X(_06599_));
 sky130_fd_sc_hd__o211ai_4 _34559_ (.A1(_06583_),
    .A2(_06587_),
    .B1(_06588_),
    .C1(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__nor2_1 _34560_ (.A(_06583_),
    .B(_06587_),
    .Y(_06602_));
 sky130_fd_sc_hd__a21oi_2 _34561_ (.A1(_06598_),
    .A2(_06585_),
    .B1(_06586_),
    .Y(_06603_));
 sky130_fd_sc_hd__o21bai_2 _34562_ (.A1(_06602_),
    .A2(_06603_),
    .B1_N(_06588_),
    .Y(_06604_));
 sky130_fd_sc_hd__o21bai_4 _34563_ (.A1(_05391_),
    .A2(_05357_),
    .B1_N(_05393_),
    .Y(_06605_));
 sky130_fd_sc_hd__a21oi_2 _34564_ (.A1(_06600_),
    .A2(_06604_),
    .B1(_06605_),
    .Y(_06606_));
 sky130_fd_sc_hd__clkbuf_2 _34565_ (.A(_06588_),
    .X(_06607_));
 sky130_fd_sc_hd__nand2_1 _34566_ (.A(_06599_),
    .B(_06607_),
    .Y(_06608_));
 sky130_fd_sc_hd__o211a_1 _34567_ (.A1(_06602_),
    .A2(_06608_),
    .B1(_06604_),
    .C1(_06605_),
    .X(_06609_));
 sky130_fd_sc_hd__o21ai_2 _34568_ (.A1(_05098_),
    .A2(_05097_),
    .B1(_05099_),
    .Y(_06610_));
 sky130_fd_sc_hd__o21ai_4 _34569_ (.A1(_06606_),
    .A2(_06609_),
    .B1(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__a21oi_2 _34570_ (.A1(_05340_),
    .A2(_05396_),
    .B1(_05339_),
    .Y(_06613_));
 sky130_fd_sc_hd__a21o_1 _34571_ (.A1(_06600_),
    .A2(_06604_),
    .B1(_06605_),
    .X(_06614_));
 sky130_fd_sc_hd__nand3_2 _34572_ (.A(_06605_),
    .B(_06600_),
    .C(_06604_),
    .Y(_06615_));
 sky130_fd_sc_hd__o21a_1 _34573_ (.A1(_05098_),
    .A2(_05097_),
    .B1(_05099_),
    .X(_06616_));
 sky130_fd_sc_hd__nand3_2 _34574_ (.A(_06614_),
    .B(_06615_),
    .C(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__nand3_2 _34575_ (.A(_06611_),
    .B(_06613_),
    .C(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__o21ai_2 _34576_ (.A1(_06078_),
    .A2(_05108_),
    .B1(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__a2bb2oi_2 _34577_ (.A1_N(_05339_),
    .A2_N(_05397_),
    .B1(_06617_),
    .B2(_06611_),
    .Y(_06620_));
 sky130_fd_sc_hd__o21ai_2 _34578_ (.A1(_05126_),
    .A2(_05125_),
    .B1(_05117_),
    .Y(_06621_));
 sky130_fd_sc_hd__nand3_1 _34579_ (.A(_06614_),
    .B(_06615_),
    .C(_06610_),
    .Y(_06622_));
 sky130_fd_sc_hd__o21bai_1 _34580_ (.A1(_06606_),
    .A2(_06609_),
    .B1_N(_06610_),
    .Y(_06624_));
 sky130_fd_sc_hd__o211ai_4 _34581_ (.A1(_05339_),
    .A2(_05397_),
    .B1(_06622_),
    .C1(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__nor2_1 _34582_ (.A(_06078_),
    .B(_05106_),
    .Y(_06626_));
 sky130_fd_sc_hd__inv_2 _34583_ (.A(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__a21o_1 _34584_ (.A1(_06618_),
    .A2(_06625_),
    .B1(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__o211ai_2 _34585_ (.A1(_06619_),
    .A2(_06620_),
    .B1(_06621_),
    .C1(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__a21oi_1 _34586_ (.A1(_06618_),
    .A2(_06625_),
    .B1(_06627_),
    .Y(_06630_));
 sky130_fd_sc_hd__o211a_1 _34587_ (.A1(_06078_),
    .A2(_05108_),
    .B1(_06618_),
    .C1(_06625_),
    .X(_06631_));
 sky130_fd_sc_hd__o21bai_2 _34588_ (.A1(_06630_),
    .A2(_06631_),
    .B1_N(_06621_),
    .Y(_06632_));
 sky130_fd_sc_hd__buf_1 _34589_ (.A(_22110_),
    .X(_06633_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34590_ (.A(_19217_),
    .X(_06635_));
 sky130_fd_sc_hd__nand2_2 _34591_ (.A(_22129_),
    .B(_22110_),
    .Y(_06636_));
 sky130_fd_sc_hd__or2_1 _34592_ (.A(_22129_),
    .B(_22110_),
    .X(_06637_));
 sky130_fd_sc_hd__a22o_1 _34593_ (.A1(_19849_),
    .A2(_22130_),
    .B1(_06636_),
    .B2(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__o21a_1 _34594_ (.A1(_06633_),
    .A2(_06635_),
    .B1(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__nor2_1 _34595_ (.A(_02019_),
    .B(_03066_),
    .Y(_06640_));
 sky130_fd_sc_hd__and2_1 _34596_ (.A(_02019_),
    .B(_03066_),
    .X(_06641_));
 sky130_fd_sc_hd__or3_1 _34597_ (.A(_06640_),
    .B(_05137_),
    .C(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34598_ (.A(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__buf_1 _34599_ (.A(_24241_),
    .X(_06644_));
 sky130_fd_sc_hd__a2bb2o_1 _34600_ (.A1_N(_06641_),
    .A2_N(_06640_),
    .B1(_06644_),
    .B2(_03565_),
    .X(_06646_));
 sky130_fd_sc_hd__and3_1 _34601_ (.A(_06639_),
    .B(_06643_),
    .C(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__a21oi_2 _34602_ (.A1(_06643_),
    .A2(_06646_),
    .B1(_06639_),
    .Y(_06648_));
 sky130_fd_sc_hd__o2bb2ai_1 _34603_ (.A1_N(_06629_),
    .A2_N(_06632_),
    .B1(_06647_),
    .B2(_06648_),
    .Y(_06649_));
 sky130_fd_sc_hd__inv_2 _34604_ (.A(_06639_),
    .Y(_06650_));
 sky130_fd_sc_hd__and3_1 _34605_ (.A(_06650_),
    .B(_06643_),
    .C(_06646_),
    .X(_06651_));
 sky130_fd_sc_hd__nand2_1 _34606_ (.A(_06642_),
    .B(_06646_),
    .Y(_06652_));
 sky130_fd_sc_hd__o211a_1 _34607_ (.A1(_06633_),
    .A2(_06635_),
    .B1(_06638_),
    .C1(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__buf_4 _34608_ (.A(_06629_),
    .X(_06654_));
 sky130_fd_sc_hd__clkbuf_2 _34609_ (.A(_06632_),
    .X(_06655_));
 sky130_fd_sc_hd__o211ai_1 _34610_ (.A1(_06651_),
    .A2(_06653_),
    .B1(_06654_),
    .C1(_06655_),
    .Y(_06657_));
 sky130_fd_sc_hd__nand3b_1 _34611_ (.A_N(_06077_),
    .B(_06649_),
    .C(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__clkbuf_2 _34612_ (.A(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__o2bb2ai_2 _34613_ (.A1_N(_06654_),
    .A2_N(_06655_),
    .B1(_06651_),
    .B2(_06653_),
    .Y(_06660_));
 sky130_fd_sc_hd__o211ai_4 _34614_ (.A1(_06647_),
    .A2(_06648_),
    .B1(_06654_),
    .C1(_06655_),
    .Y(_06661_));
 sky130_fd_sc_hd__a21o_1 _34615_ (.A1(_05146_),
    .A2(_05147_),
    .B1(_05128_),
    .X(_06662_));
 sky130_fd_sc_hd__inv_2 _34616_ (.A(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__a31oi_4 _34617_ (.A1(_06660_),
    .A2(_06661_),
    .A3(_06077_),
    .B1(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand2_2 _34618_ (.A(_05998_),
    .B(_06001_),
    .Y(_06665_));
 sky130_fd_sc_hd__o21ba_2 _34619_ (.A1(net83),
    .A2(_05399_),
    .B1_N(_05280_),
    .X(_06666_));
 sky130_fd_sc_hd__and2b_1 _34620_ (.A_N(_05588_),
    .B(_05589_),
    .X(_06668_));
 sky130_fd_sc_hd__clkbuf_2 _34621_ (.A(\delay_line[36][11] ),
    .X(_06669_));
 sky130_fd_sc_hd__buf_1 _34622_ (.A(\delay_line[36][12] ),
    .X(_06670_));
 sky130_fd_sc_hd__or2b_1 _34623_ (.A(_05295_),
    .B_N(_06670_),
    .X(_06671_));
 sky130_fd_sc_hd__or2b_1 _34624_ (.A(\delay_line[36][12] ),
    .B_N(_05295_),
    .X(_06672_));
 sky130_fd_sc_hd__nor3_1 _34625_ (.A(_05298_),
    .B(_05299_),
    .C(_03688_),
    .Y(_06673_));
 sky130_fd_sc_hd__o2bb2a_1 _34626_ (.A1_N(_06671_),
    .A2_N(_06672_),
    .B1(_06673_),
    .B2(_05298_),
    .X(_06674_));
 sky130_fd_sc_hd__a21oi_1 _34627_ (.A1(_05297_),
    .A2(_05300_),
    .B1(_05298_),
    .Y(_06675_));
 sky130_fd_sc_hd__and3_1 _34628_ (.A(_06675_),
    .B(_06672_),
    .C(_06671_),
    .X(_06676_));
 sky130_fd_sc_hd__a2111oi_1 _34629_ (.A1(_06669_),
    .A2(_05302_),
    .B1(_05305_),
    .C1(_06674_),
    .D1(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__and4_1 _34630_ (.A(_06669_),
    .B(_03688_),
    .C(_03690_),
    .D(_03692_),
    .X(_06679_));
 sky130_fd_sc_hd__o22a_1 _34631_ (.A1(_06674_),
    .A2(_06676_),
    .B1(_06679_),
    .B2(_05305_),
    .X(_06680_));
 sky130_fd_sc_hd__nor3_1 _34632_ (.A(_05328_),
    .B(_05329_),
    .C(_05331_),
    .Y(_06681_));
 sky130_fd_sc_hd__xor2_1 _34633_ (.A(net299),
    .B(\delay_line[35][15] ),
    .X(_06682_));
 sky130_fd_sc_hd__or2_1 _34634_ (.A(_05320_),
    .B(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__nand2_1 _34635_ (.A(_05320_),
    .B(_06682_),
    .Y(_06684_));
 sky130_fd_sc_hd__nor3b_1 _34636_ (.A(_05313_),
    .B(_05314_),
    .C_N(_03703_),
    .Y(_06685_));
 sky130_fd_sc_hd__a221oi_1 _34637_ (.A1(_05320_),
    .A2(net299),
    .B1(_06683_),
    .B2(_06684_),
    .C1(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__inv_2 _34638_ (.A(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__o211ai_2 _34639_ (.A1(_05314_),
    .A2(_06685_),
    .B1(_06683_),
    .C1(_06684_),
    .Y(_06688_));
 sky130_fd_sc_hd__and3_1 _34640_ (.A(_06687_),
    .B(_06688_),
    .C(_05318_),
    .X(_06690_));
 sky130_fd_sc_hd__a21oi_1 _34641_ (.A1(_06687_),
    .A2(_06688_),
    .B1(_05318_),
    .Y(_06691_));
 sky130_fd_sc_hd__nor3_1 _34642_ (.A(_25098_),
    .B(_06690_),
    .C(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__o21a_1 _34643_ (.A1(_06690_),
    .A2(_06691_),
    .B1(_25098_),
    .X(_06693_));
 sky130_fd_sc_hd__nor2_1 _34644_ (.A(net226),
    .B(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__nor2_1 _34645_ (.A(_05322_),
    .B(_05325_),
    .Y(_06695_));
 sky130_fd_sc_hd__xor2_1 _34646_ (.A(_06694_),
    .B(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__o21ba_1 _34647_ (.A1(_05328_),
    .A2(_06681_),
    .B1_N(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__and3b_1 _34648_ (.A_N(_05328_),
    .B(_05333_),
    .C(_06696_),
    .X(_06698_));
 sky130_fd_sc_hd__or4_1 _34649_ (.A(net131),
    .B(_06680_),
    .C(_06697_),
    .D(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__o22ai_2 _34650_ (.A1(net129),
    .A2(_06680_),
    .B1(_06697_),
    .B2(_06698_),
    .Y(_06701_));
 sky130_fd_sc_hd__xnor2_1 _34651_ (.A(_05284_),
    .B(net291),
    .Y(_06702_));
 sky130_fd_sc_hd__and3b_1 _34652_ (.A_N(_02732_),
    .B(_05284_),
    .C(_05287_),
    .X(_06703_));
 sky130_fd_sc_hd__a21oi_1 _34653_ (.A1(_03682_),
    .A2(\delay_line[37][14] ),
    .B1(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__xnor2_2 _34654_ (.A(_06702_),
    .B(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__inv_2 _34655_ (.A(\delay_line[37][14] ),
    .Y(_06706_));
 sky130_fd_sc_hd__o22ai_2 _34656_ (.A1(_06706_),
    .A2(_05286_),
    .B1(_05290_),
    .B2(_05292_),
    .Y(_06707_));
 sky130_fd_sc_hd__xnor2_2 _34657_ (.A(_06705_),
    .B(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__a21oi_1 _34658_ (.A1(_06699_),
    .A2(_06701_),
    .B1(_06708_),
    .Y(_06709_));
 sky130_fd_sc_hd__and3_1 _34659_ (.A(_06708_),
    .B(_06699_),
    .C(_06701_),
    .X(_06710_));
 sky130_fd_sc_hd__o32ai_2 _34660_ (.A1(_05305_),
    .A2(_05310_),
    .A3(_05334_),
    .B1(_05335_),
    .B2(_05294_),
    .Y(_06712_));
 sky130_fd_sc_hd__o21ai_1 _34661_ (.A1(_06709_),
    .A2(_06710_),
    .B1(_06712_),
    .Y(_06713_));
 sky130_fd_sc_hd__or3_1 _34662_ (.A(_06709_),
    .B(_06712_),
    .C(_06710_),
    .X(_06714_));
 sky130_fd_sc_hd__nand2_2 _34663_ (.A(_06713_),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__or3b_1 _34664_ (.A(_05380_),
    .B(_05383_),
    .C_N(_05385_),
    .X(_06716_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34665_ (.A(\delay_line[38][13] ),
    .X(_06717_));
 sky130_fd_sc_hd__nor2_1 _34666_ (.A(_05380_),
    .B(_05382_),
    .Y(_06718_));
 sky130_fd_sc_hd__xor2_2 _34667_ (.A(net285),
    .B(net284),
    .X(_06719_));
 sky130_fd_sc_hd__a311oi_1 _34668_ (.A1(_02686_),
    .A2(_06717_),
    .A3(_06718_),
    .B1(_06719_),
    .C1(_05383_),
    .Y(_06720_));
 sky130_fd_sc_hd__and3_1 _34669_ (.A(_02686_),
    .B(\delay_line[38][13] ),
    .C(_06718_),
    .X(_06721_));
 sky130_fd_sc_hd__o21a_1 _34670_ (.A1(_05382_),
    .A2(_06721_),
    .B1(_06719_),
    .X(_06723_));
 sky130_fd_sc_hd__or2_1 _34671_ (.A(_06720_),
    .B(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__a21oi_1 _34672_ (.A1(_05389_),
    .A2(_06716_),
    .B1(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__and3_1 _34673_ (.A(_05389_),
    .B(_06724_),
    .C(_06716_),
    .X(_06726_));
 sky130_fd_sc_hd__nor2_1 _34674_ (.A(_06725_),
    .B(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__and2b_1 _34675_ (.A_N(_05368_),
    .B(_05371_),
    .X(_06728_));
 sky130_fd_sc_hd__a21o_1 _34676_ (.A1(_05363_),
    .A2(_05364_),
    .B1(\delay_line[39][15] ),
    .X(_06729_));
 sky130_fd_sc_hd__nand3_1 _34677_ (.A(_05363_),
    .B(_05364_),
    .C(\delay_line[39][15] ),
    .Y(_06730_));
 sky130_fd_sc_hd__a21oi_1 _34678_ (.A1(_05360_),
    .A2(_05362_),
    .B1(_05366_),
    .Y(_06731_));
 sky130_fd_sc_hd__a21oi_2 _34679_ (.A1(_06729_),
    .A2(_06730_),
    .B1(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__inv_2 _34680_ (.A(_06732_),
    .Y(_06734_));
 sky130_fd_sc_hd__nand3_1 _34681_ (.A(_06731_),
    .B(_06729_),
    .C(_06730_),
    .Y(_06735_));
 sky130_fd_sc_hd__a21oi_1 _34682_ (.A1(_06734_),
    .A2(_06735_),
    .B1(_05358_),
    .Y(_06736_));
 sky130_fd_sc_hd__and3_1 _34683_ (.A(_06734_),
    .B(_06735_),
    .C(_05358_),
    .X(_06737_));
 sky130_fd_sc_hd__nor3_1 _34684_ (.A(_06728_),
    .B(_06736_),
    .C(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__o21a_1 _34685_ (.A1(_06736_),
    .A2(_06737_),
    .B1(_06728_),
    .X(_06739_));
 sky130_fd_sc_hd__or2_1 _34686_ (.A(_06738_),
    .B(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__and3_1 _34687_ (.A(_05375_),
    .B(_05378_),
    .C(_06740_),
    .X(_06741_));
 sky130_fd_sc_hd__inv_2 _34688_ (.A(_05375_),
    .Y(_06742_));
 sky130_fd_sc_hd__nor2_1 _34689_ (.A(_06742_),
    .B(_05377_),
    .Y(_06743_));
 sky130_fd_sc_hd__nor2_1 _34690_ (.A(_06740_),
    .B(_06743_),
    .Y(_06745_));
 sky130_fd_sc_hd__nor2_1 _34691_ (.A(_06741_),
    .B(_06745_),
    .Y(_06746_));
 sky130_fd_sc_hd__nor2_1 _34692_ (.A(_06727_),
    .B(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__nand2_1 _34693_ (.A(_06727_),
    .B(_06746_),
    .Y(_06748_));
 sky130_fd_sc_hd__inv_2 _34694_ (.A(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__nor2_2 _34695_ (.A(_06747_),
    .B(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__buf_1 _34696_ (.A(\delay_line[40][14] ),
    .X(_06751_));
 sky130_fd_sc_hd__clkbuf_2 _34697_ (.A(\delay_line[40][15] ),
    .X(_06752_));
 sky130_fd_sc_hd__nor2_1 _34698_ (.A(_06751_),
    .B(_06752_),
    .Y(_06753_));
 sky130_fd_sc_hd__and2_1 _34699_ (.A(_06751_),
    .B(\delay_line[40][15] ),
    .X(_06754_));
 sky130_fd_sc_hd__a2bb2o_1 _34700_ (.A1_N(_06753_),
    .A2_N(_06754_),
    .B1(_05342_),
    .B2(_06751_),
    .X(_06756_));
 sky130_fd_sc_hd__nand2_2 _34701_ (.A(_05341_),
    .B(_06751_),
    .Y(_06757_));
 sky130_fd_sc_hd__or2_1 _34702_ (.A(_06752_),
    .B(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__and3_1 _34703_ (.A(_06756_),
    .B(_06758_),
    .C(_03659_),
    .X(_06759_));
 sky130_fd_sc_hd__a21oi_1 _34704_ (.A1(_06756_),
    .A2(_06758_),
    .B1(_03659_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_1 _34705_ (.A(_05346_),
    .B(_03658_),
    .Y(_06761_));
 sky130_fd_sc_hd__o211a_1 _34706_ (.A1(_06759_),
    .A2(_06760_),
    .B1(_05347_),
    .C1(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__a211o_1 _34707_ (.A1(_05347_),
    .A2(_06761_),
    .B1(_06759_),
    .C1(_06760_),
    .X(_06763_));
 sky130_fd_sc_hd__or2b_2 _34708_ (.A(_06762_),
    .B_N(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__o21ba_2 _34709_ (.A1(_05351_),
    .A2(_05354_),
    .B1_N(_05352_),
    .X(_06765_));
 sky130_fd_sc_hd__xor2_4 _34710_ (.A(_06764_),
    .B(_06765_),
    .X(_06767_));
 sky130_fd_sc_hd__xnor2_4 _34711_ (.A(_06750_),
    .B(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__xor2_4 _34712_ (.A(_06715_),
    .B(_06768_),
    .X(_06769_));
 sky130_fd_sc_hd__and3b_2 _34713_ (.A_N(_05451_),
    .B(_05485_),
    .C(_05453_),
    .X(_06770_));
 sky130_fd_sc_hd__and2_1 _34714_ (.A(_05165_),
    .B(_05186_),
    .X(_06771_));
 sky130_fd_sc_hd__nor2_1 _34715_ (.A(_05186_),
    .B(_05165_),
    .Y(_06772_));
 sky130_fd_sc_hd__buf_1 _34716_ (.A(_01079_),
    .X(_06773_));
 sky130_fd_sc_hd__buf_1 _34717_ (.A(_02883_),
    .X(_06774_));
 sky130_fd_sc_hd__nor2_1 _34718_ (.A(_06773_),
    .B(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__and2_1 _34719_ (.A(_06773_),
    .B(_02883_),
    .X(_06776_));
 sky130_fd_sc_hd__buf_1 _34720_ (.A(\delay_line[34][13] ),
    .X(_06778_));
 sky130_fd_sc_hd__nor2_1 _34721_ (.A(_06778_),
    .B(net303),
    .Y(_06779_));
 sky130_fd_sc_hd__and2_1 _34722_ (.A(_06778_),
    .B(net303),
    .X(_06780_));
 sky130_fd_sc_hd__and4bb_1 _34723_ (.A_N(_06779_),
    .B_N(_06780_),
    .C(_02883_),
    .D(net304),
    .X(_06781_));
 sky130_fd_sc_hd__o2bb2a_1 _34724_ (.A1_N(_06774_),
    .A2_N(net304),
    .B1(_06779_),
    .B2(_06780_),
    .X(_06782_));
 sky130_fd_sc_hd__o22ai_1 _34725_ (.A1(_06775_),
    .A2(_06776_),
    .B1(_06781_),
    .B2(_06782_),
    .Y(_06783_));
 sky130_fd_sc_hd__or4_1 _34726_ (.A(_06775_),
    .B(_06776_),
    .C(_06781_),
    .D(_06782_),
    .X(_06784_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34727_ (.A(_05166_),
    .X(_06785_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34728_ (.A(_06778_),
    .X(_06786_));
 sky130_fd_sc_hd__o211a_1 _34729_ (.A1(_06785_),
    .A2(_05167_),
    .B1(_06773_),
    .C1(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__a211oi_1 _34730_ (.A1(_06783_),
    .A2(_06784_),
    .B1(_06787_),
    .C1(_05171_),
    .Y(_06789_));
 sky130_fd_sc_hd__o211a_1 _34731_ (.A1(_06787_),
    .A2(_05171_),
    .B1(_06783_),
    .C1(_06784_),
    .X(_06790_));
 sky130_fd_sc_hd__nor4_1 _34732_ (.A(_06771_),
    .B(_06772_),
    .C(_06789_),
    .D(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__o22a_1 _34733_ (.A1(_06771_),
    .A2(_06772_),
    .B1(_06789_),
    .B2(_06790_),
    .X(_06792_));
 sky130_fd_sc_hd__a211o_1 _34734_ (.A1(_05173_),
    .A2(_05176_),
    .B1(net225),
    .C1(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__o221ai_1 _34735_ (.A1(_05175_),
    .A2(_05177_),
    .B1(_06792_),
    .B2(net225),
    .C1(_05173_),
    .Y(_06794_));
 sky130_fd_sc_hd__and2_1 _34736_ (.A(_06793_),
    .B(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__xnor2_1 _34737_ (.A(_05162_),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__and3_1 _34738_ (.A(_05181_),
    .B(_05182_),
    .C(_06796_),
    .X(_06797_));
 sky130_fd_sc_hd__a21oi_1 _34739_ (.A1(_05181_),
    .A2(_05182_),
    .B1(_06796_),
    .Y(_06798_));
 sky130_fd_sc_hd__or2_1 _34740_ (.A(_06797_),
    .B(_06798_),
    .X(_06800_));
 sky130_fd_sc_hd__nand2_1 _34741_ (.A(_05188_),
    .B(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__nand2_1 _34742_ (.A(_05185_),
    .B(_05188_),
    .Y(_06802_));
 sky130_fd_sc_hd__nor2_1 _34743_ (.A(_03759_),
    .B(_03763_),
    .Y(_06803_));
 sky130_fd_sc_hd__o21a_1 _34744_ (.A1(_06802_),
    .A2(_06803_),
    .B1(_05188_),
    .X(_06804_));
 sky130_fd_sc_hd__nor2_1 _34745_ (.A(_06800_),
    .B(_06804_),
    .Y(_06805_));
 sky130_fd_sc_hd__o21bai_1 _34746_ (.A1(_05189_),
    .A2(_06801_),
    .B1_N(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__o211ai_1 _34747_ (.A1(_05236_),
    .A2(_05239_),
    .B1(_05259_),
    .C1(_05261_),
    .Y(_06807_));
 sky130_fd_sc_hd__nand2_1 _34748_ (.A(_05261_),
    .B(_06807_),
    .Y(_06808_));
 sky130_fd_sc_hd__a2bb2o_1 _34749_ (.A1_N(_05251_),
    .A2_N(_05255_),
    .B1(_02836_),
    .B2(_23358_),
    .X(_06809_));
 sky130_fd_sc_hd__or3b_1 _34750_ (.A(_20666_),
    .B(_24922_),
    .C_N(_05242_),
    .X(_06811_));
 sky130_fd_sc_hd__clkbuf_2 _34751_ (.A(_05241_),
    .X(_06812_));
 sky130_fd_sc_hd__a21o_1 _34752_ (.A1(_06812_),
    .A2(_05242_),
    .B1(_02848_),
    .X(_06813_));
 sky130_fd_sc_hd__and4_1 _34753_ (.A(_03780_),
    .B(_06811_),
    .C(_02840_),
    .D(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__inv_2 _34754_ (.A(_06814_),
    .Y(_06815_));
 sky130_fd_sc_hd__a22o_1 _34755_ (.A1(_05237_),
    .A2(_03780_),
    .B1(_06811_),
    .B2(_06813_),
    .X(_06816_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34756_ (.A(\delay_line[33][11] ),
    .X(_06817_));
 sky130_fd_sc_hd__xnor2_1 _34757_ (.A(_24922_),
    .B(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__or2_1 _34758_ (.A(net309),
    .B(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__nand2_1 _34759_ (.A(net309),
    .B(_06818_),
    .Y(_06820_));
 sky130_fd_sc_hd__a21bo_1 _34760_ (.A1(_06819_),
    .A2(_06820_),
    .B1_N(_05246_),
    .X(_06822_));
 sky130_fd_sc_hd__nand3b_1 _34761_ (.A_N(_05246_),
    .B(_06819_),
    .C(_06820_),
    .Y(_06823_));
 sky130_fd_sc_hd__and4_1 _34762_ (.A(_06815_),
    .B(_06816_),
    .C(_06822_),
    .D(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__a22oi_1 _34763_ (.A1(_06815_),
    .A2(_06816_),
    .B1(_06822_),
    .B2(_06823_),
    .Y(_06825_));
 sky130_fd_sc_hd__o32a_1 _34764_ (.A1(_03775_),
    .A2(_05245_),
    .A3(_05246_),
    .B1(_05247_),
    .B2(_05256_),
    .X(_06826_));
 sky130_fd_sc_hd__o21ai_1 _34765_ (.A1(_06824_),
    .A2(_06825_),
    .B1(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__nor3_1 _34766_ (.A(_06826_),
    .B(_06824_),
    .C(_06825_),
    .Y(_06828_));
 sky130_fd_sc_hd__inv_2 _34767_ (.A(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__and3_1 _34768_ (.A(_06809_),
    .B(_06827_),
    .C(_06829_),
    .X(_06830_));
 sky130_fd_sc_hd__a21o_1 _34769_ (.A1(_06827_),
    .A2(_06829_),
    .B1(_06809_),
    .X(_06831_));
 sky130_fd_sc_hd__and2b_1 _34770_ (.A_N(_06830_),
    .B(_06831_),
    .X(_06833_));
 sky130_fd_sc_hd__xnor2_1 _34771_ (.A(_06808_),
    .B(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__nor2_1 _34772_ (.A(_05267_),
    .B(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__and2_1 _34773_ (.A(_05267_),
    .B(_06834_),
    .X(_06836_));
 sky130_fd_sc_hd__nor2_1 _34774_ (.A(_06835_),
    .B(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__o21ai_2 _34775_ (.A1(_05269_),
    .A2(_05270_),
    .B1(_05266_),
    .Y(_06838_));
 sky130_fd_sc_hd__xnor2_1 _34776_ (.A(_06837_),
    .B(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__nand2_1 _34777_ (.A(_02805_),
    .B(_21126_),
    .Y(_06840_));
 sky130_fd_sc_hd__and3_1 _34778_ (.A(_05212_),
    .B(_06840_),
    .C(_24971_),
    .X(_06841_));
 sky130_fd_sc_hd__buf_2 _34779_ (.A(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__o2bb2a_1 _34780_ (.A1_N(_24971_),
    .A2_N(_06840_),
    .B1(_03826_),
    .B2(_05211_),
    .X(_06844_));
 sky130_fd_sc_hd__nand3_1 _34781_ (.A(_05202_),
    .B(_05206_),
    .C(_05207_),
    .Y(_06845_));
 sky130_fd_sc_hd__and2_1 _34782_ (.A(\delay_line[32][13] ),
    .B(\delay_line[32][15] ),
    .X(_06846_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34783_ (.A(\delay_line[32][15] ),
    .X(_06847_));
 sky130_fd_sc_hd__nor2_1 _34784_ (.A(_03811_),
    .B(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__o21a_1 _34785_ (.A1(_06846_),
    .A2(_06848_),
    .B1(_05196_),
    .X(_06849_));
 sky130_fd_sc_hd__nor3_1 _34786_ (.A(_05196_),
    .B(_06846_),
    .C(_06848_),
    .Y(_06850_));
 sky130_fd_sc_hd__o2bb2a_1 _34787_ (.A1_N(_05197_),
    .A2_N(_05198_),
    .B1(_06849_),
    .B2(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__inv_2 _34788_ (.A(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__nand2_1 _34789_ (.A(_05197_),
    .B(_05198_),
    .Y(_06853_));
 sky130_fd_sc_hd__or3_1 _34790_ (.A(_06849_),
    .B(_06850_),
    .C(_06853_),
    .X(_06855_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34791_ (.A(_03809_),
    .X(_06856_));
 sky130_fd_sc_hd__and3_1 _34792_ (.A(_06852_),
    .B(_06855_),
    .C(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__a21oi_1 _34793_ (.A1(_06852_),
    .A2(_06855_),
    .B1(_06856_),
    .Y(_06858_));
 sky130_fd_sc_hd__a211oi_2 _34794_ (.A1(_05202_),
    .A2(_06845_),
    .B1(_06857_),
    .C1(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__o211a_1 _34795_ (.A1(_06857_),
    .A2(_06858_),
    .B1(_05202_),
    .C1(_06845_),
    .X(_06860_));
 sky130_fd_sc_hd__or4_1 _34796_ (.A(_06842_),
    .B(_06844_),
    .C(_06859_),
    .D(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__o22ai_2 _34797_ (.A1(_06842_),
    .A2(_06844_),
    .B1(_06859_),
    .B2(_06860_),
    .Y(_06862_));
 sky130_fd_sc_hd__a211oi_2 _34798_ (.A1(_06861_),
    .A2(_06862_),
    .B1(_05210_),
    .C1(net169),
    .Y(_06863_));
 sky130_fd_sc_hd__o211ai_2 _34799_ (.A1(_05210_),
    .A2(net169),
    .B1(_06861_),
    .C1(_06862_),
    .Y(_06864_));
 sky130_fd_sc_hd__inv_2 _34800_ (.A(_06864_),
    .Y(_06866_));
 sky130_fd_sc_hd__nor3_1 _34801_ (.A(_05214_),
    .B(_06863_),
    .C(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__o21a_1 _34802_ (.A1(_06863_),
    .A2(_06866_),
    .B1(_05214_),
    .X(_06868_));
 sky130_fd_sc_hd__o21ai_1 _34803_ (.A1(_03823_),
    .A2(_03831_),
    .B1(_05223_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand4_2 _34804_ (.A(_03824_),
    .B(_05224_),
    .C(_03825_),
    .D(_02815_),
    .Y(_06870_));
 sky130_fd_sc_hd__o211a_1 _34805_ (.A1(_06867_),
    .A2(_06868_),
    .B1(_06869_),
    .C1(_06870_),
    .X(_06871_));
 sky130_fd_sc_hd__a211oi_1 _34806_ (.A1(_06869_),
    .A2(_06870_),
    .B1(_06867_),
    .C1(_06868_),
    .Y(_06872_));
 sky130_fd_sc_hd__nor2_1 _34807_ (.A(_06871_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__xor2_2 _34808_ (.A(_05228_),
    .B(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__a311o_1 _34809_ (.A1(_02826_),
    .A2(_02817_),
    .A3(_03837_),
    .B1(_05225_),
    .C1(_03836_),
    .X(_06875_));
 sky130_fd_sc_hd__inv_2 _34810_ (.A(_05228_),
    .Y(_06877_));
 sky130_fd_sc_hd__a21boi_1 _34811_ (.A1(_06875_),
    .A2(_06877_),
    .B1_N(_03844_),
    .Y(_06878_));
 sky130_fd_sc_hd__a21o_1 _34812_ (.A1(_03841_),
    .A2(_03844_),
    .B1(_03808_),
    .X(_06879_));
 sky130_fd_sc_hd__a22oi_2 _34813_ (.A1(_03841_),
    .A2(_03808_),
    .B1(_03807_),
    .B2(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__and3b_1 _34814_ (.A_N(_03844_),
    .B(_06875_),
    .C(_06877_),
    .X(_06881_));
 sky130_fd_sc_hd__o21bai_2 _34815_ (.A1(_06878_),
    .A2(_06880_),
    .B1_N(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__xnor2_2 _34816_ (.A(_06874_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__and2_1 _34817_ (.A(_06839_),
    .B(_06883_),
    .X(_06884_));
 sky130_fd_sc_hd__nor2_1 _34818_ (.A(_06839_),
    .B(_06883_),
    .Y(_06885_));
 sky130_fd_sc_hd__nor2_1 _34819_ (.A(_06884_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__xnor2_1 _34820_ (.A(_06806_),
    .B(_06886_),
    .Y(_06888_));
 sky130_fd_sc_hd__o21a_1 _34821_ (.A1(_06770_),
    .A2(_05487_),
    .B1(_06888_),
    .X(_06889_));
 sky130_fd_sc_hd__nor3_1 _34822_ (.A(_06770_),
    .B(_05487_),
    .C(_06888_),
    .Y(_06890_));
 sky130_fd_sc_hd__nor2_1 _34823_ (.A(_06889_),
    .B(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__or2b_1 _34824_ (.A(_05191_),
    .B_N(_05273_),
    .X(_06892_));
 sky130_fd_sc_hd__o21ai_2 _34825_ (.A1(_05235_),
    .A2(_05272_),
    .B1(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__xor2_1 _34826_ (.A(_06891_),
    .B(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__inv_2 _34827_ (.A(_05277_),
    .Y(_06895_));
 sky130_fd_sc_hd__o21ai_1 _34828_ (.A1(_05276_),
    .A2(_06895_),
    .B1(_05275_),
    .Y(_06896_));
 sky130_fd_sc_hd__nand2_1 _34829_ (.A(_06894_),
    .B(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__or2_1 _34830_ (.A(_06896_),
    .B(_06894_),
    .X(_06899_));
 sky130_fd_sc_hd__and2_1 _34831_ (.A(_06897_),
    .B(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__xnor2_1 _34832_ (.A(_06769_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__o21bai_1 _34833_ (.A1(_05586_),
    .A2(_06668_),
    .B1_N(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__or3b_1 _34834_ (.A(_05586_),
    .B(_06668_),
    .C_N(_06901_),
    .X(_06903_));
 sky130_fd_sc_hd__nand2_2 _34835_ (.A(_06902_),
    .B(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__xnor2_4 _34836_ (.A(_06666_),
    .B(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__o32a_4 _34837_ (.A1(_05487_),
    .A2(_05488_),
    .A3(_05584_),
    .B1(_05583_),
    .B2(_05492_),
    .X(_06906_));
 sky130_fd_sc_hd__or3_1 _34838_ (.A(_05463_),
    .B(_05466_),
    .C(_05462_),
    .X(_06907_));
 sky130_fd_sc_hd__xor2_2 _34839_ (.A(_04378_),
    .B(_04383_),
    .X(_06908_));
 sky130_fd_sc_hd__and2b_1 _34840_ (.A_N(net319),
    .B(_06908_),
    .X(_06910_));
 sky130_fd_sc_hd__and2b_1 _34841_ (.A_N(_06908_),
    .B(net319),
    .X(_06911_));
 sky130_fd_sc_hd__o211ai_1 _34842_ (.A1(_06910_),
    .A2(_06911_),
    .B1(_05459_),
    .C1(_05455_),
    .Y(_06912_));
 sky130_fd_sc_hd__a211o_1 _34843_ (.A1(_05459_),
    .A2(_05455_),
    .B1(_06910_),
    .C1(_06911_),
    .X(_06913_));
 sky130_fd_sc_hd__and3_1 _34844_ (.A(_02089_),
    .B(_02102_),
    .C(_02099_),
    .X(_06914_));
 sky130_fd_sc_hd__a211oi_1 _34845_ (.A1(_05476_),
    .A2(_02099_),
    .B1(_02103_),
    .C1(_02107_),
    .Y(_06915_));
 sky130_fd_sc_hd__or4_2 _34846_ (.A(_19336_),
    .B(_06914_),
    .C(_23246_),
    .D(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__a2bb2o_1 _34847_ (.A1_N(_06915_),
    .A2_N(_06914_),
    .B1(_20350_),
    .B2(_04399_),
    .X(_06917_));
 sky130_fd_sc_hd__and4_1 _34848_ (.A(_06912_),
    .B(_06913_),
    .C(_06916_),
    .D(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34849_ (.A(_06912_),
    .X(_06919_));
 sky130_fd_sc_hd__a22oi_2 _34850_ (.A1(_06919_),
    .A2(_06913_),
    .B1(_06916_),
    .B2(_06917_),
    .Y(_06921_));
 sky130_fd_sc_hd__a211oi_2 _34851_ (.A1(_05461_),
    .A2(_06907_),
    .B1(_06918_),
    .C1(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__o221a_1 _34852_ (.A1(_05463_),
    .A2(_05466_),
    .B1(_06921_),
    .B2(_06918_),
    .C1(_05461_),
    .X(_06923_));
 sky130_fd_sc_hd__buf_1 _34853_ (.A(_04378_),
    .X(_06924_));
 sky130_fd_sc_hd__buf_1 _34854_ (.A(_06924_),
    .X(_06925_));
 sky130_fd_sc_hd__o2bb2a_1 _34855_ (.A1_N(_06925_),
    .A2_N(_02092_),
    .B1(_24394_),
    .B2(_05464_),
    .X(_06926_));
 sky130_fd_sc_hd__o21a_1 _34856_ (.A1(_06922_),
    .A2(_06923_),
    .B1(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__nor3_1 _34857_ (.A(_06926_),
    .B(_06922_),
    .C(_06923_),
    .Y(_06928_));
 sky130_fd_sc_hd__or2_1 _34858_ (.A(_06927_),
    .B(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__or3b_1 _34859_ (.A(_05472_),
    .B(_05474_),
    .C_N(_06929_),
    .X(_06930_));
 sky130_fd_sc_hd__o21bai_2 _34860_ (.A1(_05472_),
    .A2(_05474_),
    .B1_N(_06929_),
    .Y(_06932_));
 sky130_fd_sc_hd__and2_1 _34861_ (.A(_06930_),
    .B(_06932_),
    .X(_06933_));
 sky130_fd_sc_hd__inv_2 _34862_ (.A(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__and3_1 _34863_ (.A(_05481_),
    .B(_04403_),
    .C(_05479_),
    .X(_06935_));
 sky130_fd_sc_hd__a21oi_1 _34864_ (.A1(_05484_),
    .A2(_05483_),
    .B1(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__or2_1 _34865_ (.A(_06934_),
    .B(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__a221o_1 _34866_ (.A1(_06930_),
    .A2(_06932_),
    .B1(_05484_),
    .B2(_05483_),
    .C1(_06935_),
    .X(_06938_));
 sky130_fd_sc_hd__a21oi_1 _34867_ (.A1(_06937_),
    .A2(_06938_),
    .B1(_05479_),
    .Y(_06939_));
 sky130_fd_sc_hd__and3_1 _34868_ (.A(_05479_),
    .B(_06937_),
    .C(_06938_),
    .X(_06940_));
 sky130_fd_sc_hd__buf_1 _34869_ (.A(\delay_line[29][13] ),
    .X(_06941_));
 sky130_fd_sc_hd__or2b_1 _34870_ (.A(net321),
    .B_N(_06941_),
    .X(_06943_));
 sky130_fd_sc_hd__or2b_1 _34871_ (.A(\delay_line[29][13] ),
    .B_N(\delay_line[29][9] ),
    .X(_06944_));
 sky130_fd_sc_hd__and2_1 _34872_ (.A(_06943_),
    .B(_06944_),
    .X(_06945_));
 sky130_fd_sc_hd__a21oi_1 _34873_ (.A1(_04408_),
    .A2(_05448_),
    .B1(_05445_),
    .Y(_06946_));
 sky130_fd_sc_hd__xor2_1 _34874_ (.A(_06945_),
    .B(_06946_),
    .X(_06947_));
 sky130_fd_sc_hd__or4bb_1 _34875_ (.A(_05445_),
    .B(_05446_),
    .C_N(_04407_),
    .D_N(_04411_),
    .X(_06948_));
 sky130_fd_sc_hd__and3_1 _34876_ (.A(_05453_),
    .B(_06947_),
    .C(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__a21oi_1 _34877_ (.A1(_05453_),
    .A2(_06948_),
    .B1(_06947_),
    .Y(_06950_));
 sky130_fd_sc_hd__nor2_1 _34878_ (.A(_06949_),
    .B(_06950_),
    .Y(_06951_));
 sky130_fd_sc_hd__o21ai_1 _34879_ (.A1(_06939_),
    .A2(_06940_),
    .B1(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__or3_1 _34880_ (.A(_06951_),
    .B(_06939_),
    .C(_06940_),
    .X(_06954_));
 sky130_fd_sc_hd__o211a_1 _34881_ (.A1(_04365_),
    .A2(_04368_),
    .B1(_05435_),
    .C1(_05437_),
    .X(_06955_));
 sky130_fd_sc_hd__o21bai_1 _34882_ (.A1(_04348_),
    .A2(_05434_),
    .B1_N(_05433_),
    .Y(_06956_));
 sky130_fd_sc_hd__clkbuf_2 _34883_ (.A(_23207_),
    .X(_06957_));
 sky130_fd_sc_hd__nand2_1 _34884_ (.A(_06957_),
    .B(_20313_),
    .Y(_06958_));
 sky130_fd_sc_hd__and4b_1 _34885_ (.A_N(_02144_),
    .B(_23214_),
    .C(_06958_),
    .D(_21264_),
    .X(_06959_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34886_ (.A(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__o2bb2a_1 _34887_ (.A1_N(_23214_),
    .A2_N(_06958_),
    .B1(_02144_),
    .B2(_05423_),
    .X(_06961_));
 sky130_fd_sc_hd__and2b_1 _34888_ (.A_N(_04351_),
    .B(_05409_),
    .X(_06962_));
 sky130_fd_sc_hd__o21ai_2 _34889_ (.A1(_05415_),
    .A2(_06962_),
    .B1(_05410_),
    .Y(_06963_));
 sky130_fd_sc_hd__xor2_2 _34890_ (.A(\delay_line[31][15] ),
    .B(_06963_),
    .X(_06965_));
 sky130_fd_sc_hd__a2111o_1 _34891_ (.A1(_05412_),
    .A2(_05416_),
    .B1(_04352_),
    .C1(_05417_),
    .D1(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__nand2_1 _34892_ (.A(_05419_),
    .B(_06965_),
    .Y(_06967_));
 sky130_fd_sc_hd__nand2_1 _34893_ (.A(_06966_),
    .B(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__o21ai_1 _34894_ (.A1(_06960_),
    .A2(_06961_),
    .B1(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__or3_1 _34895_ (.A(_06960_),
    .B(_06961_),
    .C(_06968_),
    .X(_06970_));
 sky130_fd_sc_hd__a211o_1 _34896_ (.A1(_06969_),
    .A2(_06970_),
    .B1(_05430_),
    .C1(_05431_),
    .X(_06971_));
 sky130_fd_sc_hd__o211ai_2 _34897_ (.A1(_05430_),
    .A2(_05431_),
    .B1(_06969_),
    .C1(_06970_),
    .Y(_06972_));
 sky130_fd_sc_hd__nand3_1 _34898_ (.A(_06971_),
    .B(_06972_),
    .C(_05426_),
    .Y(_06973_));
 sky130_fd_sc_hd__a32o_1 _34899_ (.A1(_04346_),
    .A2(_05422_),
    .A3(_05424_),
    .B1(_06971_),
    .B2(_06972_),
    .X(_06974_));
 sky130_fd_sc_hd__and2_1 _34900_ (.A(_06973_),
    .B(_06974_),
    .X(_06976_));
 sky130_fd_sc_hd__or2_1 _34901_ (.A(_06956_),
    .B(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__nand2_1 _34902_ (.A(_06976_),
    .B(_06956_),
    .Y(_06978_));
 sky130_fd_sc_hd__and2_1 _34903_ (.A(_06977_),
    .B(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__o21bai_2 _34904_ (.A1(_05442_),
    .A2(_05443_),
    .B1_N(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__o21bai_2 _34905_ (.A1(_05442_),
    .A2(_05443_),
    .B1_N(_05440_),
    .Y(_06981_));
 sky130_fd_sc_hd__xor2_1 _34906_ (.A(_06979_),
    .B(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__nor2_1 _34907_ (.A(_06955_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__a21oi_2 _34908_ (.A1(_06955_),
    .A2(_06980_),
    .B1(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__a21oi_2 _34909_ (.A1(_06952_),
    .A2(_06954_),
    .B1(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__o311a_1 _34910_ (.A1(_06951_),
    .A2(_06939_),
    .A3(_06940_),
    .B1(_06984_),
    .C1(_06952_),
    .X(_06987_));
 sky130_fd_sc_hd__o21a_1 _34911_ (.A1(_05582_),
    .A2(_05553_),
    .B1(_05552_),
    .X(_06988_));
 sky130_fd_sc_hd__buf_1 _34912_ (.A(_05560_),
    .X(_06989_));
 sky130_fd_sc_hd__nor2_1 _34913_ (.A(_06989_),
    .B(_05559_),
    .Y(_06990_));
 sky130_fd_sc_hd__o21ai_1 _34914_ (.A1(_05565_),
    .A2(_06990_),
    .B1(_05564_),
    .Y(_06991_));
 sky130_fd_sc_hd__inv_2 _34915_ (.A(\delay_line[28][15] ),
    .Y(_06992_));
 sky130_fd_sc_hd__nor2_1 _34916_ (.A(_06989_),
    .B(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__and3b_1 _34917_ (.A_N(_05561_),
    .B(_06992_),
    .C(_05560_),
    .X(_06994_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34918_ (.A(\delay_line[28][15] ),
    .X(_06995_));
 sky130_fd_sc_hd__and3_1 _34919_ (.A(_05561_),
    .B(_05560_),
    .C(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__o31a_1 _34920_ (.A1(_06993_),
    .A2(_06994_),
    .A3(_06996_),
    .B1(_01031_),
    .X(_06998_));
 sky130_fd_sc_hd__buf_1 _34921_ (.A(_05561_),
    .X(_06999_));
 sky130_fd_sc_hd__a2111oi_1 _34922_ (.A1(_06999_),
    .A2(_06995_),
    .B1(_06993_),
    .C1(_06994_),
    .D1(_01031_),
    .Y(_07000_));
 sky130_fd_sc_hd__or3_2 _34923_ (.A(_06991_),
    .B(_06998_),
    .C(net267),
    .X(_07001_));
 sky130_fd_sc_hd__o21ai_1 _34924_ (.A1(_06998_),
    .A2(net266),
    .B1(_06991_),
    .Y(_07002_));
 sky130_fd_sc_hd__a21o_1 _34925_ (.A1(_07001_),
    .A2(_07002_),
    .B1(_05565_),
    .X(_07003_));
 sky130_fd_sc_hd__nand3_2 _34926_ (.A(_07001_),
    .B(_07002_),
    .C(_05565_),
    .Y(_07004_));
 sky130_fd_sc_hd__o211a_1 _34927_ (.A1(_05569_),
    .A2(_05571_),
    .B1(_07003_),
    .C1(_07004_),
    .X(_07005_));
 sky130_fd_sc_hd__a211oi_1 _34928_ (.A1(_07003_),
    .A2(_07004_),
    .B1(_05569_),
    .C1(_05571_),
    .Y(_07006_));
 sky130_fd_sc_hd__nor4_1 _34929_ (.A(_07005_),
    .B(_05573_),
    .C(_05574_),
    .D(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__o22a_1 _34930_ (.A1(_07005_),
    .A2(_07006_),
    .B1(_05573_),
    .B2(_05574_),
    .X(_07009_));
 sky130_fd_sc_hd__nor2_1 _34931_ (.A(_07007_),
    .B(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__a21o_1 _34932_ (.A1(_04281_),
    .A2(_05575_),
    .B1(_05581_),
    .X(_07011_));
 sky130_fd_sc_hd__xnor2_1 _34933_ (.A(_07010_),
    .B(_07011_),
    .Y(_07012_));
 sky130_fd_sc_hd__clkbuf_2 _34934_ (.A(_05531_),
    .X(_07013_));
 sky130_fd_sc_hd__a32oi_2 _34935_ (.A1(_02203_),
    .A2(_04301_),
    .A3(_05540_),
    .B1(_05542_),
    .B2(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__inv_2 _34936_ (.A(net334),
    .Y(_07015_));
 sky130_fd_sc_hd__nor2_1 _34937_ (.A(net337),
    .B(_00994_),
    .Y(_07016_));
 sky130_fd_sc_hd__and2_1 _34938_ (.A(net337),
    .B(\delay_line[26][10] ),
    .X(_07017_));
 sky130_fd_sc_hd__or3b_2 _34939_ (.A(_07016_),
    .B(_07017_),
    .C_N(_20397_),
    .X(_07018_));
 sky130_fd_sc_hd__o21bai_1 _34940_ (.A1(_07016_),
    .A2(_07017_),
    .B1_N(_20397_),
    .Y(_07020_));
 sky130_fd_sc_hd__nand2_1 _34941_ (.A(_07018_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__a21oi_1 _34942_ (.A1(_05533_),
    .A2(_05534_),
    .B1(_07021_),
    .Y(_07022_));
 sky130_fd_sc_hd__and3_1 _34943_ (.A(_05533_),
    .B(_05534_),
    .C(_07021_),
    .X(_07023_));
 sky130_fd_sc_hd__nor2_1 _34944_ (.A(_07022_),
    .B(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__a21oi_1 _34945_ (.A1(_04298_),
    .A2(_05540_),
    .B1(_05538_),
    .Y(_07025_));
 sky130_fd_sc_hd__xor2_1 _34946_ (.A(_07024_),
    .B(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__xor2_1 _34947_ (.A(_07015_),
    .B(_07026_),
    .X(_07027_));
 sky130_fd_sc_hd__and2b_1 _34948_ (.A_N(_07014_),
    .B(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__and2b_1 _34949_ (.A_N(_07027_),
    .B(_07014_),
    .X(_07029_));
 sky130_fd_sc_hd__nor2_1 _34950_ (.A(_07028_),
    .B(_07029_),
    .Y(_07031_));
 sky130_fd_sc_hd__o21bai_1 _34951_ (.A1(_05547_),
    .A2(_05550_),
    .B1_N(_05544_),
    .Y(_07032_));
 sky130_fd_sc_hd__xnor2_1 _34952_ (.A(_07031_),
    .B(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__nand2_1 _34953_ (.A(_04315_),
    .B(net329),
    .Y(_07034_));
 sky130_fd_sc_hd__inv_2 _34954_ (.A(net329),
    .Y(_07035_));
 sky130_fd_sc_hd__nand2_1 _34955_ (.A(_07035_),
    .B(_04318_),
    .Y(_07036_));
 sky130_fd_sc_hd__and3_1 _34956_ (.A(_05496_),
    .B(_07034_),
    .C(_07036_),
    .X(_07037_));
 sky130_fd_sc_hd__a21oi_1 _34957_ (.A1(_07034_),
    .A2(_07036_),
    .B1(_05496_),
    .Y(_07038_));
 sky130_fd_sc_hd__or2_1 _34958_ (.A(_07037_),
    .B(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__clkbuf_2 _34959_ (.A(_07035_),
    .X(_07040_));
 sky130_fd_sc_hd__mux2_1 _34960_ (.A0(_07039_),
    .A1(_07040_),
    .S(_05497_),
    .X(_07042_));
 sky130_fd_sc_hd__or2_1 _34961_ (.A(_23157_),
    .B(_07042_),
    .X(_07043_));
 sky130_fd_sc_hd__nand2_1 _34962_ (.A(_23157_),
    .B(_07042_),
    .Y(_07044_));
 sky130_fd_sc_hd__and3_1 _34963_ (.A(_05504_),
    .B(_21241_),
    .C(_05505_),
    .X(_07045_));
 sky130_fd_sc_hd__a211oi_2 _34964_ (.A1(_07043_),
    .A2(_07044_),
    .B1(_05503_),
    .C1(_07045_),
    .Y(_07046_));
 sky130_fd_sc_hd__o211ai_2 _34965_ (.A1(_05503_),
    .A2(_07045_),
    .B1(_07043_),
    .C1(_07044_),
    .Y(_07047_));
 sky130_fd_sc_hd__inv_2 _34966_ (.A(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__nor3_1 _34967_ (.A(_07046_),
    .B(_05505_),
    .C(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__o32a_1 _34968_ (.A1(_20378_),
    .A2(_21237_),
    .A3(_21240_),
    .B1(_07048_),
    .B2(_07046_),
    .X(_07050_));
 sky130_fd_sc_hd__o221a_1 _34969_ (.A1(_23147_),
    .A2(_05515_),
    .B1(_07049_),
    .B2(_07050_),
    .C1(_05514_),
    .X(_07051_));
 sky130_fd_sc_hd__or4_1 _34970_ (.A(_19276_),
    .B(_20375_),
    .C(_20376_),
    .D(_05515_),
    .X(_07053_));
 sky130_fd_sc_hd__a211o_1 _34971_ (.A1(_05514_),
    .A2(_07053_),
    .B1(_07049_),
    .C1(_07050_),
    .X(_07054_));
 sky130_fd_sc_hd__inv_2 _34972_ (.A(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__a2111oi_1 _34973_ (.A1(_05493_),
    .A2(_05494_),
    .B1(_05516_),
    .C1(_07051_),
    .D1(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__o21a_1 _34974_ (.A1(_07051_),
    .A2(_07055_),
    .B1(_05518_),
    .X(_07057_));
 sky130_fd_sc_hd__nor2_1 _34975_ (.A(net127),
    .B(_07057_),
    .Y(_07058_));
 sky130_fd_sc_hd__a21oi_1 _34976_ (.A1(_05522_),
    .A2(_05523_),
    .B1(_05520_),
    .Y(_07059_));
 sky130_fd_sc_hd__xor2_1 _34977_ (.A(_07058_),
    .B(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__xnor2_1 _34978_ (.A(_07033_),
    .B(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__nand2_1 _34979_ (.A(_07012_),
    .B(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__or2_1 _34980_ (.A(_07012_),
    .B(_07061_),
    .X(_07064_));
 sky130_fd_sc_hd__nand2_1 _34981_ (.A(_07062_),
    .B(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__xor2_1 _34982_ (.A(_06988_),
    .B(_07065_),
    .X(_07066_));
 sky130_fd_sc_hd__or3b_1 _34983_ (.A(_06985_),
    .B(_06987_),
    .C_N(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__o21bai_1 _34984_ (.A1(_06985_),
    .A2(_06987_),
    .B1_N(_07066_),
    .Y(_07068_));
 sky130_fd_sc_hd__and2_2 _34985_ (.A(_07067_),
    .B(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__a21o_1 _34986_ (.A1(_05985_),
    .A2(_05860_),
    .B1(_05984_),
    .X(_07070_));
 sky130_fd_sc_hd__and2_1 _34987_ (.A(_07069_),
    .B(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__nor2_1 _34988_ (.A(_07070_),
    .B(_07069_),
    .Y(_07072_));
 sky130_fd_sc_hd__nor3_1 _34989_ (.A(_06906_),
    .B(_07071_),
    .C(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__o21a_1 _34990_ (.A1(_07071_),
    .A2(_07072_),
    .B1(_06906_),
    .X(_07075_));
 sky130_fd_sc_hd__o21a_1 _34991_ (.A1(_04158_),
    .A2(_05895_),
    .B1(_05896_),
    .X(_07076_));
 sky130_fd_sc_hd__nor2_1 _34992_ (.A(_05892_),
    .B(_05893_),
    .Y(_07077_));
 sky130_fd_sc_hd__nand2_1 _34993_ (.A(_20484_),
    .B(_05888_),
    .Y(_07078_));
 sky130_fd_sc_hd__a21bo_1 _34994_ (.A1(_05871_),
    .A2(_05870_),
    .B1_N(_05866_),
    .X(_07079_));
 sky130_fd_sc_hd__or2_2 _34995_ (.A(_05868_),
    .B(\delay_line[25][15] ),
    .X(_07080_));
 sky130_fd_sc_hd__buf_1 _34996_ (.A(\delay_line[25][15] ),
    .X(_07081_));
 sky130_fd_sc_hd__nand2_2 _34997_ (.A(_05868_),
    .B(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__inv_2 _34998_ (.A(_05862_),
    .Y(_07083_));
 sky130_fd_sc_hd__inv_2 _34999_ (.A(net340),
    .Y(_07084_));
 sky130_fd_sc_hd__o2bb2ai_1 _35000_ (.A1_N(_07080_),
    .A2_N(_07082_),
    .B1(_07083_),
    .B2(_07084_),
    .Y(_07086_));
 sky130_fd_sc_hd__nand4_1 _35001_ (.A(_07080_),
    .B(_07082_),
    .C(_05862_),
    .D(_05863_),
    .Y(_07087_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35002_ (.A(_24511_),
    .X(_07088_));
 sky130_fd_sc_hd__a21o_1 _35003_ (.A1(_07086_),
    .A2(_07087_),
    .B1(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__nand3_1 _35004_ (.A(_07087_),
    .B(_07088_),
    .C(_07086_),
    .Y(_07090_));
 sky130_fd_sc_hd__nand3_1 _35005_ (.A(_07079_),
    .B(_07089_),
    .C(_07090_),
    .Y(_07091_));
 sky130_fd_sc_hd__buf_1 _35006_ (.A(_07091_),
    .X(_07092_));
 sky130_fd_sc_hd__a21o_1 _35007_ (.A1(_07089_),
    .A2(_07090_),
    .B1(_07079_),
    .X(_07093_));
 sky130_fd_sc_hd__or3b_1 _35008_ (.A(_21561_),
    .B(_21566_),
    .C_N(_05880_),
    .X(_07094_));
 sky130_fd_sc_hd__o21a_1 _35009_ (.A1(_05880_),
    .A2(_05878_),
    .B1(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__a21oi_1 _35010_ (.A1(_07092_),
    .A2(_07093_),
    .B1(_07095_),
    .Y(_07097_));
 sky130_fd_sc_hd__a32oi_4 _35011_ (.A1(_05872_),
    .A2(_05873_),
    .A3(_05875_),
    .B1(_05879_),
    .B2(_05882_),
    .Y(_07098_));
 sky130_fd_sc_hd__a31o_1 _35012_ (.A1(_07092_),
    .A2(_07093_),
    .A3(_07095_),
    .B1(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__and3_1 _35013_ (.A(_07092_),
    .B(_07093_),
    .C(_07095_),
    .X(_07100_));
 sky130_fd_sc_hd__o21ai_1 _35014_ (.A1(_07100_),
    .A2(_07097_),
    .B1(_07098_),
    .Y(_07101_));
 sky130_fd_sc_hd__o21ai_1 _35015_ (.A1(_07097_),
    .A2(_07099_),
    .B1(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__xnor2_1 _35016_ (.A(_07078_),
    .B(_07102_),
    .Y(_07103_));
 sky130_fd_sc_hd__xor2_2 _35017_ (.A(_07077_),
    .B(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__xor2_2 _35018_ (.A(_05890_),
    .B(_07104_),
    .X(_07105_));
 sky130_fd_sc_hd__xor2_2 _35019_ (.A(_07076_),
    .B(_07105_),
    .X(_07106_));
 sky130_fd_sc_hd__o21bai_2 _35020_ (.A1(_05900_),
    .A2(_05902_),
    .B1_N(_05903_),
    .Y(_07108_));
 sky130_fd_sc_hd__xnor2_2 _35021_ (.A(_07106_),
    .B(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__or4b_1 _35022_ (.A(_17106_),
    .B(_18318_),
    .C(_05932_),
    .D_N(_06887_),
    .X(_07110_));
 sky130_fd_sc_hd__a21oi_1 _35023_ (.A1(_05918_),
    .A2(_05919_),
    .B1(_05921_),
    .Y(_07111_));
 sky130_fd_sc_hd__o21ai_1 _35024_ (.A1(_20454_),
    .A2(_17095_),
    .B1(_18318_),
    .Y(_07112_));
 sky130_fd_sc_hd__buf_1 _35025_ (.A(_21599_),
    .X(_07113_));
 sky130_fd_sc_hd__and3_1 _35026_ (.A(_07113_),
    .B(_20454_),
    .C(_18317_),
    .X(_07114_));
 sky130_fd_sc_hd__buf_1 _35027_ (.A(_02363_),
    .X(_07115_));
 sky130_fd_sc_hd__a21o_1 _35028_ (.A1(_00517_),
    .A2(_20450_),
    .B1(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__or3b_1 _35029_ (.A(_00512_),
    .B(_07113_),
    .C_N(_02363_),
    .X(_07117_));
 sky130_fd_sc_hd__inv_2 _35030_ (.A(net351),
    .Y(_07119_));
 sky130_fd_sc_hd__nand2_1 _35031_ (.A(_02367_),
    .B(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35032_ (.A(\delay_line[22][13] ),
    .X(_07121_));
 sky130_fd_sc_hd__nand2_1 _35033_ (.A(_00518_),
    .B(net351),
    .Y(_07122_));
 sky130_fd_sc_hd__nand4_2 _35034_ (.A(_07120_),
    .B(_07121_),
    .C(_00514_),
    .D(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__a22o_1 _35035_ (.A1(_00514_),
    .A2(_07121_),
    .B1(_07122_),
    .B2(_07120_),
    .X(_07124_));
 sky130_fd_sc_hd__nand4_2 _35036_ (.A(_07116_),
    .B(_07117_),
    .C(_07123_),
    .D(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__a22o_1 _35037_ (.A1(_07116_),
    .A2(_07117_),
    .B1(_07123_),
    .B2(_07124_),
    .X(_07126_));
 sky130_fd_sc_hd__nand2_1 _35038_ (.A(_05915_),
    .B(_05918_),
    .Y(_07127_));
 sky130_fd_sc_hd__a21oi_2 _35039_ (.A1(_07125_),
    .A2(_07126_),
    .B1(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__and3_1 _35040_ (.A(_07127_),
    .B(_07125_),
    .C(_07126_),
    .X(_07130_));
 sky130_fd_sc_hd__o22a_1 _35041_ (.A1(_00517_),
    .A2(_07114_),
    .B1(_07128_),
    .B2(_07130_),
    .X(_07131_));
 sky130_fd_sc_hd__clkbuf_2 _35042_ (.A(_07113_),
    .X(_07132_));
 sky130_fd_sc_hd__a2111oi_4 _35043_ (.A1(_07132_),
    .A2(_18318_),
    .B1(_00517_),
    .C1(_07128_),
    .D1(_07130_),
    .Y(_07133_));
 sky130_fd_sc_hd__o221a_1 _35044_ (.A1(_07111_),
    .A2(_07112_),
    .B1(_07131_),
    .B2(_07133_),
    .C1(_05924_),
    .X(_07134_));
 sky130_fd_sc_hd__or3b_1 _35045_ (.A(_07112_),
    .B(_07111_),
    .C_N(_05924_),
    .X(_07135_));
 sky130_fd_sc_hd__a211oi_2 _35046_ (.A1(_05924_),
    .A2(_07135_),
    .B1(_07133_),
    .C1(_07131_),
    .Y(_07136_));
 sky130_fd_sc_hd__nor3_2 _35047_ (.A(_05923_),
    .B(_07134_),
    .C(_07136_),
    .Y(_07137_));
 sky130_fd_sc_hd__o32a_1 _35048_ (.A1(_17106_),
    .A2(_04174_),
    .A3(_20454_),
    .B1(_07134_),
    .B2(_07136_),
    .X(_07138_));
 sky130_fd_sc_hd__a211oi_2 _35049_ (.A1(_05930_),
    .A2(_07110_),
    .B1(_07137_),
    .C1(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__o221a_1 _35050_ (.A1(_04192_),
    .A2(_05932_),
    .B1(_07137_),
    .B2(_07138_),
    .C1(_05930_),
    .X(_07141_));
 sky130_fd_sc_hd__nor2_1 _35051_ (.A(_07139_),
    .B(_07141_),
    .Y(_07142_));
 sky130_fd_sc_hd__or2b_1 _35052_ (.A(_05907_),
    .B_N(_05933_),
    .X(_07143_));
 sky130_fd_sc_hd__o21ai_1 _35053_ (.A1(_05934_),
    .A2(_05935_),
    .B1(_07143_),
    .Y(_07144_));
 sky130_fd_sc_hd__nor2_1 _35054_ (.A(_07142_),
    .B(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__and2_1 _35055_ (.A(_07144_),
    .B(_07142_),
    .X(_07146_));
 sky130_fd_sc_hd__or3_1 _35056_ (.A(_02336_),
    .B(_04211_),
    .C(_04207_),
    .X(_07147_));
 sky130_fd_sc_hd__o21ai_1 _35057_ (.A1(_04211_),
    .A2(_04207_),
    .B1(_02336_),
    .Y(_07148_));
 sky130_fd_sc_hd__nand2_1 _35058_ (.A(_07147_),
    .B(_07148_),
    .Y(_07149_));
 sky130_fd_sc_hd__and3_1 _35059_ (.A(_05949_),
    .B(_05950_),
    .C(_05951_),
    .X(_07150_));
 sky130_fd_sc_hd__and3_1 _35060_ (.A(_05952_),
    .B(_05956_),
    .C(_05959_),
    .X(_07152_));
 sky130_fd_sc_hd__buf_1 _35061_ (.A(\delay_line[24][11] ),
    .X(_07153_));
 sky130_fd_sc_hd__nor2_1 _35062_ (.A(_00559_),
    .B(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__and2_1 _35063_ (.A(\delay_line[24][10] ),
    .B(_07153_),
    .X(_07155_));
 sky130_fd_sc_hd__o21bai_1 _35064_ (.A1(_07154_),
    .A2(_07155_),
    .B1_N(_24583_),
    .Y(_07156_));
 sky130_fd_sc_hd__nand2_1 _35065_ (.A(_00551_),
    .B(_02317_),
    .Y(_07157_));
 sky130_fd_sc_hd__nand3b_1 _35066_ (.A_N(_07154_),
    .B(_07157_),
    .C(_24583_),
    .Y(_07158_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35067_ (.A(\delay_line[24][14] ),
    .X(_07159_));
 sky130_fd_sc_hd__nand3_1 _35068_ (.A(_07156_),
    .B(_07158_),
    .C(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__a21o_1 _35069_ (.A1(_07156_),
    .A2(_07158_),
    .B1(_07159_),
    .X(_07161_));
 sky130_fd_sc_hd__nand3_1 _35070_ (.A(_05954_),
    .B(_07160_),
    .C(_07161_),
    .Y(_07163_));
 sky130_fd_sc_hd__clkbuf_2 _35071_ (.A(_05947_),
    .X(_07164_));
 sky130_fd_sc_hd__a32o_1 _35072_ (.A1(_07164_),
    .A2(_05943_),
    .A3(_05946_),
    .B1(_07160_),
    .B2(_07161_),
    .X(_07165_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35073_ (.A(_05957_),
    .X(_07166_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35074_ (.A(_00560_),
    .X(_07167_));
 sky130_fd_sc_hd__a21oi_1 _35075_ (.A1(_07166_),
    .A2(_07167_),
    .B1(_22891_),
    .Y(_07168_));
 sky130_fd_sc_hd__o21a_1 _35076_ (.A1(_05957_),
    .A2(_07167_),
    .B1(_22891_),
    .X(_07169_));
 sky130_fd_sc_hd__o2bb2ai_1 _35077_ (.A1_N(_07163_),
    .A2_N(_07165_),
    .B1(_07168_),
    .B2(_07169_),
    .Y(_07170_));
 sky130_fd_sc_hd__clkbuf_2 _35078_ (.A(_22891_),
    .X(_07171_));
 sky130_fd_sc_hd__o2111ai_2 _35079_ (.A1(_07171_),
    .A2(_05944_),
    .B1(_05941_),
    .C1(_07163_),
    .D1(_07165_),
    .Y(_07172_));
 sky130_fd_sc_hd__o211ai_1 _35080_ (.A1(_07150_),
    .A2(_07152_),
    .B1(_07170_),
    .C1(_07172_),
    .Y(_07174_));
 sky130_fd_sc_hd__a211o_1 _35081_ (.A1(_07170_),
    .A2(_07172_),
    .B1(_07150_),
    .C1(_07152_),
    .X(_07175_));
 sky130_fd_sc_hd__nand2_1 _35082_ (.A(_07174_),
    .B(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__xnor2_1 _35083_ (.A(_07149_),
    .B(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__a21oi_1 _35084_ (.A1(_05963_),
    .A2(_05966_),
    .B1(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__and3_1 _35085_ (.A(_05963_),
    .B(_05966_),
    .C(_07177_),
    .X(_07179_));
 sky130_fd_sc_hd__o32a_2 _35086_ (.A1(_22876_),
    .A2(_02318_),
    .A3(_22871_),
    .B1(_07178_),
    .B2(_07179_),
    .X(_07180_));
 sky130_fd_sc_hd__a211o_1 _35087_ (.A1(_05963_),
    .A2(_07177_),
    .B1(_05938_),
    .C1(_07178_),
    .X(_07181_));
 sky130_fd_sc_hd__inv_2 _35088_ (.A(_07181_),
    .Y(_07182_));
 sky130_fd_sc_hd__a21o_1 _35089_ (.A1(_05970_),
    .A2(_05971_),
    .B1(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__o211a_1 _35090_ (.A1(_07182_),
    .A2(_07180_),
    .B1(_05970_),
    .C1(_05971_),
    .X(_07185_));
 sky130_fd_sc_hd__o21bai_1 _35091_ (.A1(_07180_),
    .A2(_07183_),
    .B1_N(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__and3_1 _35092_ (.A(_05937_),
    .B(_05971_),
    .C(_05973_),
    .X(_07187_));
 sky130_fd_sc_hd__a21oi_2 _35093_ (.A1(_05977_),
    .A2(_05976_),
    .B1(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__xnor2_1 _35094_ (.A(_07186_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__nor3_1 _35095_ (.A(_07145_),
    .B(_07146_),
    .C(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__o21a_1 _35096_ (.A1(_07145_),
    .A2(_07146_),
    .B1(_07189_),
    .X(_07191_));
 sky130_fd_sc_hd__or2_1 _35097_ (.A(_07190_),
    .B(_07191_),
    .X(_07192_));
 sky130_fd_sc_hd__nor2_1 _35098_ (.A(_07109_),
    .B(_07192_),
    .Y(_07193_));
 sky130_fd_sc_hd__nand2_1 _35099_ (.A(_07109_),
    .B(_07192_),
    .Y(_07194_));
 sky130_fd_sc_hd__or2b_1 _35100_ (.A(_07193_),
    .B_N(_07194_),
    .X(_07196_));
 sky130_fd_sc_hd__a21oi_1 _35101_ (.A1(_05725_),
    .A2(_05729_),
    .B1(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__and3_1 _35102_ (.A(_05725_),
    .B(_05729_),
    .C(_07196_),
    .X(_07198_));
 sky130_fd_sc_hd__a21bo_1 _35103_ (.A1(_05905_),
    .A2(_05980_),
    .B1_N(_05979_),
    .X(_07199_));
 sky130_fd_sc_hd__o21ba_1 _35104_ (.A1(_07197_),
    .A2(_07198_),
    .B1_N(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__or3b_1 _35105_ (.A(_07197_),
    .B(_07198_),
    .C_N(_07199_),
    .X(_07201_));
 sky130_fd_sc_hd__or2b_4 _35106_ (.A(_07200_),
    .B_N(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__o211a_1 _35107_ (.A1(_05752_),
    .A2(_05754_),
    .B1(_03901_),
    .C1(_05756_),
    .X(_07203_));
 sky130_fd_sc_hd__nor2_1 _35108_ (.A(_03901_),
    .B(_05758_),
    .Y(_07204_));
 sky130_fd_sc_hd__nand2_1 _35109_ (.A(_05749_),
    .B(_05760_),
    .Y(_07205_));
 sky130_fd_sc_hd__nor2_1 _35110_ (.A(_00828_),
    .B(_02489_),
    .Y(_07207_));
 sky130_fd_sc_hd__and2_1 _35111_ (.A(net382),
    .B(net381),
    .X(_07208_));
 sky130_fd_sc_hd__o21ai_1 _35112_ (.A1(_07207_),
    .A2(_07208_),
    .B1(_05739_),
    .Y(_07209_));
 sky130_fd_sc_hd__inv_2 _35113_ (.A(\delay_line[16][11] ),
    .Y(_07210_));
 sky130_fd_sc_hd__nand2_1 _35114_ (.A(_02497_),
    .B(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__nand3b_1 _35115_ (.A_N(_07208_),
    .B(_05753_),
    .C(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__a21o_1 _35116_ (.A1(_07209_),
    .A2(_07212_),
    .B1(net380),
    .X(_07213_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35117_ (.A(net380),
    .X(_07214_));
 sky130_fd_sc_hd__nand3_1 _35118_ (.A(_07212_),
    .B(_07214_),
    .C(_07209_),
    .Y(_07215_));
 sky130_fd_sc_hd__nand3_1 _35119_ (.A(_07213_),
    .B(_05746_),
    .C(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__a32o_1 _35120_ (.A1(_05747_),
    .A2(_05741_),
    .A3(_05743_),
    .B1(_07215_),
    .B2(_07213_),
    .X(_07218_));
 sky130_fd_sc_hd__o21ai_1 _35121_ (.A1(_05753_),
    .A2(_00834_),
    .B1(_23026_),
    .Y(_07219_));
 sky130_fd_sc_hd__o21a_1 _35122_ (.A1(_05752_),
    .A2(_05738_),
    .B1(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__a21o_1 _35123_ (.A1(_07216_),
    .A2(_07218_),
    .B1(_07220_),
    .X(_07221_));
 sky130_fd_sc_hd__o2111ai_2 _35124_ (.A1(_05752_),
    .A2(_05738_),
    .B1(_07216_),
    .C1(_07218_),
    .D1(_07219_),
    .Y(_07222_));
 sky130_fd_sc_hd__nand3_2 _35125_ (.A(_07205_),
    .B(_07221_),
    .C(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__a21o_1 _35126_ (.A1(_07221_),
    .A2(_07222_),
    .B1(_07205_),
    .X(_07224_));
 sky130_fd_sc_hd__and4bb_1 _35127_ (.A_N(_07203_),
    .B_N(_07204_),
    .C(_07223_),
    .D(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__a2bb2oi_1 _35128_ (.A1_N(_07203_),
    .A2_N(_07204_),
    .B1(_07223_),
    .B2(_07224_),
    .Y(_07226_));
 sky130_fd_sc_hd__a211o_1 _35129_ (.A1(_05761_),
    .A2(_05763_),
    .B1(_07225_),
    .C1(_07226_),
    .X(_07227_));
 sky130_fd_sc_hd__nand2_1 _35130_ (.A(_05759_),
    .B(_05760_),
    .Y(_07229_));
 sky130_fd_sc_hd__o31a_1 _35131_ (.A1(_02500_),
    .A2(_03883_),
    .A3(_03886_),
    .B1(_03896_),
    .X(_07230_));
 sky130_fd_sc_hd__o221ai_2 _35132_ (.A1(_07229_),
    .A2(_07230_),
    .B1(_07226_),
    .B2(_07225_),
    .C1(_05763_),
    .Y(_07231_));
 sky130_fd_sc_hd__nand4_1 _35133_ (.A(_07227_),
    .B(_03875_),
    .C(_03913_),
    .D(_07231_),
    .Y(_07232_));
 sky130_fd_sc_hd__inv_2 _35134_ (.A(_07232_),
    .Y(_07233_));
 sky130_fd_sc_hd__a22oi_1 _35135_ (.A1(_03913_),
    .A2(_03875_),
    .B1(_07231_),
    .B2(_07227_),
    .Y(_07234_));
 sky130_fd_sc_hd__inv_2 _35136_ (.A(_05769_),
    .Y(_07235_));
 sky130_fd_sc_hd__o211a_1 _35137_ (.A1(_07233_),
    .A2(_07234_),
    .B1(_05768_),
    .C1(_07235_),
    .X(_07236_));
 sky130_fd_sc_hd__a211o_1 _35138_ (.A1(_05768_),
    .A2(_07235_),
    .B1(_07233_),
    .C1(_07234_),
    .X(_07237_));
 sky130_fd_sc_hd__or2b_2 _35139_ (.A(_07236_),
    .B_N(_07237_),
    .X(_07238_));
 sky130_fd_sc_hd__o21ai_2 _35140_ (.A1(_05847_),
    .A2(_05848_),
    .B1(_03917_),
    .Y(_07240_));
 sky130_fd_sc_hd__a211oi_2 _35141_ (.A1(_03911_),
    .A2(_03912_),
    .B1(_05769_),
    .C1(_05770_),
    .Y(_07241_));
 sky130_fd_sc_hd__a21oi_4 _35142_ (.A1(_07240_),
    .A2(_05772_),
    .B1(_07241_),
    .Y(_07242_));
 sky130_fd_sc_hd__xnor2_4 _35143_ (.A(_07238_),
    .B(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__o21ai_1 _35144_ (.A1(_03981_),
    .A2(_05836_),
    .B1(_05837_),
    .Y(_07244_));
 sky130_fd_sc_hd__and3_1 _35145_ (.A(_05803_),
    .B(_05822_),
    .C(_05827_),
    .X(_07245_));
 sky130_fd_sc_hd__buf_1 _35146_ (.A(_05801_),
    .X(_07246_));
 sky130_fd_sc_hd__o21ai_1 _35147_ (.A1(_05824_),
    .A2(_05825_),
    .B1(_05817_),
    .Y(_07247_));
 sky130_fd_sc_hd__a21bo_1 _35148_ (.A1(_05811_),
    .A2(_05813_),
    .B1_N(_05808_),
    .X(_07248_));
 sky130_fd_sc_hd__buf_1 _35149_ (.A(\delay_line[15][15] ),
    .X(_07249_));
 sky130_fd_sc_hd__nor2_2 _35150_ (.A(_03954_),
    .B(_07249_),
    .Y(_07251_));
 sky130_fd_sc_hd__and2_1 _35151_ (.A(_03954_),
    .B(\delay_line[15][15] ),
    .X(_07252_));
 sky130_fd_sc_hd__nor3_2 _35152_ (.A(_05807_),
    .B(_07251_),
    .C(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__inv_2 _35153_ (.A(_03957_),
    .Y(_07254_));
 sky130_fd_sc_hd__inv_2 _35154_ (.A(\delay_line[15][14] ),
    .Y(_07255_));
 sky130_fd_sc_hd__o22a_1 _35155_ (.A1(_07254_),
    .A2(_07255_),
    .B1(_07251_),
    .B2(_07252_),
    .X(_07256_));
 sky130_fd_sc_hd__or3b_1 _35156_ (.A(_07253_),
    .B(_07256_),
    .C_N(_24745_),
    .X(_07257_));
 sky130_fd_sc_hd__nor2_1 _35157_ (.A(_07253_),
    .B(_07256_),
    .Y(_07258_));
 sky130_fd_sc_hd__or2_1 _35158_ (.A(_24745_),
    .B(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__nand3_1 _35159_ (.A(_07248_),
    .B(_07257_),
    .C(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__a21o_1 _35160_ (.A1(_07257_),
    .A2(_07259_),
    .B1(_07248_),
    .X(_07262_));
 sky130_fd_sc_hd__or2_1 _35161_ (.A(_05819_),
    .B(_03960_),
    .X(_07263_));
 sky130_fd_sc_hd__o31a_1 _35162_ (.A1(_21455_),
    .A2(_05823_),
    .A3(_21451_),
    .B1(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__and3_1 _35163_ (.A(_07260_),
    .B(_07262_),
    .C(_07264_),
    .X(_07265_));
 sky130_fd_sc_hd__a21oi_1 _35164_ (.A1(_07260_),
    .A2(_07262_),
    .B1(_07264_),
    .Y(_07266_));
 sky130_fd_sc_hd__a211o_1 _35165_ (.A1(_05826_),
    .A2(_07247_),
    .B1(_07265_),
    .C1(_07266_),
    .X(_07267_));
 sky130_fd_sc_hd__o211ai_2 _35166_ (.A1(_07265_),
    .A2(_07266_),
    .B1(_05826_),
    .C1(_07247_),
    .Y(_07268_));
 sky130_fd_sc_hd__o2111ai_2 _35167_ (.A1(_21454_),
    .A2(_05819_),
    .B1(_07246_),
    .C1(_07267_),
    .D1(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__a22o_1 _35168_ (.A1(_07246_),
    .A2(_20597_),
    .B1(_07268_),
    .B2(_07267_),
    .X(_07270_));
 sky130_fd_sc_hd__o211a_1 _35169_ (.A1(_07245_),
    .A2(_05835_),
    .B1(_07269_),
    .C1(_07270_),
    .X(_07271_));
 sky130_fd_sc_hd__a211oi_1 _35170_ (.A1(_07269_),
    .A2(_07270_),
    .B1(_07245_),
    .C1(_05835_),
    .Y(_07273_));
 sky130_fd_sc_hd__or3_1 _35171_ (.A(_07271_),
    .B(_05802_),
    .C(_07273_),
    .X(_07274_));
 sky130_fd_sc_hd__o21ai_1 _35172_ (.A1(_07273_),
    .A2(_07271_),
    .B1(_05802_),
    .Y(_07275_));
 sky130_fd_sc_hd__nand3_1 _35173_ (.A(_07244_),
    .B(_07274_),
    .C(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__a21o_1 _35174_ (.A1(_07274_),
    .A2(_07275_),
    .B1(_07244_),
    .X(_07277_));
 sky130_fd_sc_hd__and2_1 _35175_ (.A(_07276_),
    .B(_07277_),
    .X(_07278_));
 sky130_fd_sc_hd__and2b_1 _35176_ (.A_N(_05839_),
    .B(_05840_),
    .X(_07279_));
 sky130_fd_sc_hd__o21bai_1 _35177_ (.A1(_05841_),
    .A2(_05842_),
    .B1_N(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__nor2_1 _35178_ (.A(_07278_),
    .B(_07280_),
    .Y(_07281_));
 sky130_fd_sc_hd__inv_2 _35179_ (.A(_07281_),
    .Y(_07282_));
 sky130_fd_sc_hd__or2_1 _35180_ (.A(_05775_),
    .B(_05793_),
    .X(_07284_));
 sky130_fd_sc_hd__buf_1 _35181_ (.A(_23054_),
    .X(_07285_));
 sky130_fd_sc_hd__buf_1 _35182_ (.A(_24783_),
    .X(_07286_));
 sky130_fd_sc_hd__a21oi_1 _35183_ (.A1(_07285_),
    .A2(_07286_),
    .B1(_03922_),
    .Y(_07287_));
 sky130_fd_sc_hd__and3_1 _35184_ (.A(_03922_),
    .B(_07285_),
    .C(_07286_),
    .X(_07288_));
 sky130_fd_sc_hd__nor2_1 _35185_ (.A(_07286_),
    .B(_00749_),
    .Y(_07289_));
 sky130_fd_sc_hd__and2_1 _35186_ (.A(_24783_),
    .B(\delay_line[14][10] ),
    .X(_07290_));
 sky130_fd_sc_hd__or3b_1 _35187_ (.A(_07289_),
    .B(_07290_),
    .C_N(net389),
    .X(_07291_));
 sky130_fd_sc_hd__o21bai_1 _35188_ (.A1(_07289_),
    .A2(_07290_),
    .B1_N(net389),
    .Y(_07292_));
 sky130_fd_sc_hd__clkbuf_2 _35189_ (.A(\delay_line[14][13] ),
    .X(_07293_));
 sky130_fd_sc_hd__nor2_1 _35190_ (.A(_05779_),
    .B(_05780_),
    .Y(_07295_));
 sky130_fd_sc_hd__and4_1 _35191_ (.A(_07291_),
    .B(_07292_),
    .C(_07293_),
    .D(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__a22oi_1 _35192_ (.A1(_07293_),
    .A2(_07295_),
    .B1(_07291_),
    .B2(_07292_),
    .Y(_07297_));
 sky130_fd_sc_hd__or4_1 _35193_ (.A(_07287_),
    .B(_07288_),
    .C(_07296_),
    .D(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__o22ai_1 _35194_ (.A1(_07287_),
    .A2(_07288_),
    .B1(_07296_),
    .B2(_07297_),
    .Y(_07299_));
 sky130_fd_sc_hd__nand2_1 _35195_ (.A(_07298_),
    .B(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__o311a_1 _35196_ (.A1(_05776_),
    .A2(_05787_),
    .A3(_05784_),
    .B1(_07300_),
    .C1(_05783_),
    .X(_07301_));
 sky130_fd_sc_hd__inv_2 _35197_ (.A(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__a21o_1 _35198_ (.A1(_05783_),
    .A2(_05786_),
    .B1(_07300_),
    .X(_07303_));
 sky130_fd_sc_hd__and3_1 _35199_ (.A(_07302_),
    .B(_07303_),
    .C(_05787_),
    .X(_07304_));
 sky130_fd_sc_hd__a21oi_1 _35200_ (.A1(_07302_),
    .A2(_07303_),
    .B1(_05787_),
    .Y(_07306_));
 sky130_fd_sc_hd__a211oi_2 _35201_ (.A1(_05792_),
    .A2(_07284_),
    .B1(_07304_),
    .C1(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__o221a_1 _35202_ (.A1(_05775_),
    .A2(_05793_),
    .B1(_07304_),
    .B2(_07306_),
    .C1(_05792_),
    .X(_07308_));
 sky130_fd_sc_hd__a21oi_1 _35203_ (.A1(_05798_),
    .A2(_05797_),
    .B1(_05796_),
    .Y(_07309_));
 sky130_fd_sc_hd__nor3_1 _35204_ (.A(_07307_),
    .B(_07308_),
    .C(_07309_),
    .Y(_07310_));
 sky130_fd_sc_hd__o21a_1 _35205_ (.A1(_07307_),
    .A2(_07308_),
    .B1(_07309_),
    .X(_07311_));
 sky130_fd_sc_hd__nor2_1 _35206_ (.A(_07310_),
    .B(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand2_1 _35207_ (.A(_07280_),
    .B(_07278_),
    .Y(_07313_));
 sky130_fd_sc_hd__and3_1 _35208_ (.A(_07282_),
    .B(_07312_),
    .C(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__a21oi_1 _35209_ (.A1(_07313_),
    .A2(_07282_),
    .B1(_07312_),
    .Y(_07315_));
 sky130_fd_sc_hd__nor2_1 _35210_ (.A(_07314_),
    .B(_07315_),
    .Y(_07317_));
 sky130_fd_sc_hd__xor2_4 _35211_ (.A(_07243_),
    .B(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__a21oi_1 _35212_ (.A1(_05800_),
    .A2(_05844_),
    .B1(_05846_),
    .Y(_07319_));
 sky130_fd_sc_hd__nand2_1 _35213_ (.A(_07318_),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__or2_1 _35214_ (.A(_07319_),
    .B(_07318_),
    .X(_07321_));
 sky130_fd_sc_hd__or2_1 _35215_ (.A(_05595_),
    .B(_05638_),
    .X(_07322_));
 sky130_fd_sc_hd__or3b_1 _35216_ (.A(_05597_),
    .B(_05599_),
    .C_N(_05628_),
    .X(_07323_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35217_ (.A(_04089_),
    .X(_07324_));
 sky130_fd_sc_hd__a21o_1 _35218_ (.A1(_18350_),
    .A2(_07324_),
    .B1(_05598_),
    .X(_07325_));
 sky130_fd_sc_hd__o21a_1 _35219_ (.A1(_05616_),
    .A2(_05619_),
    .B1(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__inv_2 _35220_ (.A(_05613_),
    .Y(_07328_));
 sky130_fd_sc_hd__buf_1 _35221_ (.A(\delay_line[21][14] ),
    .X(_07329_));
 sky130_fd_sc_hd__nor2_1 _35222_ (.A(_05600_),
    .B(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__and2_1 _35223_ (.A(\delay_line[21][13] ),
    .B(\delay_line[21][14] ),
    .X(_07331_));
 sky130_fd_sc_hd__a211oi_2 _35224_ (.A1(_04103_),
    .A2(_05605_),
    .B1(_07330_),
    .C1(_07331_),
    .Y(_07332_));
 sky130_fd_sc_hd__and3_2 _35225_ (.A(_04103_),
    .B(_05600_),
    .C(_07329_),
    .X(_07333_));
 sky130_fd_sc_hd__or3_2 _35226_ (.A(_24635_),
    .B(_07332_),
    .C(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__o21ai_2 _35227_ (.A1(_07332_),
    .A2(_07333_),
    .B1(_24635_),
    .Y(_07335_));
 sky130_fd_sc_hd__buf_1 _35228_ (.A(_05605_),
    .X(_07336_));
 sky130_fd_sc_hd__nor2_1 _35229_ (.A(_07336_),
    .B(_05606_),
    .Y(_07337_));
 sky130_fd_sc_hd__a221o_1 _35230_ (.A1(_05609_),
    .A2(_05604_),
    .B1(_07334_),
    .B2(_07335_),
    .C1(_07337_),
    .X(_07339_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35231_ (.A(_22986_),
    .X(_07340_));
 sky130_fd_sc_hd__buf_1 _35232_ (.A(_22987_),
    .X(_07341_));
 sky130_fd_sc_hd__or3b_1 _35233_ (.A(_07340_),
    .B(_07341_),
    .C_N(_21423_),
    .X(_07342_));
 sky130_fd_sc_hd__nor2_1 _35234_ (.A(_22986_),
    .B(_07341_),
    .Y(_07343_));
 sky130_fd_sc_hd__or2_1 _35235_ (.A(_04089_),
    .B(_07343_),
    .X(_07344_));
 sky130_fd_sc_hd__a21oi_1 _35236_ (.A1(_04090_),
    .A2(_05616_),
    .B1(_05614_),
    .Y(_07345_));
 sky130_fd_sc_hd__a21oi_1 _35237_ (.A1(_07342_),
    .A2(_07344_),
    .B1(_07345_),
    .Y(_07346_));
 sky130_fd_sc_hd__and3_1 _35238_ (.A(_07345_),
    .B(_07342_),
    .C(_07344_),
    .X(_07347_));
 sky130_fd_sc_hd__nor2_1 _35239_ (.A(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35240_ (.A(_04100_),
    .X(_07350_));
 sky130_fd_sc_hd__nor2_2 _35241_ (.A(_05602_),
    .B(_05603_),
    .Y(_07351_));
 sky130_fd_sc_hd__o21a_1 _35242_ (.A1(_07350_),
    .A2(_07351_),
    .B1(_22992_),
    .X(_07352_));
 sky130_fd_sc_hd__o211ai_2 _35243_ (.A1(_07337_),
    .A2(_07352_),
    .B1(_07334_),
    .C1(_07335_),
    .Y(_07353_));
 sky130_fd_sc_hd__nand3_1 _35244_ (.A(_07339_),
    .B(_07348_),
    .C(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__a21o_1 _35245_ (.A1(_07353_),
    .A2(_07339_),
    .B1(_07348_),
    .X(_07355_));
 sky130_fd_sc_hd__o2111a_1 _35246_ (.A1(_05622_),
    .A2(_07328_),
    .B1(_07354_),
    .C1(_07355_),
    .D1(_05611_),
    .X(_07356_));
 sky130_fd_sc_hd__o21ai_1 _35247_ (.A1(_05622_),
    .A2(_07328_),
    .B1(_05611_),
    .Y(_07357_));
 sky130_fd_sc_hd__nand2_1 _35248_ (.A(_07354_),
    .B(_07355_),
    .Y(_07358_));
 sky130_fd_sc_hd__and2_1 _35249_ (.A(_07357_),
    .B(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__or3_1 _35250_ (.A(_07326_),
    .B(_07356_),
    .C(_07359_),
    .X(_07361_));
 sky130_fd_sc_hd__o21ai_1 _35251_ (.A1(_07356_),
    .A2(_07359_),
    .B1(_07326_),
    .Y(_07362_));
 sky130_fd_sc_hd__a22oi_2 _35252_ (.A1(_05629_),
    .A2(_07323_),
    .B1(_07361_),
    .B2(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand4_2 _35253_ (.A(_05629_),
    .B(_07323_),
    .C(_07361_),
    .D(_07362_),
    .Y(_07364_));
 sky130_fd_sc_hd__and4b_1 _35254_ (.A_N(_07363_),
    .B(_05597_),
    .C(_18351_),
    .D(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__inv_2 _35255_ (.A(_07364_),
    .Y(_07366_));
 sky130_fd_sc_hd__o2bb2a_1 _35256_ (.A1_N(_18351_),
    .A2_N(_05597_),
    .B1(_07366_),
    .B2(_07363_),
    .X(_07367_));
 sky130_fd_sc_hd__a211oi_1 _35257_ (.A1(_05637_),
    .A2(_07322_),
    .B1(_07365_),
    .C1(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__o221a_1 _35258_ (.A1(_05595_),
    .A2(_05638_),
    .B1(_07365_),
    .B2(_07367_),
    .C1(_05637_),
    .X(_07369_));
 sky130_fd_sc_hd__or2_2 _35259_ (.A(_07368_),
    .B(_07369_),
    .X(_07370_));
 sky130_fd_sc_hd__o21a_1 _35260_ (.A1(_05593_),
    .A2(_04121_),
    .B1(_05639_),
    .X(_07372_));
 sky130_fd_sc_hd__a21oi_4 _35261_ (.A1(_05641_),
    .A2(_05640_),
    .B1(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__xnor2_4 _35262_ (.A(_07370_),
    .B(_07373_),
    .Y(_07374_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35263_ (.A(_19395_),
    .X(_07375_));
 sky130_fd_sc_hd__clkbuf_2 _35264_ (.A(_21356_),
    .X(_07376_));
 sky130_fd_sc_hd__and3_1 _35265_ (.A(_07376_),
    .B(_21354_),
    .C(_18385_),
    .X(_07377_));
 sky130_fd_sc_hd__buf_1 _35266_ (.A(_21358_),
    .X(_07378_));
 sky130_fd_sc_hd__a21o_1 _35267_ (.A1(_19394_),
    .A2(_20542_),
    .B1(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__or3b_1 _35268_ (.A(_19390_),
    .B(_21356_),
    .C_N(_21363_),
    .X(_07380_));
 sky130_fd_sc_hd__clkbuf_2 _35269_ (.A(\delay_line[18][14] ),
    .X(_07381_));
 sky130_fd_sc_hd__nor2_1 _35270_ (.A(net373),
    .B(_07381_),
    .Y(_07383_));
 sky130_fd_sc_hd__and2_1 _35271_ (.A(net373),
    .B(\delay_line[18][14] ),
    .X(_07384_));
 sky130_fd_sc_hd__or3_1 _35272_ (.A(_07383_),
    .B(_05648_),
    .C(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__o21ai_1 _35273_ (.A1(_07384_),
    .A2(_07383_),
    .B1(_05648_),
    .Y(_07386_));
 sky130_fd_sc_hd__nand4_1 _35274_ (.A(_07379_),
    .B(_07380_),
    .C(_07385_),
    .D(_07386_),
    .Y(_07387_));
 sky130_fd_sc_hd__a22o_1 _35275_ (.A1(_07379_),
    .A2(_07380_),
    .B1(_07385_),
    .B2(_07386_),
    .X(_07388_));
 sky130_fd_sc_hd__a21o_1 _35276_ (.A1(_05654_),
    .A2(_05651_),
    .B1(net277),
    .X(_07389_));
 sky130_fd_sc_hd__a21oi_1 _35277_ (.A1(_07387_),
    .A2(_07388_),
    .B1(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__and3_1 _35278_ (.A(_07389_),
    .B(_07387_),
    .C(_07388_),
    .X(_07391_));
 sky130_fd_sc_hd__nor4_1 _35279_ (.A(_07375_),
    .B(_07377_),
    .C(_07390_),
    .D(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__buf_1 _35280_ (.A(_20542_),
    .X(_07394_));
 sky130_fd_sc_hd__or3_1 _35281_ (.A(_07394_),
    .B(_19395_),
    .C(_18389_),
    .X(_07395_));
 sky130_fd_sc_hd__o2bb2a_1 _35282_ (.A1_N(_21354_),
    .A2_N(_07395_),
    .B1(_07390_),
    .B2(_07391_),
    .X(_07396_));
 sky130_fd_sc_hd__o211a_1 _35283_ (.A1(net200),
    .A2(_07396_),
    .B1(_05659_),
    .C1(_05662_),
    .X(_07397_));
 sky130_fd_sc_hd__a211oi_1 _35284_ (.A1(_05659_),
    .A2(_05662_),
    .B1(net200),
    .C1(_07396_),
    .Y(_07398_));
 sky130_fd_sc_hd__nor2_1 _35285_ (.A(_07397_),
    .B(_07398_),
    .Y(_07399_));
 sky130_fd_sc_hd__xor2_1 _35286_ (.A(_05663_),
    .B(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__o31a_1 _35287_ (.A1(_18385_),
    .A2(_00708_),
    .A3(_05668_),
    .B1(_05666_),
    .X(_07401_));
 sky130_fd_sc_hd__xor2_1 _35288_ (.A(_07400_),
    .B(_07401_),
    .X(_07402_));
 sky130_fd_sc_hd__a21oi_1 _35289_ (.A1(_05671_),
    .A2(_05724_),
    .B1(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__and3_1 _35290_ (.A(_05671_),
    .B(_05724_),
    .C(_07402_),
    .X(_07405_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35291_ (.A(_00668_),
    .X(_07406_));
 sky130_fd_sc_hd__o221a_1 _35292_ (.A1(_20575_),
    .A2(_07406_),
    .B1(_20548_),
    .B2(_20549_),
    .C1(_20574_),
    .X(_07407_));
 sky130_fd_sc_hd__nor2_1 _35293_ (.A(_05680_),
    .B(_22953_),
    .Y(_07408_));
 sky130_fd_sc_hd__buf_1 _35294_ (.A(_20553_),
    .X(_07409_));
 sky130_fd_sc_hd__nand2_1 _35295_ (.A(_19405_),
    .B(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__a31o_1 _35296_ (.A1(_07410_),
    .A2(_20569_),
    .A3(_21376_),
    .B1(_00668_),
    .X(_07411_));
 sky130_fd_sc_hd__o21a_1 _35297_ (.A1(_07408_),
    .A2(_05683_),
    .B1(_07411_),
    .X(_07412_));
 sky130_fd_sc_hd__o21ai_1 _35298_ (.A1(_05684_),
    .A2(_05685_),
    .B1(_05699_),
    .Y(_07413_));
 sky130_fd_sc_hd__buf_1 _35299_ (.A(\delay_line[19][14] ),
    .X(_07414_));
 sky130_fd_sc_hd__clkbuf_2 _35300_ (.A(_07414_),
    .X(_07416_));
 sky130_fd_sc_hd__or3b_2 _35301_ (.A(_07416_),
    .B(_05692_),
    .C_N(_04045_),
    .X(_07417_));
 sky130_fd_sc_hd__buf_1 _35302_ (.A(net369),
    .X(_07418_));
 sky130_fd_sc_hd__nor2_1 _35303_ (.A(_07418_),
    .B(_07414_),
    .Y(_07419_));
 sky130_fd_sc_hd__and2_1 _35304_ (.A(net369),
    .B(_07414_),
    .X(_07420_));
 sky130_fd_sc_hd__o21bai_4 _35305_ (.A1(_07419_),
    .A2(_07420_),
    .B1_N(_05688_),
    .Y(_07421_));
 sky130_fd_sc_hd__a21o_1 _35306_ (.A1(_07417_),
    .A2(_07421_),
    .B1(_24660_),
    .X(_07422_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35307_ (.A(_24660_),
    .X(_07423_));
 sky130_fd_sc_hd__nand3_1 _35308_ (.A(_07417_),
    .B(_07421_),
    .C(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__clkbuf_2 _35309_ (.A(_05692_),
    .X(_07425_));
 sky130_fd_sc_hd__clkbuf_2 _35310_ (.A(_22946_),
    .X(_07427_));
 sky130_fd_sc_hd__a22o_1 _35311_ (.A1(_07425_),
    .A2(_05691_),
    .B1(_05690_),
    .B2(_07427_),
    .X(_07428_));
 sky130_fd_sc_hd__a21o_1 _35312_ (.A1(_07422_),
    .A2(_07424_),
    .B1(_07428_),
    .X(_07429_));
 sky130_fd_sc_hd__o21a_1 _35313_ (.A1(_19405_),
    .A2(_05680_),
    .B1(_22950_),
    .X(_07430_));
 sky130_fd_sc_hd__clkbuf_2 _35314_ (.A(_22949_),
    .X(_07431_));
 sky130_fd_sc_hd__nor3_2 _35315_ (.A(_20553_),
    .B(_22947_),
    .C(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35316_ (.A(_22947_),
    .X(_07433_));
 sky130_fd_sc_hd__o21a_1 _35317_ (.A1(_07433_),
    .A2(_07431_),
    .B1(_07409_),
    .X(_07434_));
 sky130_fd_sc_hd__nor2_1 _35318_ (.A(_07432_),
    .B(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__xor2_2 _35319_ (.A(_07430_),
    .B(_07435_),
    .X(_07436_));
 sky130_fd_sc_hd__nand3_1 _35320_ (.A(_07428_),
    .B(_07422_),
    .C(_07424_),
    .Y(_07438_));
 sky130_fd_sc_hd__nand3_1 _35321_ (.A(_07429_),
    .B(_07436_),
    .C(_07438_),
    .Y(_07439_));
 sky130_fd_sc_hd__a21o_1 _35322_ (.A1(_07438_),
    .A2(_07429_),
    .B1(_07436_),
    .X(_07440_));
 sky130_fd_sc_hd__nand4_1 _35323_ (.A(_05696_),
    .B(_07413_),
    .C(_07439_),
    .D(_07440_),
    .Y(_07441_));
 sky130_fd_sc_hd__a22o_1 _35324_ (.A1(_05696_),
    .A2(_07413_),
    .B1(_07439_),
    .B2(_07440_),
    .X(_07442_));
 sky130_fd_sc_hd__nand2_1 _35325_ (.A(_07441_),
    .B(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__xor2_1 _35326_ (.A(_07412_),
    .B(_07443_),
    .X(_07444_));
 sky130_fd_sc_hd__a31o_1 _35327_ (.A1(_05703_),
    .A2(_05704_),
    .A3(_04054_),
    .B1(_05679_),
    .X(_07445_));
 sky130_fd_sc_hd__nand3_1 _35328_ (.A(_07444_),
    .B(_07445_),
    .C(_05706_),
    .Y(_07446_));
 sky130_fd_sc_hd__a21o_1 _35329_ (.A1(_05706_),
    .A2(_07445_),
    .B1(_07444_),
    .X(_07447_));
 sky130_fd_sc_hd__nand2_1 _35330_ (.A(_07446_),
    .B(_07447_),
    .Y(_07449_));
 sky130_fd_sc_hd__xor2_1 _35331_ (.A(_07407_),
    .B(_07449_),
    .X(_07450_));
 sky130_fd_sc_hd__and2_1 _35332_ (.A(_05713_),
    .B(_07450_),
    .X(_07451_));
 sky130_fd_sc_hd__nand4_1 _35333_ (.A(_05712_),
    .B(_05713_),
    .C(_20575_),
    .D(_04064_),
    .Y(_07452_));
 sky130_fd_sc_hd__a21oi_1 _35334_ (.A1(_05713_),
    .A2(_07452_),
    .B1(_07450_),
    .Y(_07453_));
 sky130_fd_sc_hd__a21o_1 _35335_ (.A1(_07451_),
    .A2(_07452_),
    .B1(_07453_),
    .X(_07454_));
 sky130_fd_sc_hd__a21oi_1 _35336_ (.A1(_05676_),
    .A2(_05717_),
    .B1(_05721_),
    .Y(_07455_));
 sky130_fd_sc_hd__nor2_1 _35337_ (.A(_07454_),
    .B(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__and2_1 _35338_ (.A(_07455_),
    .B(_07454_),
    .X(_07457_));
 sky130_fd_sc_hd__o22ai_1 _35339_ (.A1(_07403_),
    .A2(_07405_),
    .B1(_07456_),
    .B2(_07457_),
    .Y(_07458_));
 sky130_fd_sc_hd__or4_1 _35340_ (.A(_07403_),
    .B(_07405_),
    .C(_07456_),
    .D(_07457_),
    .X(_07460_));
 sky130_fd_sc_hd__nand2_2 _35341_ (.A(_07458_),
    .B(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__xnor2_4 _35342_ (.A(_07374_),
    .B(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__a21boi_4 _35343_ (.A1(_07320_),
    .A2(_07321_),
    .B1_N(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__nand3b_2 _35344_ (.A_N(_07462_),
    .B(_07320_),
    .C(_07321_),
    .Y(_07464_));
 sky130_fd_sc_hd__o21ai_2 _35345_ (.A1(_05853_),
    .A2(_05858_),
    .B1(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__inv_2 _35346_ (.A(_07463_),
    .Y(_07466_));
 sky130_fd_sc_hd__a221oi_4 _35347_ (.A1(_05851_),
    .A2(_05852_),
    .B1(_07466_),
    .B2(_07464_),
    .C1(_05858_),
    .Y(_07467_));
 sky130_fd_sc_hd__o21bai_2 _35348_ (.A1(_07463_),
    .A2(_07465_),
    .B1_N(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__xor2_4 _35349_ (.A(_07202_),
    .B(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__xnor2_1 _35350_ (.A(_05989_),
    .B(_07469_),
    .Y(_07471_));
 sky130_fd_sc_hd__o21a_1 _35351_ (.A1(_07073_),
    .A2(_07075_),
    .B1(_07471_),
    .X(_07472_));
 sky130_fd_sc_hd__nor3_1 _35352_ (.A(_07073_),
    .B(_07075_),
    .C(_07471_),
    .Y(_07473_));
 sky130_fd_sc_hd__o221a_1 _35353_ (.A1(_05592_),
    .A2(_05992_),
    .B1(_07472_),
    .B2(_07473_),
    .C1(_05994_),
    .X(_07474_));
 sky130_fd_sc_hd__o21a_1 _35354_ (.A1(_05592_),
    .A2(_05992_),
    .B1(_05994_),
    .X(_07475_));
 sky130_fd_sc_hd__or3_1 _35355_ (.A(_07475_),
    .B(_07472_),
    .C(_07473_),
    .X(_07476_));
 sky130_fd_sc_hd__or2b_2 _35356_ (.A(_07474_),
    .B_N(_07476_),
    .X(_07477_));
 sky130_fd_sc_hd__xnor2_4 _35357_ (.A(_06905_),
    .B(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__xnor2_4 _35358_ (.A(_06665_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__inv_2 _35359_ (.A(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__nand3_1 _35360_ (.A(_06660_),
    .B(_06661_),
    .C(_06077_),
    .Y(_07482_));
 sky130_fd_sc_hd__a21oi_1 _35361_ (.A1(_06658_),
    .A2(_07482_),
    .B1(_06662_),
    .Y(_07483_));
 sky130_fd_sc_hd__a211oi_2 _35362_ (.A1(_06659_),
    .A2(_06664_),
    .B1(_07480_),
    .C1(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__buf_4 _35363_ (.A(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__a21o_2 _35364_ (.A1(_05998_),
    .A2(_06001_),
    .B1(_07478_),
    .X(_07486_));
 sky130_fd_sc_hd__inv_2 _35365_ (.A(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__o311a_1 _35366_ (.A1(_06000_),
    .A2(_05405_),
    .A3(_05407_),
    .B1(_07478_),
    .C1(_05998_),
    .X(_07488_));
 sky130_fd_sc_hd__nand2_1 _35367_ (.A(_06661_),
    .B(_06077_),
    .Y(_07489_));
 sky130_fd_sc_hd__or2_1 _35368_ (.A(_06647_),
    .B(_06648_),
    .X(_07490_));
 sky130_fd_sc_hd__a21oi_1 _35369_ (.A1(_06654_),
    .A2(_06655_),
    .B1(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__o211a_1 _35370_ (.A1(_07489_),
    .A2(_07491_),
    .B1(_06662_),
    .C1(_06659_),
    .X(_07493_));
 sky130_fd_sc_hd__o22ai_2 _35371_ (.A1(_07487_),
    .A2(_07488_),
    .B1(_07493_),
    .B2(_07483_),
    .Y(_07494_));
 sky130_fd_sc_hd__o21ai_2 _35372_ (.A1(_06005_),
    .A2(_06009_),
    .B1(_07494_),
    .Y(_07495_));
 sky130_fd_sc_hd__a31o_1 _35373_ (.A1(_05150_),
    .A2(_05151_),
    .A3(_05152_),
    .B1(_05154_),
    .X(_07496_));
 sky130_fd_sc_hd__buf_1 _35374_ (.A(\delay_line[17][14] ),
    .X(_07497_));
 sky130_fd_sc_hd__or2b_2 _35375_ (.A(_07497_),
    .B_N(_03001_),
    .X(_07498_));
 sky130_fd_sc_hd__or3_1 _35376_ (.A(_04551_),
    .B(_04552_),
    .C(_04550_),
    .X(_07499_));
 sky130_fd_sc_hd__o211a_1 _35377_ (.A1(_25264_),
    .A2(_01429_),
    .B1(_07498_),
    .C1(_07499_),
    .X(_07500_));
 sky130_fd_sc_hd__a21oi_1 _35378_ (.A1(_01429_),
    .A2(_25264_),
    .B1(_07498_),
    .Y(_07501_));
 sky130_fd_sc_hd__clkbuf_2 _35379_ (.A(_04574_),
    .X(_07502_));
 sky130_fd_sc_hd__o211a_1 _35380_ (.A1(_07500_),
    .A2(_07501_),
    .B1(_04573_),
    .C1(_07502_),
    .X(_07504_));
 sky130_fd_sc_hd__a211oi_1 _35381_ (.A1(_04573_),
    .A2(_07502_),
    .B1(_07500_),
    .C1(_07501_),
    .Y(_07505_));
 sky130_fd_sc_hd__o21a_1 _35382_ (.A1(_04556_),
    .A2(_04564_),
    .B1(_04565_),
    .X(_07506_));
 sky130_fd_sc_hd__buf_1 _35383_ (.A(\delay_line[17][15] ),
    .X(_07507_));
 sky130_fd_sc_hd__nor2_1 _35384_ (.A(_07497_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__and2_1 _35385_ (.A(_07497_),
    .B(\delay_line[17][15] ),
    .X(_07509_));
 sky130_fd_sc_hd__nor2_1 _35386_ (.A(_01422_),
    .B(_23569_),
    .Y(_07510_));
 sky130_fd_sc_hd__and2_1 _35387_ (.A(_23569_),
    .B(_01422_),
    .X(_07511_));
 sky130_fd_sc_hd__or4_1 _35388_ (.A(_07508_),
    .B(_07509_),
    .C(_07510_),
    .D(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__o22ai_1 _35389_ (.A1(_07508_),
    .A2(_07509_),
    .B1(_07510_),
    .B2(_07511_),
    .Y(_07513_));
 sky130_fd_sc_hd__nand2_1 _35390_ (.A(_07512_),
    .B(_07513_),
    .Y(_07515_));
 sky130_fd_sc_hd__a21oi_4 _35391_ (.A1(_23682_),
    .A2(_01448_),
    .B1(_01447_),
    .Y(_07516_));
 sky130_fd_sc_hd__nor2_1 _35392_ (.A(_07516_),
    .B(_01451_),
    .Y(_07517_));
 sky130_fd_sc_hd__and2_1 _35393_ (.A(_01451_),
    .B(_07516_),
    .X(_07518_));
 sky130_fd_sc_hd__or3_1 _35394_ (.A(_01423_),
    .B(_07517_),
    .C(_07518_),
    .X(_07519_));
 sky130_fd_sc_hd__buf_1 _35395_ (.A(_01423_),
    .X(_07520_));
 sky130_fd_sc_hd__o21ai_1 _35396_ (.A1(_07517_),
    .A2(_07518_),
    .B1(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__nor3_1 _35397_ (.A(_25260_),
    .B(_04560_),
    .C(_04561_),
    .Y(_07522_));
 sky130_fd_sc_hd__a211oi_1 _35398_ (.A1(_07519_),
    .A2(_07521_),
    .B1(_04560_),
    .C1(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__o211ai_2 _35399_ (.A1(_04560_),
    .A2(_07522_),
    .B1(_07519_),
    .C1(_07521_),
    .Y(_07524_));
 sky130_fd_sc_hd__and2b_1 _35400_ (.A_N(_07523_),
    .B(_07524_),
    .X(_07526_));
 sky130_fd_sc_hd__xor2_1 _35401_ (.A(_07515_),
    .B(_07526_),
    .X(_07527_));
 sky130_fd_sc_hd__xor2_1 _35402_ (.A(_07506_),
    .B(_07527_),
    .X(_07528_));
 sky130_fd_sc_hd__nor3_1 _35403_ (.A(_07504_),
    .B(_07505_),
    .C(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__o21a_1 _35404_ (.A1(_07504_),
    .A2(_07505_),
    .B1(_07528_),
    .X(_07530_));
 sky130_fd_sc_hd__or2_1 _35405_ (.A(_07529_),
    .B(_07530_),
    .X(_07531_));
 sky130_fd_sc_hd__o21ba_1 _35406_ (.A1(_04523_),
    .A2(_03043_),
    .B1_N(_04543_),
    .X(_07532_));
 sky130_fd_sc_hd__nor4_1 _35407_ (.A(_19849_),
    .B(_15163_),
    .C(_04532_),
    .D(_04534_),
    .Y(_07533_));
 sky130_fd_sc_hd__or2_1 _35408_ (.A(_07533_),
    .B(_04538_),
    .X(_07534_));
 sky130_fd_sc_hd__nand3b_1 _35409_ (.A_N(_05135_),
    .B(_05138_),
    .C(_05139_),
    .Y(_07535_));
 sky130_fd_sc_hd__nand2_2 _35410_ (.A(_04526_),
    .B(_04525_),
    .Y(_07537_));
 sky130_fd_sc_hd__nor2_1 _35411_ (.A(net362),
    .B(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35412_ (.A(_04526_),
    .X(_07539_));
 sky130_fd_sc_hd__clkbuf_2 _35413_ (.A(_04525_),
    .X(_07540_));
 sky130_fd_sc_hd__nand2_2 _35414_ (.A(net363),
    .B(net362),
    .Y(_07541_));
 sky130_fd_sc_hd__and2b_1 _35415_ (.A_N(net363),
    .B(net362),
    .X(_07542_));
 sky130_fd_sc_hd__a21o_1 _35416_ (.A1(_04525_),
    .A2(_07541_),
    .B1(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__a21oi_1 _35417_ (.A1(_07539_),
    .A2(_07540_),
    .B1(_07543_),
    .Y(_07544_));
 sky130_fd_sc_hd__xnor2_1 _35418_ (.A(_25217_),
    .B(_03035_),
    .Y(_07545_));
 sky130_fd_sc_hd__o21a_1 _35419_ (.A1(_07538_),
    .A2(_07544_),
    .B1(_07545_),
    .X(_07546_));
 sky130_fd_sc_hd__clkbuf_4 _35420_ (.A(_07542_),
    .X(_07548_));
 sky130_fd_sc_hd__a21oi_4 _35421_ (.A1(_07540_),
    .A2(_07541_),
    .B1(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__clkbuf_2 _35422_ (.A(_07545_),
    .X(_07550_));
 sky130_fd_sc_hd__a211oi_4 _35423_ (.A1(_07549_),
    .A2(_07537_),
    .B1(_07538_),
    .C1(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__or4_1 _35424_ (.A(_22130_),
    .B(_07546_),
    .C(_05133_),
    .D(_07551_),
    .X(_07552_));
 sky130_fd_sc_hd__o22ai_2 _35425_ (.A1(_05133_),
    .A2(_00435_),
    .B1(_07546_),
    .B2(_07551_),
    .Y(_07553_));
 sky130_fd_sc_hd__o211a_1 _35426_ (.A1(_04527_),
    .A2(_04532_),
    .B1(_07552_),
    .C1(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__a211oi_2 _35427_ (.A1(_07552_),
    .A2(_07553_),
    .B1(_04527_),
    .C1(_04532_),
    .Y(_07555_));
 sky130_fd_sc_hd__a211o_1 _35428_ (.A1(_05138_),
    .A2(_07535_),
    .B1(_07554_),
    .C1(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__o211ai_2 _35429_ (.A1(_07554_),
    .A2(_07555_),
    .B1(_05138_),
    .C1(_07535_),
    .Y(_07557_));
 sky130_fd_sc_hd__and3_1 _35430_ (.A(_07534_),
    .B(_07556_),
    .C(_07557_),
    .X(_07559_));
 sky130_fd_sc_hd__a21oi_1 _35431_ (.A1(_07556_),
    .A2(_07557_),
    .B1(_07534_),
    .Y(_07560_));
 sky130_fd_sc_hd__nor2_1 _35432_ (.A(_07559_),
    .B(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__o21a_1 _35433_ (.A1(_04542_),
    .A2(_07532_),
    .B1(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__clkbuf_2 _35434_ (.A(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__or3_1 _35435_ (.A(_04542_),
    .B(_07532_),
    .C(_07561_),
    .X(_07564_));
 sky130_fd_sc_hd__inv_2 _35436_ (.A(_07564_),
    .Y(_07565_));
 sky130_fd_sc_hd__nor3_1 _35437_ (.A(_07531_),
    .B(_07563_),
    .C(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__o21a_1 _35438_ (.A1(_07565_),
    .A2(_07562_),
    .B1(_07531_),
    .X(_07567_));
 sky130_fd_sc_hd__or2_1 _35439_ (.A(_07566_),
    .B(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__a21o_1 _35440_ (.A1(_05157_),
    .A2(_07496_),
    .B1(_07568_),
    .X(_07570_));
 sky130_fd_sc_hd__clkbuf_2 _35441_ (.A(_07566_),
    .X(_07571_));
 sky130_fd_sc_hd__o211ai_2 _35442_ (.A1(_07571_),
    .A2(_07567_),
    .B1(_07496_),
    .C1(_05157_),
    .Y(_07572_));
 sky130_fd_sc_hd__o211ai_1 _35443_ (.A1(_03048_),
    .A2(_03053_),
    .B1(_04544_),
    .C1(_04545_),
    .Y(_07573_));
 sky130_fd_sc_hd__o21ai_2 _35444_ (.A1(_04547_),
    .A2(_04587_),
    .B1(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__a21oi_2 _35445_ (.A1(_07570_),
    .A2(_07572_),
    .B1(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__nand3_2 _35446_ (.A(_07574_),
    .B(_07570_),
    .C(_07572_),
    .Y(_07576_));
 sky130_fd_sc_hd__inv_2 _35447_ (.A(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__nor2_2 _35448_ (.A(_07575_),
    .B(_07577_),
    .Y(_07578_));
 sky130_fd_sc_hd__nand2_1 _35449_ (.A(_06664_),
    .B(_06659_),
    .Y(_07579_));
 sky130_fd_sc_hd__a21o_1 _35450_ (.A1(_06659_),
    .A2(_07482_),
    .B1(_06662_),
    .X(_07581_));
 sky130_fd_sc_hd__a21oi_1 _35451_ (.A1(_07579_),
    .A2(_07581_),
    .B1(_07479_),
    .Y(_07582_));
 sky130_fd_sc_hd__a31o_1 _35452_ (.A1(_05155_),
    .A2(_05158_),
    .A3(_06006_),
    .B1(_06005_),
    .X(_07583_));
 sky130_fd_sc_hd__o21bai_4 _35453_ (.A1(_07485_),
    .A2(_07582_),
    .B1_N(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__o211ai_1 _35454_ (.A1(_07485_),
    .A2(_07495_),
    .B1(_07578_),
    .C1(_07584_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand3_4 _35455_ (.A(_07581_),
    .B(_07479_),
    .C(_07579_),
    .Y(_07586_));
 sky130_fd_sc_hd__o211a_1 _35456_ (.A1(_06005_),
    .A2(_06009_),
    .B1(_07586_),
    .C1(_07494_),
    .X(_07587_));
 sky130_fd_sc_hd__a21oi_1 _35457_ (.A1(_07586_),
    .A2(_07494_),
    .B1(_07583_),
    .Y(_07588_));
 sky130_fd_sc_hd__o22ai_1 _35458_ (.A1(_07575_),
    .A2(_07577_),
    .B1(_07587_),
    .B2(_07588_),
    .Y(_07589_));
 sky130_fd_sc_hd__nand3_2 _35459_ (.A(_06076_),
    .B(_07585_),
    .C(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__o21ai_1 _35460_ (.A1(_07587_),
    .A2(_07588_),
    .B1(_07578_),
    .Y(_07592_));
 sky130_fd_sc_hd__o221ai_4 _35461_ (.A1(_07575_),
    .A2(_07577_),
    .B1(_07485_),
    .B2(_07495_),
    .C1(_07584_),
    .Y(_07593_));
 sky130_fd_sc_hd__nand3b_1 _35462_ (.A_N(_06076_),
    .B(_07592_),
    .C(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__nand3_1 _35463_ (.A(_03608_),
    .B(_04451_),
    .C(_04591_),
    .Y(_07595_));
 sky130_fd_sc_hd__and2_1 _35464_ (.A(_04594_),
    .B(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35465_ (.A(_25240_),
    .X(_07597_));
 sky130_fd_sc_hd__o21bai_1 _35466_ (.A1(_18812_),
    .A2(_18813_),
    .B1_N(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__or3b_1 _35467_ (.A(_18812_),
    .B(_18813_),
    .C_N(_07597_),
    .X(_07599_));
 sky130_fd_sc_hd__o21ai_2 _35468_ (.A1(_25238_),
    .A2(_18725_),
    .B1(_18726_),
    .Y(_07600_));
 sky130_fd_sc_hd__a21oi_1 _35469_ (.A1(_07598_),
    .A2(_07599_),
    .B1(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__and3_1 _35470_ (.A(_07600_),
    .B(_07598_),
    .C(_07599_),
    .X(_07603_));
 sky130_fd_sc_hd__o211ai_1 _35471_ (.A1(_07601_),
    .A2(_07603_),
    .B1(_04578_),
    .C1(_04583_),
    .Y(_07604_));
 sky130_fd_sc_hd__inv_2 _35472_ (.A(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__a211oi_2 _35473_ (.A1(_04578_),
    .A2(_04583_),
    .B1(_07601_),
    .C1(_07603_),
    .Y(_07606_));
 sky130_fd_sc_hd__or3_2 _35474_ (.A(_07605_),
    .B(_06028_),
    .C(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__o21ai_2 _35475_ (.A1(_07606_),
    .A2(_07605_),
    .B1(_06028_),
    .Y(_07608_));
 sky130_fd_sc_hd__a211oi_4 _35476_ (.A1(_07607_),
    .A2(_07608_),
    .B1(_04571_),
    .C1(_04586_),
    .Y(_07609_));
 sky130_fd_sc_hd__o211a_2 _35477_ (.A1(_04571_),
    .A2(_04586_),
    .B1(_07607_),
    .C1(_07608_),
    .X(_07610_));
 sky130_fd_sc_hd__o221ai_4 _35478_ (.A1(_04477_),
    .A2(_06032_),
    .B1(_07609_),
    .B2(_07610_),
    .C1(_06033_),
    .Y(_07611_));
 sky130_fd_sc_hd__a211o_1 _35479_ (.A1(_06033_),
    .A2(_06036_),
    .B1(_07609_),
    .C1(_07610_),
    .X(_07612_));
 sky130_fd_sc_hd__nand2_1 _35480_ (.A(_07611_),
    .B(_07612_),
    .Y(_07614_));
 sky130_fd_sc_hd__or2_2 _35481_ (.A(_06038_),
    .B(_06043_),
    .X(_07615_));
 sky130_fd_sc_hd__xnor2_1 _35482_ (.A(_07614_),
    .B(_07615_),
    .Y(_07616_));
 sky130_fd_sc_hd__o21a_1 _35483_ (.A1(_04592_),
    .A2(_07596_),
    .B1(_07616_),
    .X(_07617_));
 sky130_fd_sc_hd__a211oi_1 _35484_ (.A1(_04594_),
    .A2(_07595_),
    .B1(_07616_),
    .C1(_04592_),
    .Y(_07618_));
 sky130_fd_sc_hd__nor2_1 _35485_ (.A(_07617_),
    .B(_07618_),
    .Y(_07619_));
 sky130_fd_sc_hd__o31a_1 _35486_ (.A1(_06044_),
    .A2(_06042_),
    .A3(_06043_),
    .B1(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__o21a_1 _35487_ (.A1(_07617_),
    .A2(_07618_),
    .B1(net95),
    .X(_07621_));
 sky130_fd_sc_hd__nor2_1 _35488_ (.A(_07620_),
    .B(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__nand3_1 _35489_ (.A(_07590_),
    .B(_07594_),
    .C(_07622_),
    .Y(_07623_));
 sky130_fd_sc_hd__o2bb2ai_1 _35490_ (.A1_N(_07590_),
    .A2_N(_07594_),
    .B1(_07620_),
    .B2(_07621_),
    .Y(_07625_));
 sky130_fd_sc_hd__o2111ai_1 _35491_ (.A1(_06075_),
    .A2(_06053_),
    .B1(_06023_),
    .C1(_07623_),
    .D1(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__o21a_1 _35492_ (.A1(_06075_),
    .A2(_06053_),
    .B1(_06023_),
    .X(_07627_));
 sky130_fd_sc_hd__a21o_1 _35493_ (.A1(_07623_),
    .A2(_07625_),
    .B1(_07627_),
    .X(_07628_));
 sky130_fd_sc_hd__a22o_1 _35494_ (.A1(_06050_),
    .A2(_06074_),
    .B1(_07626_),
    .B2(_07628_),
    .X(_07629_));
 sky130_fd_sc_hd__nand4_1 _35495_ (.A(_06050_),
    .B(_06074_),
    .C(_07626_),
    .D(_07628_),
    .Y(_07630_));
 sky130_fd_sc_hd__o21a_1 _35496_ (.A1(_06062_),
    .A2(_06057_),
    .B1(_06058_),
    .X(_07631_));
 sky130_fd_sc_hd__a21o_1 _35497_ (.A1(_07629_),
    .A2(_07630_),
    .B1(_07631_),
    .X(_07632_));
 sky130_fd_sc_hd__inv_2 _35498_ (.A(_07631_),
    .Y(_07633_));
 sky130_fd_sc_hd__nand2_1 _35499_ (.A(_07629_),
    .B(_07630_),
    .Y(_07634_));
 sky130_fd_sc_hd__or2_1 _35500_ (.A(_07633_),
    .B(_07634_),
    .X(_07636_));
 sky130_fd_sc_hd__nand2_1 _35501_ (.A(_06069_),
    .B(_06066_),
    .Y(_07637_));
 sky130_fd_sc_hd__o2bb2ai_2 _35502_ (.A1_N(_06067_),
    .A2_N(_07637_),
    .B1(_07633_),
    .B2(_07634_),
    .Y(_07638_));
 sky130_fd_sc_hd__a22oi_1 _35503_ (.A1(_06067_),
    .A2(_07637_),
    .B1(_07632_),
    .B2(_07636_),
    .Y(_07639_));
 sky130_fd_sc_hd__a31o_2 _35504_ (.A1(_07632_),
    .A2(_07636_),
    .A3(_07638_),
    .B1(_07639_),
    .X(_00009_));
 sky130_fd_sc_hd__and2_2 _35505_ (.A(_07632_),
    .B(_07638_),
    .X(_07640_));
 sky130_fd_sc_hd__inv_2 _35506_ (.A(_07578_),
    .Y(_07641_));
 sky130_fd_sc_hd__o22ai_1 _35507_ (.A1(_07485_),
    .A2(_07495_),
    .B1(_07641_),
    .B2(_07588_),
    .Y(_07642_));
 sky130_fd_sc_hd__a31oi_4 _35508_ (.A1(_06611_),
    .A2(_06613_),
    .A3(_06617_),
    .B1(_06626_),
    .Y(_07643_));
 sky130_fd_sc_hd__o21ai_2 _35509_ (.A1(_06715_),
    .A2(_06768_),
    .B1(_06713_),
    .Y(_07644_));
 sky130_fd_sc_hd__o211ai_2 _35510_ (.A1(_06567_),
    .A2(_05086_),
    .B1(_06572_),
    .C1(_06596_),
    .Y(_07646_));
 sky130_fd_sc_hd__o2111ai_4 _35511_ (.A1(_05081_),
    .A2(_05084_),
    .B1(_05089_),
    .C1(_06581_),
    .D1(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__o21ai_1 _35512_ (.A1(_06566_),
    .A2(_06573_),
    .B1(_05093_),
    .Y(_07648_));
 sky130_fd_sc_hd__nand2_2 _35513_ (.A(_06581_),
    .B(_07648_),
    .Y(_07649_));
 sky130_fd_sc_hd__a31oi_4 _35514_ (.A1(_05017_),
    .A2(_06544_),
    .A3(_05053_),
    .B1(_06543_),
    .Y(_07650_));
 sky130_fd_sc_hd__o21a_1 _35515_ (.A1(_06391_),
    .A2(_06389_),
    .B1(_06393_),
    .X(_07651_));
 sky130_fd_sc_hd__a22oi_4 _35516_ (.A1(_06394_),
    .A2(_07651_),
    .B1(_06388_),
    .B2(_06476_),
    .Y(_07652_));
 sky130_fd_sc_hd__inv_2 _35517_ (.A(_06465_),
    .Y(_07653_));
 sky130_fd_sc_hd__a21o_1 _35518_ (.A1(_22509_),
    .A2(_06428_),
    .B1(_21869_),
    .X(_07654_));
 sky130_fd_sc_hd__nand3_1 _35519_ (.A(_23953_),
    .B(_01739_),
    .C(_06428_),
    .Y(_07655_));
 sky130_fd_sc_hd__and4_1 _35520_ (.A(_06406_),
    .B(_06411_),
    .C(_07654_),
    .D(_07655_),
    .X(_07657_));
 sky130_fd_sc_hd__inv_2 _35521_ (.A(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__a22o_2 _35522_ (.A1(_06406_),
    .A2(_06411_),
    .B1(_07654_),
    .B2(_07655_),
    .X(_07659_));
 sky130_fd_sc_hd__and3_1 _35523_ (.A(_07658_),
    .B(_06434_),
    .C(_07659_),
    .X(_07660_));
 sky130_fd_sc_hd__a21oi_1 _35524_ (.A1(_07659_),
    .A2(_07658_),
    .B1(_06434_),
    .Y(_07661_));
 sky130_fd_sc_hd__and4b_1 _35525_ (.A_N(_17916_),
    .B(_03369_),
    .C(_04650_),
    .D(_06419_),
    .X(_07662_));
 sky130_fd_sc_hd__a21oi_1 _35526_ (.A1(_03368_),
    .A2(_04649_),
    .B1(_06398_),
    .Y(_07663_));
 sky130_fd_sc_hd__nor2_1 _35527_ (.A(net423),
    .B(\delay_line[8][15] ),
    .Y(_07664_));
 sky130_fd_sc_hd__and2_1 _35528_ (.A(net423),
    .B(\delay_line[8][15] ),
    .X(_07665_));
 sky130_fd_sc_hd__o21bai_2 _35529_ (.A1(_07664_),
    .A2(_07665_),
    .B1_N(_03367_),
    .Y(_07666_));
 sky130_fd_sc_hd__nand2_1 _35530_ (.A(_04649_),
    .B(_06416_),
    .Y(_07668_));
 sky130_fd_sc_hd__nand3b_1 _35531_ (.A_N(_07664_),
    .B(_07668_),
    .C(_03368_),
    .Y(_07669_));
 sky130_fd_sc_hd__o211ai_2 _35532_ (.A1(_06400_),
    .A2(_07663_),
    .B1(_07666_),
    .C1(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__inv_2 _35533_ (.A(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__a221oi_2 _35534_ (.A1(_03369_),
    .A2(_06412_),
    .B1(_07666_),
    .B2(_07669_),
    .C1(_07663_),
    .Y(_07672_));
 sky130_fd_sc_hd__o21a_1 _35535_ (.A1(_07671_),
    .A2(_07672_),
    .B1(_03354_),
    .X(_07673_));
 sky130_fd_sc_hd__nor3_1 _35536_ (.A(_07672_),
    .B(_03354_),
    .C(_07671_),
    .Y(_07674_));
 sky130_fd_sc_hd__clkbuf_2 _35537_ (.A(_06412_),
    .X(_07675_));
 sky130_fd_sc_hd__xor2_2 _35538_ (.A(_22439_),
    .B(_06416_),
    .X(_07676_));
 sky130_fd_sc_hd__a311o_1 _35539_ (.A1(_06419_),
    .A2(_22543_),
    .A3(_07675_),
    .B1(_07676_),
    .C1(_06417_),
    .X(_07677_));
 sky130_fd_sc_hd__and3_1 _35540_ (.A(_06419_),
    .B(_22543_),
    .C(_07675_),
    .X(_07679_));
 sky130_fd_sc_hd__o21ai_1 _35541_ (.A1(_06417_),
    .A2(_07679_),
    .B1(_07676_),
    .Y(_07680_));
 sky130_fd_sc_hd__o211ai_1 _35542_ (.A1(_07673_),
    .A2(_07674_),
    .B1(_07677_),
    .C1(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__a211o_1 _35543_ (.A1(_07677_),
    .A2(_07680_),
    .B1(_07673_),
    .C1(_07674_),
    .X(_07682_));
 sky130_fd_sc_hd__o211a_1 _35544_ (.A1(_06423_),
    .A2(_07662_),
    .B1(_07681_),
    .C1(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__a211oi_1 _35545_ (.A1(_07681_),
    .A2(_07682_),
    .B1(_06423_),
    .C1(_07662_),
    .Y(_07684_));
 sky130_fd_sc_hd__or4_1 _35546_ (.A(_07660_),
    .B(_07661_),
    .C(_07683_),
    .D(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__o22ai_2 _35547_ (.A1(_07660_),
    .A2(_07661_),
    .B1(_07683_),
    .B2(_07684_),
    .Y(_07686_));
 sky130_fd_sc_hd__o21ba_2 _35548_ (.A1(_06446_),
    .A2(_06455_),
    .B1_N(_06454_),
    .X(_07687_));
 sky130_fd_sc_hd__nand3b_1 _35549_ (.A_N(_04840_),
    .B(_06344_),
    .C(_06345_),
    .Y(_07688_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35550_ (.A(_03265_),
    .X(_07690_));
 sky130_fd_sc_hd__clkbuf_2 _35551_ (.A(_06335_),
    .X(_07691_));
 sky130_fd_sc_hd__or3b_4 _35552_ (.A(_07690_),
    .B(_07691_),
    .C_N(_06445_),
    .X(_07692_));
 sky130_fd_sc_hd__and3_1 _35553_ (.A(_06332_),
    .B(_06333_),
    .C(_04838_),
    .X(_07693_));
 sky130_fd_sc_hd__buf_1 _35554_ (.A(\delay_line[9][15] ),
    .X(_07694_));
 sky130_fd_sc_hd__clkbuf_2 _35555_ (.A(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__nand2_2 _35556_ (.A(_04614_),
    .B(_04828_),
    .Y(_07696_));
 sky130_fd_sc_hd__nor2_1 _35557_ (.A(_04828_),
    .B(_07694_),
    .Y(_07697_));
 sky130_fd_sc_hd__and2_1 _35558_ (.A(_04828_),
    .B(_07694_),
    .X(_07698_));
 sky130_fd_sc_hd__a2bb2o_1 _35559_ (.A1_N(_07697_),
    .A2_N(_07698_),
    .B1(_06445_),
    .B2(_06335_),
    .X(_07699_));
 sky130_fd_sc_hd__o211ai_4 _35560_ (.A1(_07695_),
    .A2(_07696_),
    .B1(_25341_),
    .C1(_07699_),
    .Y(_07701_));
 sky130_fd_sc_hd__or2_2 _35561_ (.A(_07694_),
    .B(_07696_),
    .X(_07702_));
 sky130_fd_sc_hd__clkbuf_2 _35562_ (.A(_25341_),
    .X(_07703_));
 sky130_fd_sc_hd__a21o_1 _35563_ (.A1(_07699_),
    .A2(_07702_),
    .B1(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__o211a_1 _35564_ (.A1(_07693_),
    .A2(_06339_),
    .B1(_07701_),
    .C1(_07704_),
    .X(_07705_));
 sky130_fd_sc_hd__a221oi_2 _35565_ (.A1(_06334_),
    .A2(_06336_),
    .B1(_07704_),
    .B2(_07701_),
    .C1(_07693_),
    .Y(_07706_));
 sky130_fd_sc_hd__a211oi_2 _35566_ (.A1(_06453_),
    .A2(_07692_),
    .B1(_07705_),
    .C1(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__o211a_1 _35567_ (.A1(_07705_),
    .A2(_07706_),
    .B1(_06453_),
    .C1(_07692_),
    .X(_07708_));
 sky130_fd_sc_hd__a211o_1 _35568_ (.A1(_07688_),
    .A2(_06349_),
    .B1(_07707_),
    .C1(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__o211ai_2 _35569_ (.A1(_07707_),
    .A2(_07708_),
    .B1(_07688_),
    .C1(_06349_),
    .Y(_07710_));
 sky130_fd_sc_hd__and3b_1 _35570_ (.A_N(_07687_),
    .B(_07709_),
    .C(_07710_),
    .X(_07712_));
 sky130_fd_sc_hd__inv_2 _35571_ (.A(_07710_),
    .Y(_07713_));
 sky130_fd_sc_hd__o21ai_2 _35572_ (.A1(_07687_),
    .A2(_07713_),
    .B1(_07709_),
    .Y(_07714_));
 sky130_fd_sc_hd__nor2_1 _35573_ (.A(_06460_),
    .B(_06463_),
    .Y(_07715_));
 sky130_fd_sc_hd__o221ai_4 _35574_ (.A1(_07687_),
    .A2(_07712_),
    .B1(_07713_),
    .B2(_07714_),
    .C1(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__nand2_1 _35575_ (.A(_07709_),
    .B(_07710_),
    .Y(_07717_));
 sky130_fd_sc_hd__a211o_1 _35576_ (.A1(_07687_),
    .A2(_07717_),
    .B1(_07712_),
    .C1(_07715_),
    .X(_07718_));
 sky130_fd_sc_hd__nand4_2 _35577_ (.A(_07685_),
    .B(_07686_),
    .C(_07716_),
    .D(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__a22o_1 _35578_ (.A1(_07685_),
    .A2(_07686_),
    .B1(_07716_),
    .B2(_07718_),
    .X(_07720_));
 sky130_fd_sc_hd__o211a_2 _35579_ (.A1(_06373_),
    .A2(_06377_),
    .B1(_07719_),
    .C1(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__a221oi_2 _35580_ (.A1(_06374_),
    .A2(_06372_),
    .B1(_07719_),
    .B2(_07720_),
    .C1(_06377_),
    .Y(_07723_));
 sky130_fd_sc_hd__nor2_1 _35581_ (.A(_07721_),
    .B(_07723_),
    .Y(_07724_));
 sky130_fd_sc_hd__o21a_4 _35582_ (.A1(_07653_),
    .A2(_06467_),
    .B1(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__nor3_1 _35583_ (.A(_07653_),
    .B(_06467_),
    .C(_07724_),
    .Y(_07726_));
 sky130_fd_sc_hd__o21ai_2 _35584_ (.A1(_06318_),
    .A2(_06311_),
    .B1(_06383_),
    .Y(_07727_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35585_ (.A(_04796_),
    .X(_07728_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35586_ (.A(\delay_line[12][15] ),
    .X(_07729_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35587_ (.A(_00121_),
    .X(_07730_));
 sky130_fd_sc_hd__a21o_1 _35588_ (.A1(_07728_),
    .A2(_07729_),
    .B1(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__nand3_2 _35589_ (.A(_07730_),
    .B(_07728_),
    .C(_07729_),
    .Y(_07732_));
 sky130_fd_sc_hd__nand3_2 _35590_ (.A(_07731_),
    .B(_06299_),
    .C(_07732_),
    .Y(_07734_));
 sky130_fd_sc_hd__a21o_1 _35591_ (.A1(_07732_),
    .A2(_07731_),
    .B1(_06299_),
    .X(_07735_));
 sky130_fd_sc_hd__o211a_1 _35592_ (.A1(_06298_),
    .A2(_06303_),
    .B1(_07734_),
    .C1(_07735_),
    .X(_07736_));
 sky130_fd_sc_hd__clkbuf_2 _35593_ (.A(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__a211oi_4 _35594_ (.A1(_07734_),
    .A2(_07735_),
    .B1(_06298_),
    .C1(_06303_),
    .Y(_07738_));
 sky130_fd_sc_hd__a311oi_4 _35595_ (.A1(_23898_),
    .A2(_06204_),
    .A3(_06203_),
    .B1(_07737_),
    .C1(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__o2111a_1 _35596_ (.A1(_07737_),
    .A2(_07738_),
    .B1(_23898_),
    .C1(_06204_),
    .D1(_06203_),
    .X(_07740_));
 sky130_fd_sc_hd__a21oi_2 _35597_ (.A1(_06285_),
    .A2(_06290_),
    .B1(_06212_),
    .Y(_07741_));
 sky130_fd_sc_hd__inv_2 _35598_ (.A(_06308_),
    .Y(_07742_));
 sky130_fd_sc_hd__a31oi_4 _35599_ (.A1(_06212_),
    .A2(_06285_),
    .A3(_06290_),
    .B1(_07742_),
    .Y(_07743_));
 sky130_fd_sc_hd__nand2_1 _35600_ (.A(_06258_),
    .B(_04729_),
    .Y(_07745_));
 sky130_fd_sc_hd__or2b_1 _35601_ (.A(_25433_),
    .B_N(\delay_line[11][13] ),
    .X(_07746_));
 sky130_fd_sc_hd__nand2_1 _35602_ (.A(_04710_),
    .B(_06235_),
    .Y(_07747_));
 sky130_fd_sc_hd__clkbuf_2 _35603_ (.A(_07747_),
    .X(_07748_));
 sky130_fd_sc_hd__or2b_1 _35604_ (.A(_01555_),
    .B_N(net409),
    .X(_07749_));
 sky130_fd_sc_hd__nand2b_1 _35605_ (.A_N(\delay_line[11][14] ),
    .B(_06233_),
    .Y(_07750_));
 sky130_fd_sc_hd__nand2_1 _35606_ (.A(_07749_),
    .B(_07750_),
    .Y(_07751_));
 sky130_fd_sc_hd__a21oi_1 _35607_ (.A1(_07746_),
    .A2(_07748_),
    .B1(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__and3_1 _35608_ (.A(_07746_),
    .B(_07751_),
    .C(_07747_),
    .X(_07753_));
 sky130_fd_sc_hd__or2_2 _35609_ (.A(_07752_),
    .B(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__nor2_1 _35610_ (.A(_06239_),
    .B(_04715_),
    .Y(_07756_));
 sky130_fd_sc_hd__nor2_1 _35611_ (.A(_06234_),
    .B(_06237_),
    .Y(_07757_));
 sky130_fd_sc_hd__a31o_1 _35612_ (.A1(_04706_),
    .A2(_04713_),
    .A3(_06235_),
    .B1(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__a21oi_4 _35613_ (.A1(_04717_),
    .A2(_07756_),
    .B1(_07758_),
    .Y(_07759_));
 sky130_fd_sc_hd__nor2_1 _35614_ (.A(_07754_),
    .B(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__nor2_1 _35615_ (.A(_07752_),
    .B(_07753_),
    .Y(_07761_));
 sky130_fd_sc_hd__nand2_1 _35616_ (.A(_04718_),
    .B(_06248_),
    .Y(_07762_));
 sky130_fd_sc_hd__o21bai_2 _35617_ (.A1(_07762_),
    .A2(_06246_),
    .B1_N(_07758_),
    .Y(_07763_));
 sky130_fd_sc_hd__nor2_1 _35618_ (.A(_07761_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__inv_2 _35619_ (.A(net433),
    .Y(_07765_));
 sky130_fd_sc_hd__clkbuf_2 _35620_ (.A(_07765_),
    .X(_07767_));
 sky130_fd_sc_hd__or3b_2 _35621_ (.A(_07767_),
    .B(_04694_),
    .C_N(_04695_),
    .X(_07768_));
 sky130_fd_sc_hd__or2_1 _35622_ (.A(_03160_),
    .B(_07765_),
    .X(_07769_));
 sky130_fd_sc_hd__nand3b_2 _35623_ (.A_N(_03169_),
    .B(_06225_),
    .C(_06219_),
    .Y(_07770_));
 sky130_fd_sc_hd__xnor2_2 _35624_ (.A(\delay_line[4][11] ),
    .B(\delay_line[4][13] ),
    .Y(_07771_));
 sky130_fd_sc_hd__and3_1 _35625_ (.A(_07769_),
    .B(_07770_),
    .C(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__a21oi_2 _35626_ (.A1(_07769_),
    .A2(_07770_),
    .B1(_07771_),
    .Y(_07773_));
 sky130_fd_sc_hd__nor2_2 _35627_ (.A(_07772_),
    .B(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__a21oi_2 _35628_ (.A1(_06244_),
    .A2(_07768_),
    .B1(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__and3_1 _35629_ (.A(_06244_),
    .B(_07774_),
    .C(_07768_),
    .X(_07776_));
 sky130_fd_sc_hd__o22ai_2 _35630_ (.A1(_07760_),
    .A2(_07764_),
    .B1(_07775_),
    .B2(_07776_),
    .Y(_07778_));
 sky130_fd_sc_hd__nand2_1 _35631_ (.A(_06243_),
    .B(_06253_),
    .Y(_07779_));
 sky130_fd_sc_hd__and3_1 _35632_ (.A(net433),
    .B(_03162_),
    .C(_04695_),
    .X(_07780_));
 sky130_fd_sc_hd__o22ai_4 _35633_ (.A1(_07772_),
    .A2(_07773_),
    .B1(_07780_),
    .B2(_06255_),
    .Y(_07781_));
 sky130_fd_sc_hd__nand3_2 _35634_ (.A(_06244_),
    .B(_07774_),
    .C(_07768_),
    .Y(_07782_));
 sky130_fd_sc_hd__nor2_1 _35635_ (.A(_07760_),
    .B(_07764_),
    .Y(_07783_));
 sky130_fd_sc_hd__nand3_1 _35636_ (.A(_07781_),
    .B(_07782_),
    .C(_07783_),
    .Y(_07784_));
 sky130_fd_sc_hd__o211a_1 _35637_ (.A1(_06255_),
    .A2(_06256_),
    .B1(_07779_),
    .C1(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__buf_2 _35638_ (.A(\delay_line[0][15] ),
    .X(_07786_));
 sky130_fd_sc_hd__a21boi_1 _35639_ (.A1(_06243_),
    .A2(_07786_),
    .B1_N(_06252_),
    .Y(_07787_));
 sky130_fd_sc_hd__a21oi_1 _35640_ (.A1(_07778_),
    .A2(_07784_),
    .B1(_07787_),
    .Y(_07789_));
 sky130_fd_sc_hd__a21oi_1 _35641_ (.A1(_07778_),
    .A2(_07785_),
    .B1(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__a21oi_2 _35642_ (.A1(_06265_),
    .A2(_07745_),
    .B1(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__buf_2 _35643_ (.A(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__clkinvlp_2 _35644_ (.A(_06252_),
    .Y(_07793_));
 sky130_fd_sc_hd__nand2_1 _35645_ (.A(_06229_),
    .B(_06244_),
    .Y(_07794_));
 sky130_fd_sc_hd__nand2_1 _35646_ (.A(_06250_),
    .B(_06251_),
    .Y(_07795_));
 sky130_fd_sc_hd__inv_2 _35647_ (.A(_06253_),
    .Y(_07796_));
 sky130_fd_sc_hd__a21oi_1 _35648_ (.A1(_07794_),
    .A2(_07795_),
    .B1(_07796_),
    .Y(_07797_));
 sky130_fd_sc_hd__a21oi_2 _35649_ (.A1(_07781_),
    .A2(_07782_),
    .B1(_07783_),
    .Y(_07798_));
 sky130_fd_sc_hd__nand2_1 _35650_ (.A(_07783_),
    .B(_07782_),
    .Y(_07800_));
 sky130_fd_sc_hd__nor2_1 _35651_ (.A(_07775_),
    .B(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__o22ai_1 _35652_ (.A1(_07793_),
    .A2(_07797_),
    .B1(_07798_),
    .B2(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__o211ai_2 _35653_ (.A1(_07775_),
    .A2(_07800_),
    .B1(_07787_),
    .C1(_07778_),
    .Y(_07803_));
 sky130_fd_sc_hd__nand3_2 _35654_ (.A(_06265_),
    .B(_07802_),
    .C(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__buf_1 _35655_ (.A(\delay_line[13][15] ),
    .X(_07805_));
 sky130_fd_sc_hd__and3_1 _35656_ (.A(_04751_),
    .B(_07805_),
    .C(_01630_),
    .X(_07806_));
 sky130_fd_sc_hd__buf_1 _35657_ (.A(_07805_),
    .X(_07807_));
 sky130_fd_sc_hd__nor2_1 _35658_ (.A(_03191_),
    .B(_07805_),
    .Y(_07808_));
 sky130_fd_sc_hd__inv_2 _35659_ (.A(\delay_line[13][15] ),
    .Y(_07809_));
 sky130_fd_sc_hd__nor2_1 _35660_ (.A(_04751_),
    .B(_07809_),
    .Y(_07811_));
 sky130_fd_sc_hd__o2bb2a_1 _35661_ (.A1_N(_01630_),
    .A2_N(_07807_),
    .B1(_07808_),
    .B2(_07811_),
    .X(_07812_));
 sky130_fd_sc_hd__nor2_1 _35662_ (.A(_07806_),
    .B(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__o21ai_2 _35663_ (.A1(_07804_),
    .A2(_06268_),
    .B1(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__a21oi_1 _35664_ (.A1(_06273_),
    .A2(_06259_),
    .B1(_07804_),
    .Y(_07815_));
 sky130_fd_sc_hd__o22ai_4 _35665_ (.A1(_07806_),
    .A2(_07812_),
    .B1(_07815_),
    .B2(_07791_),
    .Y(_07816_));
 sky130_fd_sc_hd__a21oi_1 _35666_ (.A1(_06270_),
    .A2(_06274_),
    .B1(_06275_),
    .Y(_07817_));
 sky130_fd_sc_hd__o21ai_2 _35667_ (.A1(_06289_),
    .A2(_07817_),
    .B1(_06277_),
    .Y(_07818_));
 sky130_fd_sc_hd__o211ai_2 _35668_ (.A1(_07792_),
    .A2(_07814_),
    .B1(_07816_),
    .C1(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__o21ai_2 _35669_ (.A1(_07792_),
    .A2(_07814_),
    .B1(_07816_),
    .Y(_07820_));
 sky130_fd_sc_hd__a21boi_2 _35670_ (.A1(_06269_),
    .A2(_06294_),
    .B1_N(_06276_),
    .Y(_07822_));
 sky130_fd_sc_hd__nand2_1 _35671_ (.A(_07820_),
    .B(_07822_),
    .Y(_07823_));
 sky130_fd_sc_hd__xnor2_1 _35672_ (.A(_00096_),
    .B(\delay_line[13][14] ),
    .Y(_07824_));
 sky130_fd_sc_hd__and4b_1 _35673_ (.A_N(_00096_),
    .B(_06278_),
    .C(_06280_),
    .D(_04772_),
    .X(_07825_));
 sky130_fd_sc_hd__a21oi_2 _35674_ (.A1(_06286_),
    .A2(_07824_),
    .B1(_07825_),
    .Y(_07826_));
 sky130_fd_sc_hd__and3_1 _35675_ (.A(_01537_),
    .B(_04771_),
    .C(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__a21oi_2 _35676_ (.A1(_01537_),
    .A2(_04775_),
    .B1(_07826_),
    .Y(_07828_));
 sky130_fd_sc_hd__nor2_1 _35677_ (.A(_07827_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__nand3_1 _35678_ (.A(_07819_),
    .B(_07823_),
    .C(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__nor2_2 _35679_ (.A(_07822_),
    .B(_07820_),
    .Y(_07831_));
 sky130_fd_sc_hd__a21o_1 _35680_ (.A1(_06259_),
    .A2(_06273_),
    .B1(_07804_),
    .X(_07833_));
 sky130_fd_sc_hd__nand3b_1 _35681_ (.A_N(_07792_),
    .B(_07813_),
    .C(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__a21oi_2 _35682_ (.A1(_07834_),
    .A2(_07816_),
    .B1(_07818_),
    .Y(_07835_));
 sky130_fd_sc_hd__o22ai_4 _35683_ (.A1(_07827_),
    .A2(_07828_),
    .B1(_07831_),
    .B2(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__o211ai_4 _35684_ (.A1(_07741_),
    .A2(_07743_),
    .B1(_07830_),
    .C1(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__o21ai_1 _35685_ (.A1(_07831_),
    .A2(_07835_),
    .B1(_07829_),
    .Y(_07838_));
 sky130_fd_sc_hd__a21oi_1 _35686_ (.A1(_06291_),
    .A2(_06308_),
    .B1(_07741_),
    .Y(_07839_));
 sky130_fd_sc_hd__o211ai_1 _35687_ (.A1(_07827_),
    .A2(_07828_),
    .B1(_07819_),
    .C1(_07823_),
    .Y(_07840_));
 sky130_fd_sc_hd__nand3_1 _35688_ (.A(_07838_),
    .B(_07839_),
    .C(_07840_),
    .Y(_07841_));
 sky130_fd_sc_hd__buf_6 _35689_ (.A(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__o211ai_2 _35690_ (.A1(_07739_),
    .A2(_07740_),
    .B1(_07837_),
    .C1(_07842_),
    .Y(_07844_));
 sky130_fd_sc_hd__nor3_2 _35691_ (.A(_07738_),
    .B(_06206_),
    .C(_07736_),
    .Y(_07845_));
 sky130_fd_sc_hd__o21a_1 _35692_ (.A1(_07737_),
    .A2(_07738_),
    .B1(_06206_),
    .X(_07846_));
 sky130_fd_sc_hd__o2bb2ai_2 _35693_ (.A1_N(_07837_),
    .A2_N(_07842_),
    .B1(_07845_),
    .B2(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__nand3_2 _35694_ (.A(_07727_),
    .B(_07844_),
    .C(_07847_),
    .Y(_07848_));
 sky130_fd_sc_hd__nand2_1 _35695_ (.A(_06320_),
    .B(_06319_),
    .Y(_07849_));
 sky130_fd_sc_hd__and3_1 _35696_ (.A(_07819_),
    .B(_07823_),
    .C(_07829_),
    .X(_07850_));
 sky130_fd_sc_hd__o21ai_2 _35697_ (.A1(_07741_),
    .A2(_07743_),
    .B1(_07836_),
    .Y(_07851_));
 sky130_fd_sc_hd__o221ai_2 _35698_ (.A1(_07845_),
    .A2(_07846_),
    .B1(_07850_),
    .B2(_07851_),
    .C1(_07842_),
    .Y(_07852_));
 sky130_fd_sc_hd__o2bb2ai_1 _35699_ (.A1_N(_07837_),
    .A2_N(_07841_),
    .B1(_07739_),
    .B2(_07740_),
    .Y(_07853_));
 sky130_fd_sc_hd__nand4_2 _35700_ (.A(_06383_),
    .B(_07849_),
    .C(_07852_),
    .D(_07853_),
    .Y(_07855_));
 sky130_fd_sc_hd__buf_4 _35701_ (.A(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__o2bb2a_1 _35702_ (.A1_N(_06352_),
    .A2_N(_06367_),
    .B1(_06371_),
    .B2(_06351_),
    .X(_07857_));
 sky130_fd_sc_hd__or2_2 _35703_ (.A(_06208_),
    .B(_06210_),
    .X(_07858_));
 sky130_fd_sc_hd__or2_1 _35704_ (.A(_04842_),
    .B(_25375_),
    .X(_07859_));
 sky130_fd_sc_hd__nand2_1 _35705_ (.A(_04842_),
    .B(_25370_),
    .Y(_07860_));
 sky130_fd_sc_hd__buf_1 _35706_ (.A(\delay_line[10][13] ),
    .X(_07861_));
 sky130_fd_sc_hd__nand3_1 _35707_ (.A(_07859_),
    .B(_07860_),
    .C(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__clkbuf_2 _35708_ (.A(_07861_),
    .X(_07863_));
 sky130_fd_sc_hd__a21o_1 _35709_ (.A1(_07859_),
    .A2(_07860_),
    .B1(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__nand3b_2 _35710_ (.A_N(_06344_),
    .B(_07862_),
    .C(_07864_),
    .Y(_07866_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35711_ (.A(_03281_),
    .X(_07867_));
 sky130_fd_sc_hd__a32o_1 _35712_ (.A1(_07867_),
    .A2(_06342_),
    .A3(_06343_),
    .B1(_07862_),
    .B2(_07864_),
    .X(_07868_));
 sky130_fd_sc_hd__buf_1 _35713_ (.A(_06330_),
    .X(_07869_));
 sky130_fd_sc_hd__clkbuf_2 _35714_ (.A(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__nor2_1 _35715_ (.A(_22456_),
    .B(_06331_),
    .Y(_07871_));
 sky130_fd_sc_hd__nand2_1 _35716_ (.A(_06331_),
    .B(_22456_),
    .Y(_07872_));
 sky130_fd_sc_hd__or4b_2 _35717_ (.A(_06341_),
    .B(_23762_),
    .C(_07871_),
    .D_N(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__or2_1 _35718_ (.A(_21801_),
    .B(_06331_),
    .X(_07874_));
 sky130_fd_sc_hd__a22o_1 _35719_ (.A1(_01694_),
    .A2(_04842_),
    .B1(_07874_),
    .B2(_07872_),
    .X(_07875_));
 sky130_fd_sc_hd__or4bb_4 _35720_ (.A(_04611_),
    .B(_07870_),
    .C_N(_07873_),
    .D_N(_07875_),
    .X(_07877_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35721_ (.A(_07870_),
    .X(_07878_));
 sky130_fd_sc_hd__a2bb2o_1 _35722_ (.A1_N(_04611_),
    .A2_N(_07878_),
    .B1(_07873_),
    .B2(_07875_),
    .X(_07879_));
 sky130_fd_sc_hd__nand4_2 _35723_ (.A(_07866_),
    .B(_07868_),
    .C(_07877_),
    .D(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__a22o_1 _35724_ (.A1(_07866_),
    .A2(_07868_),
    .B1(_07877_),
    .B2(_07879_),
    .X(_07881_));
 sky130_fd_sc_hd__nand2_2 _35725_ (.A(_07880_),
    .B(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__o21a_1 _35726_ (.A1(_06353_),
    .A2(_01529_),
    .B1(_06355_),
    .X(_07883_));
 sky130_fd_sc_hd__nand2_1 _35727_ (.A(_01529_),
    .B(_06353_),
    .Y(_07884_));
 sky130_fd_sc_hd__o2bb2a_1 _35728_ (.A1_N(_07883_),
    .A2_N(_07884_),
    .B1(_06355_),
    .B2(_06202_),
    .X(_07885_));
 sky130_fd_sc_hd__a21boi_2 _35729_ (.A1(_06201_),
    .A2(_06204_),
    .B1_N(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__nor2_1 _35730_ (.A(net399),
    .B(_06200_),
    .Y(_07888_));
 sky130_fd_sc_hd__a221o_1 _35731_ (.A1(_07728_),
    .A2(_07888_),
    .B1(_06199_),
    .B2(_06202_),
    .C1(_07885_),
    .X(_07889_));
 sky130_fd_sc_hd__and3b_1 _35732_ (.A_N(_07886_),
    .B(_07889_),
    .C(_06356_),
    .X(_07890_));
 sky130_fd_sc_hd__buf_1 _35733_ (.A(_06202_),
    .X(_07891_));
 sky130_fd_sc_hd__a221oi_1 _35734_ (.A1(_07728_),
    .A2(_07888_),
    .B1(_06199_),
    .B2(_07891_),
    .C1(_07885_),
    .Y(_07892_));
 sky130_fd_sc_hd__o32a_1 _35735_ (.A1(_06365_),
    .A2(_06354_),
    .A3(_06357_),
    .B1(_07886_),
    .B2(_07892_),
    .X(_07893_));
 sky130_fd_sc_hd__a211o_1 _35736_ (.A1(_06361_),
    .A2(_06368_),
    .B1(_07890_),
    .C1(_07893_),
    .X(_07894_));
 sky130_fd_sc_hd__o211ai_1 _35737_ (.A1(_07890_),
    .A2(_07893_),
    .B1(_06361_),
    .C1(_06368_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand2_2 _35738_ (.A(_07894_),
    .B(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__xor2_4 _35739_ (.A(_07882_),
    .B(_07896_),
    .X(_07897_));
 sky130_fd_sc_hd__xnor2_2 _35740_ (.A(_07858_),
    .B(_07897_),
    .Y(_07899_));
 sky130_fd_sc_hd__nor2_4 _35741_ (.A(_07857_),
    .B(_07899_),
    .Y(_07900_));
 sky130_fd_sc_hd__and2_2 _35742_ (.A(_07899_),
    .B(_07857_),
    .X(_07901_));
 sky130_fd_sc_hd__nor2_2 _35743_ (.A(_07900_),
    .B(_07901_),
    .Y(_07902_));
 sky130_fd_sc_hd__and3_2 _35744_ (.A(_07848_),
    .B(_07856_),
    .C(_07902_),
    .X(_07903_));
 sky130_fd_sc_hd__inv_2 _35745_ (.A(_06379_),
    .Y(_07904_));
 sky130_fd_sc_hd__a31oi_4 _35746_ (.A1(_06323_),
    .A2(_06324_),
    .A3(_06325_),
    .B1(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__o2bb2ai_4 _35747_ (.A1_N(_07848_),
    .A2_N(_07856_),
    .B1(_07900_),
    .B2(_07901_),
    .Y(_07906_));
 sky130_fd_sc_hd__o21ai_4 _35748_ (.A1(_06391_),
    .A2(_07905_),
    .B1(_07906_),
    .Y(_07907_));
 sky130_fd_sc_hd__a21oi_1 _35749_ (.A1(_06327_),
    .A2(_06380_),
    .B1(_06390_),
    .Y(_07908_));
 sky130_fd_sc_hd__nor2_1 _35750_ (.A(_07845_),
    .B(_07846_),
    .Y(_07910_));
 sky130_fd_sc_hd__and3_2 _35751_ (.A(_07837_),
    .B(_07842_),
    .C(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__nand2_2 _35752_ (.A(_07727_),
    .B(_07847_),
    .Y(_07912_));
 sky130_fd_sc_hd__o221ai_4 _35753_ (.A1(_07900_),
    .A2(_07901_),
    .B1(_07911_),
    .B2(_07912_),
    .C1(_07855_),
    .Y(_07913_));
 sky130_fd_sc_hd__inv_2 _35754_ (.A(_07857_),
    .Y(_07914_));
 sky130_fd_sc_hd__nor2_1 _35755_ (.A(_07914_),
    .B(_07899_),
    .Y(_07915_));
 sky130_fd_sc_hd__and2_1 _35756_ (.A(_07914_),
    .B(_07899_),
    .X(_07916_));
 sky130_fd_sc_hd__o2bb2ai_2 _35757_ (.A1_N(_07848_),
    .A2_N(_07856_),
    .B1(_07915_),
    .B2(_07916_),
    .Y(_07917_));
 sky130_fd_sc_hd__nand3_2 _35758_ (.A(_07908_),
    .B(_07913_),
    .C(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__o221ai_4 _35759_ (.A1(_07725_),
    .A2(net100),
    .B1(_07903_),
    .B2(_07907_),
    .C1(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__o211ai_4 _35760_ (.A1(_07911_),
    .A2(_07912_),
    .B1(_07856_),
    .C1(_07902_),
    .Y(_07921_));
 sky130_fd_sc_hd__o211ai_4 _35761_ (.A1(_06391_),
    .A2(_07905_),
    .B1(_07921_),
    .C1(_07906_),
    .Y(_07922_));
 sky130_fd_sc_hd__buf_4 _35762_ (.A(_07918_),
    .X(_07923_));
 sky130_fd_sc_hd__nor4_1 _35763_ (.A(_07653_),
    .B(_06467_),
    .C(_07721_),
    .D(_07723_),
    .Y(_07924_));
 sky130_fd_sc_hd__o22a_1 _35764_ (.A1(_07653_),
    .A2(_06467_),
    .B1(_07721_),
    .B2(_07723_),
    .X(_07925_));
 sky130_fd_sc_hd__o2bb2ai_4 _35765_ (.A1_N(_07922_),
    .A2_N(_07923_),
    .B1(net106),
    .B2(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__nand3_1 _35766_ (.A(_07652_),
    .B(_07919_),
    .C(_07926_),
    .Y(_07927_));
 sky130_fd_sc_hd__buf_6 _35767_ (.A(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__o22ai_4 _35768_ (.A1(_06382_),
    .A2(_06488_),
    .B1(_06475_),
    .B2(_06484_),
    .Y(_07929_));
 sky130_fd_sc_hd__o2bb2ai_2 _35769_ (.A1_N(_07922_),
    .A2_N(_07923_),
    .B1(_07725_),
    .B2(_07726_),
    .Y(_07930_));
 sky130_fd_sc_hd__nor2_2 _35770_ (.A(_07725_),
    .B(net100),
    .Y(_07932_));
 sky130_fd_sc_hd__o211ai_2 _35771_ (.A1(_07903_),
    .A2(_07907_),
    .B1(_07923_),
    .C1(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__nand3_4 _35772_ (.A(_07929_),
    .B(_07930_),
    .C(_07933_),
    .Y(_07934_));
 sky130_fd_sc_hd__nand2_4 _35773_ (.A(_06121_),
    .B(_06189_),
    .Y(_07935_));
 sky130_fd_sc_hd__a21o_1 _35774_ (.A1(_06085_),
    .A2(_04671_),
    .B1(_06112_),
    .X(_07936_));
 sky130_fd_sc_hd__nand2_1 _35775_ (.A(_07936_),
    .B(_06116_),
    .Y(_07937_));
 sky130_fd_sc_hd__a31o_1 _35776_ (.A1(_06441_),
    .A2(_06440_),
    .A3(_06426_),
    .B1(_06424_),
    .X(_07938_));
 sky130_fd_sc_hd__a21oi_2 _35777_ (.A1(_04662_),
    .A2(_06439_),
    .B1(_06437_),
    .Y(_07939_));
 sky130_fd_sc_hd__or2b_2 _35778_ (.A(\delay_line[7][8] ),
    .B_N(\delay_line[6][15] ),
    .X(_07940_));
 sky130_fd_sc_hd__or2b_1 _35779_ (.A(_06088_),
    .B_N(\delay_line[7][8] ),
    .X(_07941_));
 sky130_fd_sc_hd__o21a_1 _35780_ (.A1(_04973_),
    .A2(_25296_),
    .B1(net425),
    .X(_07943_));
 sky130_fd_sc_hd__a211o_1 _35781_ (.A1(_07940_),
    .A2(_07941_),
    .B1(_06101_),
    .C1(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__o211ai_4 _35782_ (.A1(_06101_),
    .A2(_07943_),
    .B1(_07940_),
    .C1(_07941_),
    .Y(_07945_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35783_ (.A(_06088_),
    .X(_07946_));
 sky130_fd_sc_hd__clkbuf_2 _35784_ (.A(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__and4b_1 _35785_ (.A_N(_01912_),
    .B(_07944_),
    .C(_07945_),
    .D(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__a21boi_1 _35786_ (.A1(_07944_),
    .A2(_07945_),
    .B1_N(_06089_),
    .Y(_07949_));
 sky130_fd_sc_hd__or2_1 _35787_ (.A(\delay_line[7][11] ),
    .B(\delay_line[7][12] ),
    .X(_07950_));
 sky130_fd_sc_hd__nand2_1 _35788_ (.A(\delay_line[7][11] ),
    .B(\delay_line[7][12] ),
    .Y(_07951_));
 sky130_fd_sc_hd__a21o_1 _35789_ (.A1(_07950_),
    .A2(_07951_),
    .B1(_01909_),
    .X(_07952_));
 sky130_fd_sc_hd__nand3_1 _35790_ (.A(_07950_),
    .B(_07951_),
    .C(_01909_),
    .Y(_07954_));
 sky130_fd_sc_hd__and4bb_1 _35791_ (.A_N(_07948_),
    .B_N(_07949_),
    .C(_07952_),
    .D(_07954_),
    .X(_07955_));
 sky130_fd_sc_hd__a2bb2oi_1 _35792_ (.A1_N(_07948_),
    .A2_N(_07949_),
    .B1(_07952_),
    .B2(_07954_),
    .Y(_07956_));
 sky130_fd_sc_hd__nor2_1 _35793_ (.A(_07955_),
    .B(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__xor2_1 _35794_ (.A(_07939_),
    .B(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__xnor2_1 _35795_ (.A(_06109_),
    .B(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__nor2_1 _35796_ (.A(_07938_),
    .B(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__nand2_2 _35797_ (.A(_07959_),
    .B(_07938_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand2b_1 _35798_ (.A_N(_07960_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__o31a_1 _35799_ (.A1(_06098_),
    .A2(_06099_),
    .A3(_06104_),
    .B1(_06107_),
    .X(_07963_));
 sky130_fd_sc_hd__o21ba_2 _35800_ (.A1(_04988_),
    .A2(_06110_),
    .B1_N(_07963_),
    .X(_07965_));
 sky130_fd_sc_hd__xnor2_1 _35801_ (.A(_07962_),
    .B(_07965_),
    .Y(_07966_));
 sky130_fd_sc_hd__xnor2_1 _35802_ (.A(_07937_),
    .B(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__nand2_1 _35803_ (.A(_06134_),
    .B(_06136_),
    .Y(_07968_));
 sky130_fd_sc_hd__and3_1 _35804_ (.A(_06162_),
    .B(_04956_),
    .C(_06163_),
    .X(_07969_));
 sky130_fd_sc_hd__and4_1 _35805_ (.A(_04940_),
    .B(_06126_),
    .C(_06127_),
    .D(_04941_),
    .X(_07970_));
 sky130_fd_sc_hd__nor2_1 _35806_ (.A(net435),
    .B(net438),
    .Y(_07971_));
 sky130_fd_sc_hd__and2_1 _35807_ (.A(\delay_line[3][14] ),
    .B(net438),
    .X(_07972_));
 sky130_fd_sc_hd__nor2_1 _35808_ (.A(_07971_),
    .B(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__or2_1 _35809_ (.A(_06146_),
    .B(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__o21ai_1 _35810_ (.A1(_24040_),
    .A2(_06147_),
    .B1(_07973_),
    .Y(_07976_));
 sky130_fd_sc_hd__and2b_1 _35811_ (.A_N(\delay_line[3][13] ),
    .B(net438),
    .X(_07977_));
 sky130_fd_sc_hd__and3_1 _35812_ (.A(_07974_),
    .B(_07976_),
    .C(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__a21oi_1 _35813_ (.A1(_07974_),
    .A2(_07976_),
    .B1(_07977_),
    .Y(_07979_));
 sky130_fd_sc_hd__nor2_1 _35814_ (.A(_07978_),
    .B(_07979_),
    .Y(_07980_));
 sky130_fd_sc_hd__xnor2_1 _35815_ (.A(_06153_),
    .B(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__nor2_1 _35816_ (.A(_07970_),
    .B(_07981_),
    .Y(_07982_));
 sky130_fd_sc_hd__a21boi_2 _35817_ (.A1(_06129_),
    .A2(_06133_),
    .B1_N(_07981_),
    .Y(_07983_));
 sky130_fd_sc_hd__a21oi_1 _35818_ (.A1(_07982_),
    .A2(_06133_),
    .B1(_07983_),
    .Y(_07984_));
 sky130_fd_sc_hd__nor3_1 _35819_ (.A(_07969_),
    .B(_06166_),
    .C(_07984_),
    .Y(_07985_));
 sky130_fd_sc_hd__o21a_1 _35820_ (.A1(_07969_),
    .A2(_06166_),
    .B1(_07984_),
    .X(_07987_));
 sky130_fd_sc_hd__nor2_1 _35821_ (.A(_07985_),
    .B(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__xor2_1 _35822_ (.A(_07968_),
    .B(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__o21ba_1 _35823_ (.A1(_06177_),
    .A2(_06178_),
    .B1_N(_06181_),
    .X(_07990_));
 sky130_fd_sc_hd__a21oi_2 _35824_ (.A1(_06154_),
    .A2(_06156_),
    .B1(_01884_),
    .Y(_07991_));
 sky130_fd_sc_hd__and3_1 _35825_ (.A(_06156_),
    .B(_01884_),
    .C(_06154_),
    .X(_07992_));
 sky130_fd_sc_hd__nor3_1 _35826_ (.A(_07991_),
    .B(_07992_),
    .C(_06163_),
    .Y(_07993_));
 sky130_fd_sc_hd__o21a_1 _35827_ (.A1(_07991_),
    .A2(_07992_),
    .B1(_06163_),
    .X(_07994_));
 sky130_fd_sc_hd__nor2_1 _35828_ (.A(net250),
    .B(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__buf_1 _35829_ (.A(\delay_line[3][15] ),
    .X(_07996_));
 sky130_fd_sc_hd__nor2_1 _35830_ (.A(_01863_),
    .B(_07996_),
    .Y(_07998_));
 sky130_fd_sc_hd__and2_1 _35831_ (.A(_01863_),
    .B(_07996_),
    .X(_07999_));
 sky130_fd_sc_hd__o21ai_2 _35832_ (.A1(_07998_),
    .A2(_07999_),
    .B1(_06157_),
    .Y(_08000_));
 sky130_fd_sc_hd__or3_1 _35833_ (.A(_06157_),
    .B(_07998_),
    .C(_07999_),
    .X(_08001_));
 sky130_fd_sc_hd__and3_1 _35834_ (.A(_07995_),
    .B(_08000_),
    .C(_08001_),
    .X(_08002_));
 sky130_fd_sc_hd__o2bb2a_1 _35835_ (.A1_N(_08001_),
    .A2_N(_08000_),
    .B1(net250),
    .B2(_07994_),
    .X(_08003_));
 sky130_fd_sc_hd__or2_1 _35836_ (.A(_08002_),
    .B(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__nand3b_1 _35837_ (.A_N(_04979_),
    .B(_06094_),
    .C(_06096_),
    .Y(_08005_));
 sky130_fd_sc_hd__o21a_1 _35838_ (.A1(_01920_),
    .A2(_06168_),
    .B1(_04978_),
    .X(_08006_));
 sky130_fd_sc_hd__nor3_1 _35839_ (.A(_01920_),
    .B(_06168_),
    .C(_06097_),
    .Y(_08007_));
 sky130_fd_sc_hd__a211o_1 _35840_ (.A1(_06096_),
    .A2(_08005_),
    .B1(_08006_),
    .C1(_08007_),
    .X(_08009_));
 sky130_fd_sc_hd__clkbuf_2 _35841_ (.A(_06168_),
    .X(_08010_));
 sky130_fd_sc_hd__o21a_1 _35842_ (.A1(_03424_),
    .A2(_08010_),
    .B1(_04927_),
    .X(_08011_));
 sky130_fd_sc_hd__o211ai_2 _35843_ (.A1(_08006_),
    .A2(_08007_),
    .B1(_06096_),
    .C1(_08005_),
    .Y(_08012_));
 sky130_fd_sc_hd__and3_1 _35844_ (.A(_08009_),
    .B(_08011_),
    .C(_08012_),
    .X(_08013_));
 sky130_fd_sc_hd__a21oi_1 _35845_ (.A1(_08012_),
    .A2(_08009_),
    .B1(_08011_),
    .Y(_08014_));
 sky130_fd_sc_hd__nor2_1 _35846_ (.A(_08013_),
    .B(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__o21a_1 _35847_ (.A1(_06175_),
    .A2(_06176_),
    .B1(_06174_),
    .X(_08016_));
 sky130_fd_sc_hd__xor2_1 _35848_ (.A(_08015_),
    .B(_08016_),
    .X(_08017_));
 sky130_fd_sc_hd__or2_1 _35849_ (.A(_08004_),
    .B(_08017_),
    .X(_08018_));
 sky130_fd_sc_hd__nand2_1 _35850_ (.A(_08004_),
    .B(_08017_),
    .Y(_08020_));
 sky130_fd_sc_hd__nand2_1 _35851_ (.A(_08018_),
    .B(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__xor2_1 _35852_ (.A(_07990_),
    .B(_08021_),
    .X(_08022_));
 sky130_fd_sc_hd__xor2_1 _35853_ (.A(_07989_),
    .B(_08022_),
    .X(_08023_));
 sky130_fd_sc_hd__and2_1 _35854_ (.A(_07967_),
    .B(_08023_),
    .X(_08024_));
 sky130_fd_sc_hd__nor2_1 _35855_ (.A(_07967_),
    .B(_08023_),
    .Y(_08025_));
 sky130_fd_sc_hd__a21boi_2 _35856_ (.A1(_06396_),
    .A2(_06471_),
    .B1_N(_06472_),
    .Y(_08026_));
 sky130_fd_sc_hd__o21a_1 _35857_ (.A1(_08024_),
    .A2(_08025_),
    .B1(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__or3_2 _35858_ (.A(_08026_),
    .B(_08024_),
    .C(_08025_),
    .X(_08028_));
 sky130_fd_sc_hd__or2b_4 _35859_ (.A(_08027_),
    .B_N(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__xnor2_4 _35860_ (.A(_07935_),
    .B(_08029_),
    .Y(_08031_));
 sky130_fd_sc_hd__a21oi_1 _35861_ (.A1(_07928_),
    .A2(_07934_),
    .B1(_08031_),
    .Y(_08032_));
 sky130_fd_sc_hd__and3_1 _35862_ (.A(_07928_),
    .B(_07934_),
    .C(_08031_),
    .X(_08033_));
 sky130_fd_sc_hd__a21oi_2 _35863_ (.A1(_06489_),
    .A2(_06486_),
    .B1(_06487_),
    .Y(_08034_));
 sky130_fd_sc_hd__a21oi_1 _35864_ (.A1(_06195_),
    .A2(_06494_),
    .B1(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__o21ai_2 _35865_ (.A1(_08032_),
    .A2(_08033_),
    .B1(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__a31oi_2 _35866_ (.A1(_06486_),
    .A2(_06487_),
    .A3(_06489_),
    .B1(_06196_),
    .Y(_08037_));
 sky130_fd_sc_hd__nand2_1 _35867_ (.A(_07927_),
    .B(_07934_),
    .Y(_08038_));
 sky130_fd_sc_hd__xor2_4 _35868_ (.A(_07935_),
    .B(_08029_),
    .X(_08039_));
 sky130_fd_sc_hd__nand2_4 _35869_ (.A(_08038_),
    .B(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__nand3_4 _35870_ (.A(_07928_),
    .B(_07934_),
    .C(_08031_),
    .Y(_08042_));
 sky130_fd_sc_hd__o211ai_4 _35871_ (.A1(_08034_),
    .A2(_08037_),
    .B1(_08040_),
    .C1(_08042_),
    .Y(_08043_));
 sky130_fd_sc_hd__inv_2 _35872_ (.A(_06191_),
    .Y(_08044_));
 sky130_fd_sc_hd__o21a_1 _35873_ (.A1(_06506_),
    .A2(_06537_),
    .B1(_06536_),
    .X(_08045_));
 sky130_fd_sc_hd__clkbuf_2 _35874_ (.A(_05024_),
    .X(_08046_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _35875_ (.A(_05025_),
    .X(_08047_));
 sky130_fd_sc_hd__a211o_1 _35876_ (.A1(_08046_),
    .A2(_08047_),
    .B1(_03082_),
    .C1(_01493_),
    .X(_08048_));
 sky130_fd_sc_hd__a22o_1 _35877_ (.A1(_06514_),
    .A2(_06515_),
    .B1(_01841_),
    .B2(_05027_),
    .X(_08049_));
 sky130_fd_sc_hd__a21oi_1 _35878_ (.A1(_06509_),
    .A2(_08049_),
    .B1(_06516_),
    .Y(_08050_));
 sky130_fd_sc_hd__and4_1 _35879_ (.A(_06511_),
    .B(_06512_),
    .C(_03488_),
    .D(net439),
    .X(_08051_));
 sky130_fd_sc_hd__a31oi_1 _35880_ (.A1(_06511_),
    .A2(_06512_),
    .A3(_03488_),
    .B1(net439),
    .Y(_08053_));
 sky130_fd_sc_hd__a21o_1 _35881_ (.A1(net446),
    .A2(net445),
    .B1(_05027_),
    .X(_08054_));
 sky130_fd_sc_hd__or3_1 _35882_ (.A(_05025_),
    .B(_05024_),
    .C(_06510_),
    .X(_08055_));
 sky130_fd_sc_hd__and3_1 _35883_ (.A(_08054_),
    .B(_08055_),
    .C(_03086_),
    .X(_08056_));
 sky130_fd_sc_hd__a21oi_1 _35884_ (.A1(_08054_),
    .A2(_08055_),
    .B1(_03086_),
    .Y(_08057_));
 sky130_fd_sc_hd__nor4_1 _35885_ (.A(_08051_),
    .B(_08053_),
    .C(_08056_),
    .D(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__o22ai_1 _35886_ (.A1(_08051_),
    .A2(_08053_),
    .B1(_08056_),
    .B2(_08057_),
    .Y(_08059_));
 sky130_fd_sc_hd__inv_2 _35887_ (.A(_08059_),
    .Y(_08060_));
 sky130_fd_sc_hd__nor3_1 _35888_ (.A(_08050_),
    .B(net199),
    .C(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__o21ai_1 _35889_ (.A1(net199),
    .A2(_08060_),
    .B1(_08050_),
    .Y(_08062_));
 sky130_fd_sc_hd__inv_2 _35890_ (.A(_08062_),
    .Y(_08064_));
 sky130_fd_sc_hd__or3_1 _35891_ (.A(_08048_),
    .B(_08061_),
    .C(_08064_),
    .X(_08065_));
 sky130_fd_sc_hd__o21ai_1 _35892_ (.A1(_08061_),
    .A2(_08064_),
    .B1(_08048_),
    .Y(_08066_));
 sky130_fd_sc_hd__o211a_1 _35893_ (.A1(_06141_),
    .A2(_06145_),
    .B1(_08065_),
    .C1(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__a211oi_1 _35894_ (.A1(_08065_),
    .A2(_08066_),
    .B1(_06141_),
    .C1(_06145_),
    .Y(_08068_));
 sky130_fd_sc_hd__nor2_1 _35895_ (.A(_08067_),
    .B(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__nor3_1 _35896_ (.A(_06521_),
    .B(net168),
    .C(_08069_),
    .Y(_08070_));
 sky130_fd_sc_hd__o21a_1 _35897_ (.A1(_06521_),
    .A2(net168),
    .B1(_08069_),
    .X(_08071_));
 sky130_fd_sc_hd__nor2_1 _35898_ (.A(_08070_),
    .B(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__a21bo_1 _35899_ (.A1(_06182_),
    .A2(_06186_),
    .B1_N(_08072_),
    .X(_08073_));
 sky130_fd_sc_hd__o211ai_2 _35900_ (.A1(_08070_),
    .A2(_08071_),
    .B1(_06182_),
    .C1(_06186_),
    .Y(_08075_));
 sky130_fd_sc_hd__nand2_1 _35901_ (.A(_08073_),
    .B(_08075_),
    .Y(_08076_));
 sky130_fd_sc_hd__a21bo_1 _35902_ (.A1(_06527_),
    .A2(_06529_),
    .B1_N(_06526_),
    .X(_08077_));
 sky130_fd_sc_hd__xnor2_1 _35903_ (.A(_08076_),
    .B(_08077_),
    .Y(_08078_));
 sky130_fd_sc_hd__xor2_1 _35904_ (.A(_08045_),
    .B(_08078_),
    .X(_08079_));
 sky130_fd_sc_hd__a31o_1 _35905_ (.A1(_08044_),
    .A2(_06550_),
    .A3(_08079_),
    .B1(_06540_),
    .X(_08080_));
 sky130_fd_sc_hd__a21oi_1 _35906_ (.A1(_08044_),
    .A2(_06550_),
    .B1(_08079_),
    .Y(_08081_));
 sky130_fd_sc_hd__buf_1 _35907_ (.A(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__and3_1 _35908_ (.A(_08044_),
    .B(_06550_),
    .C(_08079_),
    .X(_08083_));
 sky130_fd_sc_hd__or2_1 _35909_ (.A(_08081_),
    .B(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__a2bb2o_1 _35910_ (.A1_N(_08080_),
    .A2_N(_08082_),
    .B1(_06540_),
    .B2(_08084_),
    .X(_08086_));
 sky130_fd_sc_hd__a21oi_1 _35911_ (.A1(_08036_),
    .A2(_08043_),
    .B1(_08086_),
    .Y(_08087_));
 sky130_fd_sc_hd__nand3_2 _35912_ (.A(_08086_),
    .B(_08036_),
    .C(_08043_),
    .Y(_08088_));
 sky130_fd_sc_hd__o211ai_1 _35913_ (.A1(_06547_),
    .A2(_06498_),
    .B1(_06560_),
    .C1(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__o21ai_1 _35914_ (.A1(_06547_),
    .A2(_06498_),
    .B1(_06560_),
    .Y(_08090_));
 sky130_fd_sc_hd__o2bb2a_2 _35915_ (.A1_N(_06540_),
    .A2_N(_08084_),
    .B1(_08080_),
    .B2(_08082_),
    .X(_08091_));
 sky130_fd_sc_hd__nand3_1 _35916_ (.A(_08036_),
    .B(_08043_),
    .C(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__nor2_1 _35917_ (.A(_08082_),
    .B(_08080_),
    .Y(_08093_));
 sky130_fd_sc_hd__o32a_1 _35918_ (.A1(_06504_),
    .A2(_06538_),
    .A3(_06539_),
    .B1(_08082_),
    .B2(_08083_),
    .X(_08094_));
 sky130_fd_sc_hd__o2bb2ai_2 _35919_ (.A1_N(_06195_),
    .A2_N(_06494_),
    .B1(_06482_),
    .B2(_06477_),
    .Y(_08095_));
 sky130_fd_sc_hd__a21oi_4 _35920_ (.A1(_08040_),
    .A2(_08042_),
    .B1(_08095_),
    .Y(_08097_));
 sky130_fd_sc_hd__o211a_1 _35921_ (.A1(_08034_),
    .A2(_08037_),
    .B1(_08040_),
    .C1(_08042_),
    .X(_08098_));
 sky130_fd_sc_hd__o22ai_1 _35922_ (.A1(_08093_),
    .A2(_08094_),
    .B1(_08097_),
    .B2(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand3_1 _35923_ (.A(_08090_),
    .B(_08092_),
    .C(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__o21ai_1 _35924_ (.A1(_08087_),
    .A2(_08089_),
    .B1(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__o21ai_2 _35925_ (.A1(_08097_),
    .A2(_08098_),
    .B1(_08091_),
    .Y(_08102_));
 sky130_fd_sc_hd__a2bb2oi_2 _35926_ (.A1_N(_06499_),
    .A2_N(_06553_),
    .B1(_06554_),
    .B2(_06556_),
    .Y(_08103_));
 sky130_fd_sc_hd__a21oi_2 _35927_ (.A1(_08088_),
    .A2(_08102_),
    .B1(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__a31o_1 _35928_ (.A1(_08102_),
    .A2(_08103_),
    .A3(_08088_),
    .B1(_07650_),
    .X(_08105_));
 sky130_fd_sc_hd__o2bb2ai_1 _35929_ (.A1_N(_07650_),
    .A2_N(_08101_),
    .B1(_08104_),
    .B2(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__o22a_1 _35930_ (.A1(_06571_),
    .A2(_06570_),
    .B1(_06578_),
    .B2(_06575_),
    .X(_08108_));
 sky130_fd_sc_hd__nand2_1 _35931_ (.A(_08106_),
    .B(_08108_),
    .Y(_08109_));
 sky130_fd_sc_hd__o22ai_2 _35932_ (.A1(_06571_),
    .A2(_06570_),
    .B1(_06578_),
    .B2(_06575_),
    .Y(_08110_));
 sky130_fd_sc_hd__nand2_1 _35933_ (.A(_08101_),
    .B(_07650_),
    .Y(_08111_));
 sky130_fd_sc_hd__a31oi_2 _35934_ (.A1(_08102_),
    .A2(_08103_),
    .A3(_08088_),
    .B1(_07650_),
    .Y(_08112_));
 sky130_fd_sc_hd__nand2_1 _35935_ (.A(_08112_),
    .B(_08100_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand3_2 _35936_ (.A(_08110_),
    .B(_08111_),
    .C(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand2_2 _35937_ (.A(_08109_),
    .B(_08114_),
    .Y(_08115_));
 sky130_fd_sc_hd__o211a_1 _35938_ (.A1(_06593_),
    .A2(_07647_),
    .B1(_07649_),
    .C1(_08115_),
    .X(_08116_));
 sky130_fd_sc_hd__nor2_1 _35939_ (.A(_05081_),
    .B(_05084_),
    .Y(_08117_));
 sky130_fd_sc_hd__nor2_1 _35940_ (.A(_08117_),
    .B(_06589_),
    .Y(_08119_));
 sky130_fd_sc_hd__nand4_2 _35941_ (.A(_06597_),
    .B(_03544_),
    .C(_08119_),
    .D(_03559_),
    .Y(_08120_));
 sky130_fd_sc_hd__a21oi_2 _35942_ (.A1(_07649_),
    .A2(_08120_),
    .B1(_08115_),
    .Y(_08121_));
 sky130_fd_sc_hd__a21oi_4 _35943_ (.A1(_06750_),
    .A2(_06767_),
    .B1(_06749_),
    .Y(_08122_));
 sky130_fd_sc_hd__o21ai_4 _35944_ (.A1(_08116_),
    .A2(_08121_),
    .B1(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__and3_1 _35945_ (.A(_06576_),
    .B(_06577_),
    .C(_06580_),
    .X(_08124_));
 sky130_fd_sc_hd__o22a_1 _35946_ (.A1(_05088_),
    .A2(_06584_),
    .B1(_06566_),
    .B2(_06573_),
    .X(_08125_));
 sky130_fd_sc_hd__o221ai_4 _35947_ (.A1(_08124_),
    .A2(_08125_),
    .B1(_06582_),
    .B2(_05094_),
    .C1(_08115_),
    .Y(_08126_));
 sky130_fd_sc_hd__o21ai_4 _35948_ (.A1(_06593_),
    .A2(_07647_),
    .B1(_07649_),
    .Y(_08127_));
 sky130_fd_sc_hd__inv_2 _35949_ (.A(_08115_),
    .Y(_08128_));
 sky130_fd_sc_hd__nand2_2 _35950_ (.A(_08127_),
    .B(_08128_),
    .Y(_08130_));
 sky130_fd_sc_hd__nand3b_4 _35951_ (.A_N(_08122_),
    .B(_08126_),
    .C(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__inv_2 _35952_ (.A(\delay_line[23][14] ),
    .Y(_08132_));
 sky130_fd_sc_hd__o22ai_4 _35953_ (.A1(_06583_),
    .A2(_06587_),
    .B1(_08132_),
    .B2(_06603_),
    .Y(_08133_));
 sky130_fd_sc_hd__a21o_1 _35954_ (.A1(_08123_),
    .A2(_08131_),
    .B1(_08133_),
    .X(_08134_));
 sky130_fd_sc_hd__nand3_1 _35955_ (.A(_08133_),
    .B(_08123_),
    .C(_08131_),
    .Y(_08135_));
 sky130_fd_sc_hd__nand3_1 _35956_ (.A(_07644_),
    .B(_08134_),
    .C(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__a21oi_2 _35957_ (.A1(_08123_),
    .A2(_08131_),
    .B1(_08133_),
    .Y(_08137_));
 sky130_fd_sc_hd__nand2_1 _35958_ (.A(_08123_),
    .B(_08131_),
    .Y(_08138_));
 sky130_fd_sc_hd__o22a_1 _35959_ (.A1(_06583_),
    .A2(_06587_),
    .B1(_08132_),
    .B2(_06603_),
    .X(_08139_));
 sky130_fd_sc_hd__nor2_2 _35960_ (.A(_08138_),
    .B(_08139_),
    .Y(_08141_));
 sky130_fd_sc_hd__inv_2 _35961_ (.A(_07644_),
    .Y(_08142_));
 sky130_fd_sc_hd__o21ai_2 _35962_ (.A1(_08137_),
    .A2(_08141_),
    .B1(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand2_1 _35963_ (.A(_06615_),
    .B(_06616_),
    .Y(_08144_));
 sky130_fd_sc_hd__nand2_1 _35964_ (.A(_06614_),
    .B(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__a21o_1 _35965_ (.A1(_08136_),
    .A2(_08143_),
    .B1(_08145_),
    .X(_08146_));
 sky130_fd_sc_hd__o2111ai_1 _35966_ (.A1(_06606_),
    .A2(_06616_),
    .B1(_08136_),
    .C1(_08143_),
    .D1(_06615_),
    .Y(_08147_));
 sky130_fd_sc_hd__nand2_1 _35967_ (.A(_08146_),
    .B(_08147_),
    .Y(_08148_));
 sky130_fd_sc_hd__o21ai_4 _35968_ (.A1(_06620_),
    .A2(_07643_),
    .B1(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand4_1 _35969_ (.A(_06614_),
    .B(_08144_),
    .C(_08136_),
    .D(_08143_),
    .Y(_08150_));
 sky130_fd_sc_hd__nor3_1 _35970_ (.A(_08142_),
    .B(_08137_),
    .C(_08141_),
    .Y(_08152_));
 sky130_fd_sc_hd__a21oi_1 _35971_ (.A1(_08134_),
    .A2(_08135_),
    .B1(_07644_),
    .Y(_08153_));
 sky130_fd_sc_hd__o21ai_1 _35972_ (.A1(_08152_),
    .A2(_08153_),
    .B1(_08145_),
    .Y(_08154_));
 sky130_fd_sc_hd__nand2_1 _35973_ (.A(_08150_),
    .B(_08154_),
    .Y(_08155_));
 sky130_fd_sc_hd__nand3_4 _35974_ (.A(_08155_),
    .B(_06619_),
    .C(_06625_),
    .Y(_08156_));
 sky130_fd_sc_hd__nand2_1 _35975_ (.A(_08149_),
    .B(_08156_),
    .Y(_08157_));
 sky130_fd_sc_hd__clkbuf_2 _35976_ (.A(_24286_),
    .X(_08158_));
 sky130_fd_sc_hd__mux2_1 _35977_ (.A0(_08158_),
    .A1(_20261_),
    .S(_06636_),
    .X(_08159_));
 sky130_fd_sc_hd__nor2_1 _35978_ (.A(_02016_),
    .B(_06588_),
    .Y(_08160_));
 sky130_fd_sc_hd__nor2_1 _35979_ (.A(_00395_),
    .B(_08132_),
    .Y(_08161_));
 sky130_fd_sc_hd__buf_1 _35980_ (.A(_03066_),
    .X(_08163_));
 sky130_fd_sc_hd__and4bb_1 _35981_ (.A_N(_08160_),
    .B_N(_08161_),
    .C(_02015_),
    .D(_08163_),
    .X(_08164_));
 sky130_fd_sc_hd__o2bb2a_1 _35982_ (.A1_N(_02015_),
    .A2_N(_08163_),
    .B1(_08160_),
    .B2(_08161_),
    .X(_08165_));
 sky130_fd_sc_hd__nor2_1 _35983_ (.A(_08164_),
    .B(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__and2_2 _35984_ (.A(_08159_),
    .B(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__nor2_1 _35985_ (.A(_08159_),
    .B(_08166_),
    .Y(_08168_));
 sky130_fd_sc_hd__nor2_1 _35986_ (.A(_08167_),
    .B(_08168_),
    .Y(_08169_));
 sky130_fd_sc_hd__nand2_1 _35987_ (.A(_08157_),
    .B(_08169_),
    .Y(_08170_));
 sky130_fd_sc_hd__o21a_2 _35988_ (.A1(_06666_),
    .A2(_06904_),
    .B1(_06902_),
    .X(_08171_));
 sky130_fd_sc_hd__o211ai_4 _35989_ (.A1(_08167_),
    .A2(_08168_),
    .B1(_08149_),
    .C1(_08156_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand3_1 _35990_ (.A(_08170_),
    .B(_08171_),
    .C(_08172_),
    .Y(_08174_));
 sky130_fd_sc_hd__clkbuf_2 _35991_ (.A(_08174_),
    .X(_08175_));
 sky130_fd_sc_hd__nand2_2 _35992_ (.A(_08156_),
    .B(_08169_),
    .Y(_08176_));
 sky130_fd_sc_hd__o211a_1 _35993_ (.A1(_06620_),
    .A2(_07643_),
    .B1(_08150_),
    .C1(_08154_),
    .X(_08177_));
 sky130_fd_sc_hd__inv_2 _35994_ (.A(_08171_),
    .Y(_08178_));
 sky130_fd_sc_hd__o2bb2ai_1 _35995_ (.A1_N(_08149_),
    .A2_N(_08156_),
    .B1(_08167_),
    .B2(_08168_),
    .Y(_08179_));
 sky130_fd_sc_hd__o211ai_1 _35996_ (.A1(_08176_),
    .A2(_08177_),
    .B1(_08178_),
    .C1(_08179_),
    .Y(_08180_));
 sky130_fd_sc_hd__clkbuf_2 _35997_ (.A(_08180_),
    .X(_08181_));
 sky130_fd_sc_hd__nand2_1 _35998_ (.A(_07643_),
    .B(_06625_),
    .Y(_08182_));
 sky130_fd_sc_hd__a21oi_1 _35999_ (.A1(_06628_),
    .A2(_08182_),
    .B1(_06621_),
    .Y(_08183_));
 sky130_fd_sc_hd__o21ai_1 _36000_ (.A1(_07490_),
    .A2(_08183_),
    .B1(_06629_),
    .Y(_08185_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36001_ (.A(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__a21oi_1 _36002_ (.A1(_08175_),
    .A2(_08181_),
    .B1(_08186_),
    .Y(_08187_));
 sky130_fd_sc_hd__clkbuf_2 _36003_ (.A(_08187_),
    .X(_08188_));
 sky130_fd_sc_hd__nand3_1 _36004_ (.A(_08186_),
    .B(_08175_),
    .C(_08181_),
    .Y(_08189_));
 sky130_fd_sc_hd__o21a_2 _36005_ (.A1(_07474_),
    .A2(_06905_),
    .B1(_07476_),
    .X(_08190_));
 sky130_fd_sc_hd__a21bo_2 _36006_ (.A1(_06769_),
    .A2(_06900_),
    .B1_N(_06897_),
    .X(_08191_));
 sky130_fd_sc_hd__clkbuf_2 _36007_ (.A(_06752_),
    .X(_08192_));
 sky130_fd_sc_hd__buf_1 _36008_ (.A(_06751_),
    .X(_08193_));
 sky130_fd_sc_hd__and3_1 _36009_ (.A(_03663_),
    .B(_08193_),
    .C(_06752_),
    .X(_08194_));
 sky130_fd_sc_hd__a21oi_2 _36010_ (.A1(_08193_),
    .A2(_08192_),
    .B1(_03663_),
    .Y(_08196_));
 sky130_fd_sc_hd__o211ai_4 _36011_ (.A1(_06752_),
    .A2(_06757_),
    .B1(_03659_),
    .C1(_06756_),
    .Y(_08197_));
 sky130_fd_sc_hd__o221ai_4 _36012_ (.A1(_08192_),
    .A2(_06757_),
    .B1(_08194_),
    .B2(_08196_),
    .C1(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__a211o_1 _36013_ (.A1(_06758_),
    .A2(_08197_),
    .B1(_08194_),
    .C1(_08196_),
    .X(_08199_));
 sky130_fd_sc_hd__o21ai_2 _36014_ (.A1(_06762_),
    .A2(_06765_),
    .B1(_06763_),
    .Y(_08200_));
 sky130_fd_sc_hd__a21oi_1 _36015_ (.A1(_08198_),
    .A2(_08199_),
    .B1(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__and3_1 _36016_ (.A(_08198_),
    .B(_08199_),
    .C(_08200_),
    .X(_08202_));
 sky130_fd_sc_hd__a21oi_1 _36017_ (.A1(_06719_),
    .A2(_06721_),
    .B1(_06725_),
    .Y(_08203_));
 sky130_fd_sc_hd__buf_1 _36018_ (.A(\delay_line[38][12] ),
    .X(_08204_));
 sky130_fd_sc_hd__xnor2_1 _36019_ (.A(_06717_),
    .B(net284),
    .Y(_08205_));
 sky130_fd_sc_hd__and3_1 _36020_ (.A(_03642_),
    .B(_05379_),
    .C(_06719_),
    .X(_08207_));
 sky130_fd_sc_hd__a211o_1 _36021_ (.A1(_08204_),
    .A2(net284),
    .B1(_08205_),
    .C1(_08207_),
    .X(_08208_));
 sky130_fd_sc_hd__a21o_1 _36022_ (.A1(_08204_),
    .A2(net284),
    .B1(_08207_),
    .X(_08209_));
 sky130_fd_sc_hd__nand2_1 _36023_ (.A(_08209_),
    .B(_08205_),
    .Y(_08210_));
 sky130_fd_sc_hd__and3_1 _36024_ (.A(_08203_),
    .B(_08208_),
    .C(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__inv_2 _36025_ (.A(_08211_),
    .Y(_08212_));
 sky130_fd_sc_hd__a21o_1 _36026_ (.A1(_08210_),
    .A2(_08208_),
    .B1(_08203_),
    .X(_08213_));
 sky130_fd_sc_hd__buf_1 _36027_ (.A(_05360_),
    .X(_08214_));
 sky130_fd_sc_hd__clkbuf_4 _36028_ (.A(\delay_line[39][15] ),
    .X(_08215_));
 sky130_fd_sc_hd__o21bai_1 _36029_ (.A1(_08214_),
    .A2(_05362_),
    .B1_N(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__a21bo_1 _36030_ (.A1(_08214_),
    .A2(_05362_),
    .B1_N(\delay_line[39][15] ),
    .X(_08218_));
 sky130_fd_sc_hd__mux2_1 _36031_ (.A0(_08216_),
    .A1(_08218_),
    .S(_05358_),
    .X(_08219_));
 sky130_fd_sc_hd__nor2_1 _36032_ (.A(_06738_),
    .B(_06745_),
    .Y(_08220_));
 sky130_fd_sc_hd__or2_1 _36033_ (.A(_08219_),
    .B(_08220_),
    .X(_08221_));
 sky130_fd_sc_hd__or3b_1 _36034_ (.A(_06738_),
    .B(_06745_),
    .C_N(_08219_),
    .X(_08222_));
 sky130_fd_sc_hd__a22o_1 _36035_ (.A1(_08212_),
    .A2(_08213_),
    .B1(_08221_),
    .B2(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__nand4_1 _36036_ (.A(_08212_),
    .B(_08213_),
    .C(_08221_),
    .D(_08222_),
    .Y(_08224_));
 sky130_fd_sc_hd__and4bb_2 _36037_ (.A_N(_08201_),
    .B_N(_08202_),
    .C(_08223_),
    .D(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__nand2_1 _36038_ (.A(_08223_),
    .B(_08224_),
    .Y(_08226_));
 sky130_fd_sc_hd__o21a_2 _36039_ (.A1(_08201_),
    .A2(_08202_),
    .B1(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__inv_2 _36040_ (.A(_06701_),
    .Y(_08229_));
 sky130_fd_sc_hd__o21a_1 _36041_ (.A1(_08229_),
    .A2(_06708_),
    .B1(_06699_),
    .X(_08230_));
 sky130_fd_sc_hd__nor2_1 _36042_ (.A(net291),
    .B(_06706_),
    .Y(_08231_));
 sky130_fd_sc_hd__nand2_1 _36043_ (.A(_06706_),
    .B(\delay_line[37][15] ),
    .Y(_08232_));
 sky130_fd_sc_hd__and2b_1 _36044_ (.A_N(_08231_),
    .B(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__inv_2 _36045_ (.A(net291),
    .Y(_08234_));
 sky130_fd_sc_hd__or3b_1 _36046_ (.A(\delay_line[37][12] ),
    .B(_06706_),
    .C_N(_06702_),
    .X(_08235_));
 sky130_fd_sc_hd__a22oi_1 _36047_ (.A1(net291),
    .A2(_06703_),
    .B1(_06707_),
    .B2(_06705_),
    .Y(_08236_));
 sky130_fd_sc_hd__o211a_1 _36048_ (.A1(_05284_),
    .A2(_08234_),
    .B1(_08235_),
    .C1(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__xor2_1 _36049_ (.A(_08233_),
    .B(_08237_),
    .X(_08238_));
 sky130_fd_sc_hd__and2b_1 _36050_ (.A_N(_05295_),
    .B(_06670_),
    .X(_08240_));
 sky130_fd_sc_hd__and3_1 _36051_ (.A(_06671_),
    .B(_06672_),
    .C(_05298_),
    .X(_08241_));
 sky130_fd_sc_hd__xnor2_1 _36052_ (.A(_06669_),
    .B(\delay_line[36][13] ),
    .Y(_08242_));
 sky130_fd_sc_hd__o21ai_1 _36053_ (.A1(_08240_),
    .A2(_08241_),
    .B1(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__or3_1 _36054_ (.A(_08240_),
    .B(_08242_),
    .C(_08241_),
    .X(_08244_));
 sky130_fd_sc_hd__nand2_1 _36055_ (.A(_08243_),
    .B(_08244_),
    .Y(_08245_));
 sky130_fd_sc_hd__a21oi_1 _36056_ (.A1(_06670_),
    .A2(_06673_),
    .B1(_06680_),
    .Y(_08246_));
 sky130_fd_sc_hd__xnor2_1 _36057_ (.A(_08245_),
    .B(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36058_ (.A(_05320_),
    .X(_08248_));
 sky130_fd_sc_hd__buf_1 _36059_ (.A(\delay_line[35][15] ),
    .X(_08249_));
 sky130_fd_sc_hd__buf_1 _36060_ (.A(net299),
    .X(_08251_));
 sky130_fd_sc_hd__or4b_1 _36061_ (.A(_08248_),
    .B(_08249_),
    .C(_05316_),
    .D_N(_08251_),
    .X(_08252_));
 sky130_fd_sc_hd__o21ai_2 _36062_ (.A1(_08248_),
    .A2(_08249_),
    .B1(_08251_),
    .Y(_08253_));
 sky130_fd_sc_hd__a21o_1 _36063_ (.A1(_08248_),
    .A2(_08249_),
    .B1(_08251_),
    .X(_08254_));
 sky130_fd_sc_hd__a21bo_1 _36064_ (.A1(_08253_),
    .A2(_08254_),
    .B1_N(_06688_),
    .X(_08255_));
 sky130_fd_sc_hd__a21boi_1 _36065_ (.A1(_08252_),
    .A2(_08255_),
    .B1_N(_01290_),
    .Y(_08256_));
 sky130_fd_sc_hd__and3b_1 _36066_ (.A_N(_01290_),
    .B(_08252_),
    .C(_08255_),
    .X(_08257_));
 sky130_fd_sc_hd__nor2_1 _36067_ (.A(_06690_),
    .B(_06692_),
    .Y(_08258_));
 sky130_fd_sc_hd__o21a_1 _36068_ (.A1(_08256_),
    .A2(_08257_),
    .B1(_08258_),
    .X(_08259_));
 sky130_fd_sc_hd__nor3_1 _36069_ (.A(_08258_),
    .B(_08256_),
    .C(_08257_),
    .Y(_08260_));
 sky130_fd_sc_hd__clkbuf_2 _36070_ (.A(_08260_),
    .X(_08262_));
 sky130_fd_sc_hd__o32ai_2 _36071_ (.A1(net226),
    .A2(_06693_),
    .A3(_06695_),
    .B1(_08259_),
    .B2(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__or4b_1 _36072_ (.A(_06695_),
    .B(_08259_),
    .C(_08260_),
    .D_N(_06694_),
    .X(_08264_));
 sky130_fd_sc_hd__a21bo_1 _36073_ (.A1(_06697_),
    .A2(_08263_),
    .B1_N(_08264_),
    .X(_08265_));
 sky130_fd_sc_hd__o21bai_1 _36074_ (.A1(_06697_),
    .A2(_08263_),
    .B1_N(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__or2_1 _36075_ (.A(_08247_),
    .B(_08266_),
    .X(_08267_));
 sky130_fd_sc_hd__nand2_1 _36076_ (.A(_08247_),
    .B(_08266_),
    .Y(_08268_));
 sky130_fd_sc_hd__nand2_1 _36077_ (.A(_08267_),
    .B(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__or2_1 _36078_ (.A(_08238_),
    .B(_08269_),
    .X(_08270_));
 sky130_fd_sc_hd__nand2_1 _36079_ (.A(_08238_),
    .B(_08269_),
    .Y(_08271_));
 sky130_fd_sc_hd__nand2_1 _36080_ (.A(_08270_),
    .B(_08271_),
    .Y(_08273_));
 sky130_fd_sc_hd__nor2_1 _36081_ (.A(_08230_),
    .B(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__nand2_1 _36082_ (.A(_08273_),
    .B(_08230_),
    .Y(_08275_));
 sky130_fd_sc_hd__or2b_1 _36083_ (.A(_08274_),
    .B_N(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__nor3_1 _36084_ (.A(_08225_),
    .B(_08227_),
    .C(_08276_),
    .Y(_08277_));
 sky130_fd_sc_hd__o21a_1 _36085_ (.A1(_08225_),
    .A2(_08227_),
    .B1(_08276_),
    .X(_08278_));
 sky130_fd_sc_hd__or2_2 _36086_ (.A(_08277_),
    .B(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__a21bo_2 _36087_ (.A1(_06954_),
    .A2(_06984_),
    .B1_N(_06952_),
    .X(_08280_));
 sky130_fd_sc_hd__or3b_1 _36088_ (.A(_01075_),
    .B(_03737_),
    .C_N(_06795_),
    .X(_08281_));
 sky130_fd_sc_hd__inv_2 _36089_ (.A(_02880_),
    .Y(_08282_));
 sky130_fd_sc_hd__buf_1 _36090_ (.A(_06774_),
    .X(_08284_));
 sky130_fd_sc_hd__and3_1 _36091_ (.A(_08282_),
    .B(_06773_),
    .C(_08284_),
    .X(_08285_));
 sky130_fd_sc_hd__buf_1 _36092_ (.A(_06773_),
    .X(_08286_));
 sky130_fd_sc_hd__a21oi_1 _36093_ (.A1(_08286_),
    .A2(_08284_),
    .B1(_08282_),
    .Y(_08287_));
 sky130_fd_sc_hd__nor2_1 _36094_ (.A(_06774_),
    .B(_06786_),
    .Y(_08288_));
 sky130_fd_sc_hd__and2_1 _36095_ (.A(_06774_),
    .B(_06778_),
    .X(_08289_));
 sky130_fd_sc_hd__inv_2 _36096_ (.A(_06778_),
    .Y(_08290_));
 sky130_fd_sc_hd__buf_1 _36097_ (.A(net304),
    .X(_08291_));
 sky130_fd_sc_hd__or3b_2 _36098_ (.A(_08290_),
    .B(_08291_),
    .C_N(net303),
    .X(_08292_));
 sky130_fd_sc_hd__nand2_1 _36099_ (.A(_08290_),
    .B(_08291_),
    .Y(_08293_));
 sky130_fd_sc_hd__clkbuf_2 _36100_ (.A(net303),
    .X(_08295_));
 sky130_fd_sc_hd__and2b_1 _36101_ (.A_N(net303),
    .B(_08291_),
    .X(_08296_));
 sky130_fd_sc_hd__a31oi_1 _36102_ (.A1(_08292_),
    .A2(_08293_),
    .A3(_08295_),
    .B1(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__o21ai_1 _36103_ (.A1(_08288_),
    .A2(_08289_),
    .B1(_08297_),
    .Y(_08298_));
 sky130_fd_sc_hd__or3_2 _36104_ (.A(_08288_),
    .B(_08289_),
    .C(_08297_),
    .X(_08299_));
 sky130_fd_sc_hd__or2b_1 _36105_ (.A(_06781_),
    .B_N(_06784_),
    .X(_08300_));
 sky130_fd_sc_hd__and3_1 _36106_ (.A(_08298_),
    .B(_08299_),
    .C(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__a21oi_1 _36107_ (.A1(_08298_),
    .A2(_08299_),
    .B1(_08300_),
    .Y(_08302_));
 sky130_fd_sc_hd__nor2_1 _36108_ (.A(_08301_),
    .B(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__or3b_1 _36109_ (.A(_08285_),
    .B(_08287_),
    .C_N(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__nor2_1 _36110_ (.A(_08285_),
    .B(_08287_),
    .Y(_08306_));
 sky130_fd_sc_hd__or2_1 _36111_ (.A(_08306_),
    .B(_08303_),
    .X(_08307_));
 sky130_fd_sc_hd__o211a_1 _36112_ (.A1(_06790_),
    .A2(_06791_),
    .B1(_08304_),
    .C1(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__a211oi_1 _36113_ (.A1(_08304_),
    .A2(_08307_),
    .B1(_06790_),
    .C1(_06791_),
    .Y(_08309_));
 sky130_fd_sc_hd__o22a_1 _36114_ (.A1(_05165_),
    .A2(_05186_),
    .B1(_08308_),
    .B2(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__nor2_1 _36115_ (.A(_08309_),
    .B(_08308_),
    .Y(_08311_));
 sky130_fd_sc_hd__and4b_1 _36116_ (.A_N(_05186_),
    .B(_05160_),
    .C(_08286_),
    .D(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__a211o_1 _36117_ (.A1(_06793_),
    .A2(_08281_),
    .B1(_08310_),
    .C1(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__o211ai_1 _36118_ (.A1(_08310_),
    .A2(_08312_),
    .B1(_06793_),
    .C1(_08281_),
    .Y(_08314_));
 sky130_fd_sc_hd__o211a_1 _36119_ (.A1(_06798_),
    .A2(_06805_),
    .B1(_08313_),
    .C1(_08314_),
    .X(_08315_));
 sky130_fd_sc_hd__a211o_1 _36120_ (.A1(_08313_),
    .A2(_08314_),
    .B1(_06798_),
    .C1(_06805_),
    .X(_08317_));
 sky130_fd_sc_hd__and2b_1 _36121_ (.A_N(_08315_),
    .B(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__a21o_1 _36122_ (.A1(_06809_),
    .A2(_06827_),
    .B1(_06828_),
    .X(_08319_));
 sky130_fd_sc_hd__buf_1 _36123_ (.A(_05252_),
    .X(_08320_));
 sky130_fd_sc_hd__buf_1 _36124_ (.A(_24922_),
    .X(_08321_));
 sky130_fd_sc_hd__clkbuf_2 _36125_ (.A(_08321_),
    .X(_08322_));
 sky130_fd_sc_hd__a31o_1 _36126_ (.A1(_03769_),
    .A2(_08320_),
    .A3(_08322_),
    .B1(_06814_),
    .X(_08323_));
 sky130_fd_sc_hd__a21oi_1 _36127_ (.A1(_02845_),
    .A2(_08321_),
    .B1(_23357_),
    .Y(_08324_));
 sky130_fd_sc_hd__and3_1 _36128_ (.A(_23364_),
    .B(_02845_),
    .C(_08321_),
    .X(_08325_));
 sky130_fd_sc_hd__nor4b_1 _36129_ (.A(_03769_),
    .B(_08324_),
    .C(_08325_),
    .D_N(_05252_),
    .Y(_08326_));
 sky130_fd_sc_hd__inv_2 _36130_ (.A(net249),
    .Y(_08328_));
 sky130_fd_sc_hd__a2bb2o_1 _36131_ (.A1_N(_08324_),
    .A2_N(_08325_),
    .B1(_02848_),
    .B2(_08320_),
    .X(_08329_));
 sky130_fd_sc_hd__nor2_1 _36132_ (.A(_06817_),
    .B(_03774_),
    .Y(_08330_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36133_ (.A(_02838_),
    .X(_08331_));
 sky130_fd_sc_hd__nor2_1 _36134_ (.A(_02845_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__or3_1 _36135_ (.A(_08330_),
    .B(_08332_),
    .C(_06820_),
    .X(_08333_));
 sky130_fd_sc_hd__a2bb2o_1 _36136_ (.A1_N(_08330_),
    .A2_N(_08332_),
    .B1(net309),
    .B2(_06818_),
    .X(_08334_));
 sky130_fd_sc_hd__and4_1 _36137_ (.A(_08328_),
    .B(_08329_),
    .C(_08333_),
    .D(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__a22oi_2 _36138_ (.A1(_08328_),
    .A2(_08329_),
    .B1(_08333_),
    .B2(_08334_),
    .Y(_08336_));
 sky130_fd_sc_hd__nand4_1 _36139_ (.A(_06815_),
    .B(_06816_),
    .C(_06822_),
    .D(_06823_),
    .Y(_08337_));
 sky130_fd_sc_hd__o211ai_2 _36140_ (.A1(_08335_),
    .A2(_08336_),
    .B1(_06822_),
    .C1(_08337_),
    .Y(_08339_));
 sky130_fd_sc_hd__a211o_1 _36141_ (.A1(_06822_),
    .A2(_08337_),
    .B1(_08335_),
    .C1(_08336_),
    .X(_08340_));
 sky130_fd_sc_hd__and3_1 _36142_ (.A(_08323_),
    .B(_08339_),
    .C(_08340_),
    .X(_08341_));
 sky130_fd_sc_hd__a21oi_1 _36143_ (.A1(_08339_),
    .A2(_08340_),
    .B1(_08323_),
    .Y(_08342_));
 sky130_fd_sc_hd__nor2_1 _36144_ (.A(_08341_),
    .B(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__xnor2_1 _36145_ (.A(_08319_),
    .B(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__and4bb_1 _36146_ (.A_N(_06830_),
    .B_N(_08344_),
    .C(_06831_),
    .D(_06808_),
    .X(_08345_));
 sky130_fd_sc_hd__a21boi_1 _36147_ (.A1(_06808_),
    .A2(_06833_),
    .B1_N(_08344_),
    .Y(_08346_));
 sky130_fd_sc_hd__nor2_1 _36148_ (.A(_08345_),
    .B(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__inv_2 _36149_ (.A(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__a21oi_1 _36150_ (.A1(_06838_),
    .A2(_06837_),
    .B1(_06835_),
    .Y(_08350_));
 sky130_fd_sc_hd__nor2_1 _36151_ (.A(_08348_),
    .B(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__a211o_1 _36152_ (.A1(_06838_),
    .A2(_06837_),
    .B1(_06835_),
    .C1(_08347_),
    .X(_08352_));
 sky130_fd_sc_hd__and2b_1 _36153_ (.A_N(_08351_),
    .B(_08352_),
    .X(_08353_));
 sky130_fd_sc_hd__a21oi_1 _36154_ (.A1(_05192_),
    .A2(_05225_),
    .B1(_06873_),
    .Y(_08354_));
 sky130_fd_sc_hd__a21oi_1 _36155_ (.A1(_05234_),
    .A2(_05230_),
    .B1(_06881_),
    .Y(_08355_));
 sky130_fd_sc_hd__and3_1 _36156_ (.A(_06873_),
    .B(_05192_),
    .C(_05225_),
    .X(_08356_));
 sky130_fd_sc_hd__o21bai_1 _36157_ (.A1(_08354_),
    .A2(_08355_),
    .B1_N(_08356_),
    .Y(_08357_));
 sky130_fd_sc_hd__xor2_2 _36158_ (.A(_21116_),
    .B(_02795_),
    .X(_08358_));
 sky130_fd_sc_hd__xnor2_1 _36159_ (.A(_24971_),
    .B(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__a21oi_1 _36160_ (.A1(_05197_),
    .A2(_06847_),
    .B1(_05195_),
    .Y(_08361_));
 sky130_fd_sc_hd__a211oi_2 _36161_ (.A1(_06855_),
    .A2(_06856_),
    .B1(_06851_),
    .C1(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__o21a_1 _36162_ (.A1(_06851_),
    .A2(_06857_),
    .B1(_08361_),
    .X(_08363_));
 sky130_fd_sc_hd__or3_2 _36163_ (.A(_08359_),
    .B(_08362_),
    .C(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__o21ai_2 _36164_ (.A1(_08362_),
    .A2(_08363_),
    .B1(_08359_),
    .Y(_08365_));
 sky130_fd_sc_hd__nor4_1 _36165_ (.A(_06842_),
    .B(_06844_),
    .C(_06859_),
    .D(_06860_),
    .Y(_08366_));
 sky130_fd_sc_hd__or2_1 _36166_ (.A(_06859_),
    .B(_08366_),
    .X(_08367_));
 sky130_fd_sc_hd__and3_1 _36167_ (.A(_08364_),
    .B(_08365_),
    .C(_08367_),
    .X(_08368_));
 sky130_fd_sc_hd__a21oi_1 _36168_ (.A1(_08364_),
    .A2(_08365_),
    .B1(_08367_),
    .Y(_08369_));
 sky130_fd_sc_hd__nor2_2 _36169_ (.A(_08368_),
    .B(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__xnor2_2 _36170_ (.A(_06842_),
    .B(_08370_),
    .Y(_08372_));
 sky130_fd_sc_hd__o21a_1 _36171_ (.A1(_05214_),
    .A2(_06863_),
    .B1(_06864_),
    .X(_08373_));
 sky130_fd_sc_hd__xor2_1 _36172_ (.A(_08372_),
    .B(_08373_),
    .X(_08374_));
 sky130_fd_sc_hd__xnor2_1 _36173_ (.A(_06872_),
    .B(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__xnor2_1 _36174_ (.A(_08357_),
    .B(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__xor2_1 _36175_ (.A(_08353_),
    .B(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__xor2_1 _36176_ (.A(_08318_),
    .B(_08377_),
    .X(_08378_));
 sky130_fd_sc_hd__xnor2_1 _36177_ (.A(_08280_),
    .B(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__o21ba_1 _36178_ (.A1(_06806_),
    .A2(_06884_),
    .B1_N(_06885_),
    .X(_08380_));
 sky130_fd_sc_hd__xor2_1 _36179_ (.A(_08379_),
    .B(_08380_),
    .X(_08381_));
 sky130_fd_sc_hd__a21o_1 _36180_ (.A1(_06891_),
    .A2(_06893_),
    .B1(_06889_),
    .X(_08383_));
 sky130_fd_sc_hd__nand2_2 _36181_ (.A(_08381_),
    .B(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__a211o_1 _36182_ (.A1(_06893_),
    .A2(_06891_),
    .B1(_06889_),
    .C1(_08381_),
    .X(_08385_));
 sky130_fd_sc_hd__nand3b_1 _36183_ (.A_N(_08279_),
    .B(_08384_),
    .C(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__a21bo_1 _36184_ (.A1(_08384_),
    .A2(_08385_),
    .B1_N(_08279_),
    .X(_08387_));
 sky130_fd_sc_hd__a21o_1 _36185_ (.A1(_07070_),
    .A2(_07069_),
    .B1(_07073_),
    .X(_08388_));
 sky130_fd_sc_hd__a21oi_1 _36186_ (.A1(_08386_),
    .A2(_08387_),
    .B1(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__and3_1 _36187_ (.A(_08388_),
    .B(_08386_),
    .C(_08387_),
    .X(_08390_));
 sky130_fd_sc_hd__nor2_1 _36188_ (.A(_08389_),
    .B(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__or2_1 _36189_ (.A(_08191_),
    .B(_08391_),
    .X(_08392_));
 sky130_fd_sc_hd__nand2_1 _36190_ (.A(_08391_),
    .B(_08191_),
    .Y(_08394_));
 sky130_fd_sc_hd__a21oi_2 _36191_ (.A1(_05989_),
    .A2(_07469_),
    .B1(_07473_),
    .Y(_08395_));
 sky130_fd_sc_hd__o22ai_4 _36192_ (.A1(_07463_),
    .A2(_07465_),
    .B1(_07202_),
    .B2(_07467_),
    .Y(_08396_));
 sky130_fd_sc_hd__o21a_4 _36193_ (.A1(_07374_),
    .A2(_07461_),
    .B1(_07460_),
    .X(_08397_));
 sky130_fd_sc_hd__or2_1 _36194_ (.A(_07077_),
    .B(_07103_),
    .X(_08398_));
 sky130_fd_sc_hd__buf_1 _36195_ (.A(_05888_),
    .X(_08399_));
 sky130_fd_sc_hd__nand4b_1 _36196_ (.A_N(_08399_),
    .B(_07104_),
    .C(_18322_),
    .D(_05889_),
    .Y(_08400_));
 sky130_fd_sc_hd__buf_1 _36197_ (.A(_05880_),
    .X(_08401_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36198_ (.A(_08401_),
    .X(_08402_));
 sky130_fd_sc_hd__and2b_1 _36199_ (.A_N(_08402_),
    .B(_05889_),
    .X(_08403_));
 sky130_fd_sc_hd__inv_2 _36200_ (.A(_05878_),
    .Y(_08405_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36201_ (.A(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__nand3_1 _36202_ (.A(_08406_),
    .B(_08401_),
    .C(_05888_),
    .Y(_08407_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36203_ (.A(_05878_),
    .X(_08408_));
 sky130_fd_sc_hd__o2111ai_2 _36204_ (.A1(_05880_),
    .A2(_08408_),
    .B1(_07091_),
    .C1(_07093_),
    .D1(_07094_),
    .Y(_08409_));
 sky130_fd_sc_hd__inv_2 _36205_ (.A(_05871_),
    .Y(_08410_));
 sky130_fd_sc_hd__clkbuf_2 _36206_ (.A(_05863_),
    .X(_08411_));
 sky130_fd_sc_hd__or2_1 _36207_ (.A(net340),
    .B(\delay_line[25][15] ),
    .X(_08412_));
 sky130_fd_sc_hd__nand2_1 _36208_ (.A(_05863_),
    .B(_07081_),
    .Y(_08413_));
 sky130_fd_sc_hd__a22o_2 _36209_ (.A1(_05868_),
    .A2(_07081_),
    .B1(_08412_),
    .B2(_08413_),
    .X(_08414_));
 sky130_fd_sc_hd__o211ai_4 _36210_ (.A1(_08411_),
    .A2(_07082_),
    .B1(_05867_),
    .C1(_08414_),
    .Y(_08416_));
 sky130_fd_sc_hd__inv_2 _36211_ (.A(\delay_line[25][13] ),
    .Y(_08417_));
 sky130_fd_sc_hd__or3b_2 _36212_ (.A(_08417_),
    .B(_05863_),
    .C_N(_07081_),
    .X(_08418_));
 sky130_fd_sc_hd__a21o_1 _36213_ (.A1(_08418_),
    .A2(_08414_),
    .B1(_05867_),
    .X(_08419_));
 sky130_fd_sc_hd__nand2_1 _36214_ (.A(_07087_),
    .B(_07090_),
    .Y(_08420_));
 sky130_fd_sc_hd__and3_1 _36215_ (.A(_08416_),
    .B(_08419_),
    .C(_08420_),
    .X(_08421_));
 sky130_fd_sc_hd__a21oi_1 _36216_ (.A1(_08416_),
    .A2(_08419_),
    .B1(_08420_),
    .Y(_08422_));
 sky130_fd_sc_hd__nor3_1 _36217_ (.A(_22816_),
    .B(_08405_),
    .C(_22813_),
    .Y(_08423_));
 sky130_fd_sc_hd__a2111oi_2 _36218_ (.A1(_08406_),
    .A2(_08410_),
    .B1(_08421_),
    .C1(_08422_),
    .D1(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__o21ai_1 _36219_ (.A1(_22813_),
    .A2(_22816_),
    .B1(_05878_),
    .Y(_08425_));
 sky130_fd_sc_hd__o221a_1 _36220_ (.A1(_08410_),
    .A2(_08408_),
    .B1(_08422_),
    .B2(_08421_),
    .C1(_08425_),
    .X(_08427_));
 sky130_fd_sc_hd__a211oi_2 _36221_ (.A1(_07092_),
    .A2(_08409_),
    .B1(_08424_),
    .C1(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__o211a_1 _36222_ (.A1(_08424_),
    .A2(_08427_),
    .B1(_07092_),
    .C1(_08409_),
    .X(_08429_));
 sky130_fd_sc_hd__o2bb2a_1 _36223_ (.A1_N(_08401_),
    .A2_N(_08407_),
    .B1(_08428_),
    .B2(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__and4bb_1 _36224_ (.A_N(_08429_),
    .B_N(_08428_),
    .C(_08407_),
    .D(_08401_),
    .X(_08431_));
 sky130_fd_sc_hd__nor2_1 _36225_ (.A(_08430_),
    .B(_08431_),
    .Y(_08432_));
 sky130_fd_sc_hd__or3_1 _36226_ (.A(_07098_),
    .B(_07100_),
    .C(_07097_),
    .X(_08433_));
 sky130_fd_sc_hd__o21ai_1 _36227_ (.A1(_07078_),
    .A2(_07102_),
    .B1(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__and2_1 _36228_ (.A(_08432_),
    .B(_08434_),
    .X(_08435_));
 sky130_fd_sc_hd__nor2_1 _36229_ (.A(_08434_),
    .B(_08432_),
    .Y(_08436_));
 sky130_fd_sc_hd__nor2_1 _36230_ (.A(_08435_),
    .B(_08436_),
    .Y(_08438_));
 sky130_fd_sc_hd__nand3_1 _36231_ (.A(_08399_),
    .B(_08403_),
    .C(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__a21o_1 _36232_ (.A1(_05888_),
    .A2(_08403_),
    .B1(_08438_),
    .X(_08440_));
 sky130_fd_sc_hd__nand2_1 _36233_ (.A(_08439_),
    .B(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__a21oi_1 _36234_ (.A1(_08398_),
    .A2(_08400_),
    .B1(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__and3_1 _36235_ (.A(_08398_),
    .B(_08400_),
    .C(_08441_),
    .X(_08443_));
 sky130_fd_sc_hd__nor2_1 _36236_ (.A(_08442_),
    .B(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__nor2_1 _36237_ (.A(_07076_),
    .B(_07105_),
    .Y(_08445_));
 sky130_fd_sc_hd__a21oi_2 _36238_ (.A1(_07108_),
    .A2(_07106_),
    .B1(_08445_),
    .Y(_08446_));
 sky130_fd_sc_hd__xnor2_2 _36239_ (.A(_08444_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__and3b_1 _36240_ (.A_N(_07115_),
    .B(_20450_),
    .C(_20454_),
    .X(_08449_));
 sky130_fd_sc_hd__buf_1 _36241_ (.A(_04177_),
    .X(_08450_));
 sky130_fd_sc_hd__a21oi_1 _36242_ (.A1(_07113_),
    .A2(_07115_),
    .B1(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__and3_1 _36243_ (.A(_07113_),
    .B(_02363_),
    .C(_04177_),
    .X(_08452_));
 sky130_fd_sc_hd__buf_1 _36244_ (.A(\delay_line[22][11] ),
    .X(_08453_));
 sky130_fd_sc_hd__or2_1 _36245_ (.A(_08453_),
    .B(net350),
    .X(_08454_));
 sky130_fd_sc_hd__nand2_1 _36246_ (.A(_08453_),
    .B(net350),
    .Y(_08455_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36247_ (.A(net351),
    .X(_08456_));
 sky130_fd_sc_hd__nand4_1 _36248_ (.A(_08454_),
    .B(_08455_),
    .C(_00518_),
    .D(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__a22o_1 _36249_ (.A1(_00518_),
    .A2(net351),
    .B1(_08454_),
    .B2(_08455_),
    .X(_08458_));
 sky130_fd_sc_hd__or4bb_1 _36250_ (.A(_08451_),
    .B(_08452_),
    .C_N(_08457_),
    .D_N(_08458_),
    .X(_08460_));
 sky130_fd_sc_hd__a2bb2o_1 _36251_ (.A1_N(_08451_),
    .A2_N(_08452_),
    .B1(_08457_),
    .B2(_08458_),
    .X(_08461_));
 sky130_fd_sc_hd__nand2_1 _36252_ (.A(_07123_),
    .B(_07125_),
    .Y(_08462_));
 sky130_fd_sc_hd__a21oi_1 _36253_ (.A1(_08460_),
    .A2(_08461_),
    .B1(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__and3_1 _36254_ (.A(_08462_),
    .B(_08460_),
    .C(_08461_),
    .X(_08464_));
 sky130_fd_sc_hd__nor4_1 _36255_ (.A(_07132_),
    .B(_08449_),
    .C(_08463_),
    .D(_08464_),
    .Y(_08465_));
 sky130_fd_sc_hd__o22a_1 _36256_ (.A1(_07132_),
    .A2(_08449_),
    .B1(_08463_),
    .B2(_08464_),
    .X(_08466_));
 sky130_fd_sc_hd__nor2_1 _36257_ (.A(_08465_),
    .B(_08466_),
    .Y(_08467_));
 sky130_fd_sc_hd__a311o_1 _36258_ (.A1(_07127_),
    .A2(_07125_),
    .A3(_07126_),
    .B1(_07133_),
    .C1(_08467_),
    .X(_08468_));
 sky130_fd_sc_hd__o21ai_1 _36259_ (.A1(_07130_),
    .A2(_07133_),
    .B1(_08467_),
    .Y(_08469_));
 sky130_fd_sc_hd__and2_1 _36260_ (.A(_08468_),
    .B(_08469_),
    .X(_08471_));
 sky130_fd_sc_hd__xor2_1 _36261_ (.A(_07114_),
    .B(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__o21a_1 _36262_ (.A1(_07136_),
    .A2(_07137_),
    .B1(_08472_),
    .X(_08473_));
 sky130_fd_sc_hd__nor3_1 _36263_ (.A(_07136_),
    .B(_07137_),
    .C(_08472_),
    .Y(_08474_));
 sky130_fd_sc_hd__nor2_1 _36264_ (.A(_08473_),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__o21a_1 _36265_ (.A1(_07139_),
    .A2(_07146_),
    .B1(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__or3_1 _36266_ (.A(_07139_),
    .B(_07146_),
    .C(_08475_),
    .X(_08477_));
 sky130_fd_sc_hd__or2b_1 _36267_ (.A(_08476_),
    .B_N(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__o21ai_2 _36268_ (.A1(_02317_),
    .A2(_04213_),
    .B1(_00551_),
    .Y(_08479_));
 sky130_fd_sc_hd__and2_1 _36269_ (.A(_07153_),
    .B(net341),
    .X(_08480_));
 sky130_fd_sc_hd__inv_2 _36270_ (.A(\delay_line[24][15] ),
    .Y(_08482_));
 sky130_fd_sc_hd__nor2_2 _36271_ (.A(_07153_),
    .B(_04213_),
    .Y(_08483_));
 sky130_fd_sc_hd__inv_2 _36272_ (.A(_00559_),
    .Y(_08484_));
 sky130_fd_sc_hd__o21ai_1 _36273_ (.A1(_08480_),
    .A2(_08483_),
    .B1(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__o211ai_1 _36274_ (.A1(_08479_),
    .A2(_08480_),
    .B1(_08482_),
    .C1(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__o21ai_2 _36275_ (.A1(_08480_),
    .A2(_08479_),
    .B1(_08485_),
    .Y(_08487_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36276_ (.A(\delay_line[24][15] ),
    .X(_08488_));
 sky130_fd_sc_hd__nand2_1 _36277_ (.A(_08487_),
    .B(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__a21o_1 _36278_ (.A1(_08486_),
    .A2(_08489_),
    .B1(_07160_),
    .X(_08490_));
 sky130_fd_sc_hd__o21a_1 _36279_ (.A1(_00560_),
    .A2(_02322_),
    .B1(_05957_),
    .X(_08491_));
 sky130_fd_sc_hd__o21ba_1 _36280_ (.A1(_05957_),
    .A2(_07155_),
    .B1_N(_08491_),
    .X(_08493_));
 sky130_fd_sc_hd__nand3_1 _36281_ (.A(_07160_),
    .B(_08486_),
    .C(_08489_),
    .Y(_08494_));
 sky130_fd_sc_hd__nand3_1 _36282_ (.A(_08490_),
    .B(_08493_),
    .C(_08494_),
    .Y(_08495_));
 sky130_fd_sc_hd__a21o_1 _36283_ (.A1(_08494_),
    .A2(_08490_),
    .B1(_08493_),
    .X(_08496_));
 sky130_fd_sc_hd__nand2_1 _36284_ (.A(_07163_),
    .B(_07172_),
    .Y(_08497_));
 sky130_fd_sc_hd__a21o_1 _36285_ (.A1(_08495_),
    .A2(_08496_),
    .B1(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__nand3_1 _36286_ (.A(_08497_),
    .B(_08495_),
    .C(_08496_),
    .Y(_08499_));
 sky130_fd_sc_hd__o211a_1 _36287_ (.A1(_07166_),
    .A2(_07167_),
    .B1(_04225_),
    .C1(_07171_),
    .X(_08500_));
 sky130_fd_sc_hd__nor2_1 _36288_ (.A(_04225_),
    .B(_07169_),
    .Y(_08501_));
 sky130_fd_sc_hd__nor2_1 _36289_ (.A(_08500_),
    .B(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__nand3_1 _36290_ (.A(_08498_),
    .B(_08499_),
    .C(_08502_),
    .Y(_08504_));
 sky130_fd_sc_hd__a21o_1 _36291_ (.A1(_08498_),
    .A2(_08499_),
    .B1(_08502_),
    .X(_08505_));
 sky130_fd_sc_hd__and2_1 _36292_ (.A(_08504_),
    .B(_08505_),
    .X(_08506_));
 sky130_fd_sc_hd__o21ai_1 _36293_ (.A1(_07149_),
    .A2(_07176_),
    .B1(_07174_),
    .Y(_08507_));
 sky130_fd_sc_hd__xnor2_1 _36294_ (.A(_08506_),
    .B(_08507_),
    .Y(_08508_));
 sky130_fd_sc_hd__nor2_1 _36295_ (.A(_07147_),
    .B(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__o31a_1 _36296_ (.A1(_02336_),
    .A2(_04211_),
    .A3(_04207_),
    .B1(_08508_),
    .X(_08510_));
 sky130_fd_sc_hd__nor2_1 _36297_ (.A(_08509_),
    .B(_08510_),
    .Y(_08511_));
 sky130_fd_sc_hd__nor3_1 _36298_ (.A(_07178_),
    .B(_07182_),
    .C(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__o21a_1 _36299_ (.A1(_07178_),
    .A2(_07182_),
    .B1(_08511_),
    .X(_08513_));
 sky130_fd_sc_hd__nor2_1 _36300_ (.A(_08512_),
    .B(_08513_),
    .Y(_08515_));
 sky130_fd_sc_hd__o22ai_4 _36301_ (.A1(_07183_),
    .A2(_07180_),
    .B1(_07185_),
    .B2(_07188_),
    .Y(_08516_));
 sky130_fd_sc_hd__xor2_2 _36302_ (.A(_08515_),
    .B(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__xnor2_2 _36303_ (.A(_08478_),
    .B(_08517_),
    .Y(_08518_));
 sky130_fd_sc_hd__xnor2_2 _36304_ (.A(_08447_),
    .B(_08518_),
    .Y(_08519_));
 sky130_fd_sc_hd__xor2_1 _36305_ (.A(_08397_),
    .B(_08519_),
    .X(_08520_));
 sky130_fd_sc_hd__o21ai_1 _36306_ (.A1(_07190_),
    .A2(_07193_),
    .B1(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__or3_1 _36307_ (.A(_07190_),
    .B(_07193_),
    .C(_08520_),
    .X(_08522_));
 sky130_fd_sc_hd__and2_1 _36308_ (.A(_08521_),
    .B(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__inv_2 _36309_ (.A(_08523_),
    .Y(_08524_));
 sky130_fd_sc_hd__o21ba_1 _36310_ (.A1(_07243_),
    .A2(_07315_),
    .B1_N(_07314_),
    .X(_08526_));
 sky130_fd_sc_hd__nand2_1 _36311_ (.A(_07227_),
    .B(_07232_),
    .Y(_08527_));
 sky130_fd_sc_hd__or4bb_1 _36312_ (.A(_07203_),
    .B(_07204_),
    .C_N(_07223_),
    .D_N(_07224_),
    .X(_08528_));
 sky130_fd_sc_hd__buf_1 _36313_ (.A(_05752_),
    .X(_08529_));
 sky130_fd_sc_hd__and3_1 _36314_ (.A(_05740_),
    .B(_08529_),
    .C(_03874_),
    .X(_08530_));
 sky130_fd_sc_hd__a21oi_1 _36315_ (.A1(_05740_),
    .A2(_08529_),
    .B1(_03874_),
    .Y(_08531_));
 sky130_fd_sc_hd__a21o_1 _36316_ (.A1(_00834_),
    .A2(_02494_),
    .B1(_05753_),
    .X(_08532_));
 sky130_fd_sc_hd__o21ai_1 _36317_ (.A1(_05739_),
    .A2(_07207_),
    .B1(_08532_),
    .Y(_08533_));
 sky130_fd_sc_hd__and3_1 _36318_ (.A(_07212_),
    .B(\delay_line[16][14] ),
    .C(_07209_),
    .X(_08534_));
 sky130_fd_sc_hd__clkbuf_2 _36319_ (.A(\delay_line[16][12] ),
    .X(_08535_));
 sky130_fd_sc_hd__o21ai_2 _36320_ (.A1(_02489_),
    .A2(_08535_),
    .B1(_00828_),
    .Y(_08537_));
 sky130_fd_sc_hd__and2_1 _36321_ (.A(net381),
    .B(\delay_line[16][12] ),
    .X(_08538_));
 sky130_fd_sc_hd__inv_2 _36322_ (.A(net379),
    .Y(_08539_));
 sky130_fd_sc_hd__nor2_2 _36323_ (.A(_02489_),
    .B(_08535_),
    .Y(_08540_));
 sky130_fd_sc_hd__o21ai_1 _36324_ (.A1(_08538_),
    .A2(_08540_),
    .B1(_02498_),
    .Y(_08541_));
 sky130_fd_sc_hd__o211a_1 _36325_ (.A1(_08537_),
    .A2(_08538_),
    .B1(_08539_),
    .C1(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__o21ai_2 _36326_ (.A1(_08538_),
    .A2(_08537_),
    .B1(_08541_),
    .Y(_08543_));
 sky130_fd_sc_hd__and2_1 _36327_ (.A(_08543_),
    .B(net379),
    .X(_08544_));
 sky130_fd_sc_hd__nor3_1 _36328_ (.A(_08534_),
    .B(_08542_),
    .C(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__o21a_1 _36329_ (.A1(_08542_),
    .A2(_08544_),
    .B1(_08534_),
    .X(_08546_));
 sky130_fd_sc_hd__or3_1 _36330_ (.A(_08533_),
    .B(_08545_),
    .C(_08546_),
    .X(_08548_));
 sky130_fd_sc_hd__o21ai_2 _36331_ (.A1(_08545_),
    .A2(_08546_),
    .B1(_08533_),
    .Y(_08549_));
 sky130_fd_sc_hd__and3_1 _36332_ (.A(_07213_),
    .B(_05746_),
    .C(_07215_),
    .X(_08550_));
 sky130_fd_sc_hd__and3_1 _36333_ (.A(_07216_),
    .B(_07218_),
    .C(_07220_),
    .X(_08551_));
 sky130_fd_sc_hd__a211oi_2 _36334_ (.A1(_08548_),
    .A2(_08549_),
    .B1(_08550_),
    .C1(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__o211ai_2 _36335_ (.A1(_08550_),
    .A2(_08551_),
    .B1(_08548_),
    .C1(_08549_),
    .Y(_08553_));
 sky130_fd_sc_hd__inv_2 _36336_ (.A(_08553_),
    .Y(_08554_));
 sky130_fd_sc_hd__nor4_1 _36337_ (.A(_08530_),
    .B(_08531_),
    .C(_08552_),
    .D(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__o22a_1 _36338_ (.A1(_08530_),
    .A2(_08531_),
    .B1(_08552_),
    .B2(_08554_),
    .X(_08556_));
 sky130_fd_sc_hd__a211o_1 _36339_ (.A1(_07223_),
    .A2(_08528_),
    .B1(_08555_),
    .C1(_08556_),
    .X(_08557_));
 sky130_fd_sc_hd__o211ai_1 _36340_ (.A1(_08555_),
    .A2(_08556_),
    .B1(_07223_),
    .C1(_08528_),
    .Y(_08559_));
 sky130_fd_sc_hd__nand4_1 _36341_ (.A(_08557_),
    .B(_03901_),
    .C(_08559_),
    .D(_05758_),
    .Y(_08560_));
 sky130_fd_sc_hd__a22o_1 _36342_ (.A1(_03901_),
    .A2(_05758_),
    .B1(_08559_),
    .B2(_08557_),
    .X(_08561_));
 sky130_fd_sc_hd__nand2_1 _36343_ (.A(_08560_),
    .B(_08561_),
    .Y(_08562_));
 sky130_fd_sc_hd__xnor2_1 _36344_ (.A(_08527_),
    .B(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__o21ai_2 _36345_ (.A1(_07236_),
    .A2(_07242_),
    .B1(_07237_),
    .Y(_08564_));
 sky130_fd_sc_hd__xnor2_1 _36346_ (.A(_08563_),
    .B(_08564_),
    .Y(_08565_));
 sky130_fd_sc_hd__o21bai_1 _36347_ (.A1(_07308_),
    .A2(_07309_),
    .B1_N(_07307_),
    .Y(_08566_));
 sky130_fd_sc_hd__and3_1 _36348_ (.A(_03923_),
    .B(_07286_),
    .C(_02405_),
    .X(_08567_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36349_ (.A(_07286_),
    .X(_08568_));
 sky130_fd_sc_hd__clkbuf_2 _36350_ (.A(_02405_),
    .X(_08570_));
 sky130_fd_sc_hd__a21oi_1 _36351_ (.A1(_08568_),
    .A2(_08570_),
    .B1(_03923_),
    .Y(_08571_));
 sky130_fd_sc_hd__inv_2 _36352_ (.A(net388),
    .Y(_08572_));
 sky130_fd_sc_hd__xor2_2 _36353_ (.A(_00749_),
    .B(\delay_line[14][11] ),
    .X(_08573_));
 sky130_fd_sc_hd__xor2_1 _36354_ (.A(_08572_),
    .B(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__or4b_1 _36355_ (.A(_07289_),
    .B(_07290_),
    .C(_08574_),
    .D_N(\delay_line[14][14] ),
    .X(_08575_));
 sky130_fd_sc_hd__nand2_1 _36356_ (.A(_08574_),
    .B(_07291_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand2_1 _36357_ (.A(_08575_),
    .B(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__or3_2 _36358_ (.A(_08567_),
    .B(_08571_),
    .C(_08577_),
    .X(_08578_));
 sky130_fd_sc_hd__o21ai_1 _36359_ (.A1(_08567_),
    .A2(_08571_),
    .B1(_08577_),
    .Y(_08579_));
 sky130_fd_sc_hd__or2b_1 _36360_ (.A(_07296_),
    .B_N(_07298_),
    .X(_08581_));
 sky130_fd_sc_hd__a21oi_1 _36361_ (.A1(_08578_),
    .A2(_08579_),
    .B1(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__and3_1 _36362_ (.A(_08581_),
    .B(_08578_),
    .C(_08579_),
    .X(_08583_));
 sky130_fd_sc_hd__nor2_1 _36363_ (.A(_08582_),
    .B(_08583_),
    .Y(_08584_));
 sky130_fd_sc_hd__xor2_1 _36364_ (.A(_07288_),
    .B(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__a21bo_1 _36365_ (.A1(_07302_),
    .A2(_05787_),
    .B1_N(_07303_),
    .X(_08586_));
 sky130_fd_sc_hd__nand2_1 _36366_ (.A(_08585_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__or2_1 _36367_ (.A(_08586_),
    .B(_08585_),
    .X(_08588_));
 sky130_fd_sc_hd__and3_2 _36368_ (.A(_08566_),
    .B(_08587_),
    .C(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__a211o_1 _36369_ (.A1(_08587_),
    .A2(_08588_),
    .B1(_07307_),
    .C1(_07310_),
    .X(_08590_));
 sky130_fd_sc_hd__inv_2 _36370_ (.A(_08590_),
    .Y(_08592_));
 sky130_fd_sc_hd__nand2_1 _36371_ (.A(_07267_),
    .B(_07269_),
    .Y(_08593_));
 sky130_fd_sc_hd__clkbuf_2 _36372_ (.A(_03960_),
    .X(_08594_));
 sky130_fd_sc_hd__or3b_2 _36373_ (.A(_08594_),
    .B(_05823_),
    .C_N(_05801_),
    .X(_08595_));
 sky130_fd_sc_hd__and2_1 _36374_ (.A(_24745_),
    .B(_07258_),
    .X(_08596_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36375_ (.A(_00781_),
    .X(_08597_));
 sky130_fd_sc_hd__buf_1 _36376_ (.A(_03954_),
    .X(_08598_));
 sky130_fd_sc_hd__or3b_1 _36377_ (.A(_08598_),
    .B(_07255_),
    .C_N(_07249_),
    .X(_08599_));
 sky130_fd_sc_hd__nand2_2 _36378_ (.A(_07252_),
    .B(_07255_),
    .Y(_08600_));
 sky130_fd_sc_hd__o211a_1 _36379_ (.A1(_05805_),
    .A2(_07249_),
    .B1(_08599_),
    .C1(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__nand2_2 _36380_ (.A(_08597_),
    .B(_08601_),
    .Y(_08603_));
 sky130_fd_sc_hd__or2_1 _36381_ (.A(_08597_),
    .B(_08601_),
    .X(_08604_));
 sky130_fd_sc_hd__o211ai_4 _36382_ (.A1(_07253_),
    .A2(_08596_),
    .B1(_08603_),
    .C1(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__nor2_1 _36383_ (.A(_07251_),
    .B(_07252_),
    .Y(_08606_));
 sky130_fd_sc_hd__a221o_1 _36384_ (.A1(_05809_),
    .A2(_08606_),
    .B1(_08603_),
    .B2(_08604_),
    .C1(_08596_),
    .X(_08607_));
 sky130_fd_sc_hd__or3b_2 _36385_ (.A(_23075_),
    .B(_23079_),
    .C_N(_08594_),
    .X(_08608_));
 sky130_fd_sc_hd__or2_1 _36386_ (.A(_08594_),
    .B(_05813_),
    .X(_08609_));
 sky130_fd_sc_hd__a22o_1 _36387_ (.A1(_08605_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__clkbuf_2 _36388_ (.A(_05813_),
    .X(_08611_));
 sky130_fd_sc_hd__o2111ai_4 _36389_ (.A1(_08594_),
    .A2(_08611_),
    .B1(_08605_),
    .C1(_08607_),
    .D1(_08608_),
    .Y(_08612_));
 sky130_fd_sc_hd__and3_1 _36390_ (.A(_07248_),
    .B(_07257_),
    .C(_07259_),
    .X(_08614_));
 sky130_fd_sc_hd__a221o_1 _36391_ (.A1(_07264_),
    .A2(_07262_),
    .B1(_08610_),
    .B2(_08612_),
    .C1(_08614_),
    .X(_08615_));
 sky130_fd_sc_hd__o211ai_4 _36392_ (.A1(_08614_),
    .A2(_07265_),
    .B1(_08612_),
    .C1(_08610_),
    .Y(_08616_));
 sky130_fd_sc_hd__a22o_1 _36393_ (.A1(_08595_),
    .A2(_05819_),
    .B1(_08615_),
    .B2(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__nand4_2 _36394_ (.A(_08615_),
    .B(_08616_),
    .C(_08595_),
    .D(_05819_),
    .Y(_08618_));
 sky130_fd_sc_hd__nand3_2 _36395_ (.A(_08593_),
    .B(_08617_),
    .C(_08618_),
    .Y(_08619_));
 sky130_fd_sc_hd__inv_2 _36396_ (.A(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__a21oi_1 _36397_ (.A1(_08617_),
    .A2(_08618_),
    .B1(_08593_),
    .Y(_08621_));
 sky130_fd_sc_hd__o2bb2a_1 _36398_ (.A1_N(_07246_),
    .A2_N(_20603_),
    .B1(_08620_),
    .B2(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__o21bai_1 _36399_ (.A1(_05802_),
    .A2(_07273_),
    .B1_N(_07271_),
    .Y(_08623_));
 sky130_fd_sc_hd__or4bb_1 _36400_ (.A(_08621_),
    .B(_20597_),
    .C_N(_07246_),
    .D_N(_08619_),
    .X(_08625_));
 sky130_fd_sc_hd__nand2_1 _36401_ (.A(_08623_),
    .B(_08625_),
    .Y(_08626_));
 sky130_fd_sc_hd__and4b_1 _36402_ (.A_N(_08621_),
    .B(_20603_),
    .C(_07246_),
    .D(_08619_),
    .X(_08627_));
 sky130_fd_sc_hd__o21bai_1 _36403_ (.A1(_08622_),
    .A2(_08627_),
    .B1_N(_08623_),
    .Y(_08628_));
 sky130_fd_sc_hd__o21ai_1 _36404_ (.A1(_08622_),
    .A2(_08626_),
    .B1(_08628_),
    .Y(_08629_));
 sky130_fd_sc_hd__a21boi_1 _36405_ (.A1(_07280_),
    .A2(_07278_),
    .B1_N(_07276_),
    .Y(_08630_));
 sky130_fd_sc_hd__xnor2_1 _36406_ (.A(_08629_),
    .B(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__or3_1 _36407_ (.A(_08589_),
    .B(_08592_),
    .C(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__o21ai_1 _36408_ (.A1(_08589_),
    .A2(_08592_),
    .B1(_08631_),
    .Y(_08633_));
 sky130_fd_sc_hd__nand2_1 _36409_ (.A(_08632_),
    .B(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__and2_1 _36410_ (.A(_08565_),
    .B(_08634_),
    .X(_08636_));
 sky130_fd_sc_hd__inv_2 _36411_ (.A(_08636_),
    .Y(_08637_));
 sky130_fd_sc_hd__or2_1 _36412_ (.A(_08565_),
    .B(_08634_),
    .X(_08638_));
 sky130_fd_sc_hd__and3b_2 _36413_ (.A_N(_08526_),
    .B(_08637_),
    .C(_08638_),
    .X(_08639_));
 sky130_fd_sc_hd__a21boi_4 _36414_ (.A1(_08637_),
    .A2(_08638_),
    .B1_N(_08526_),
    .Y(_08640_));
 sky130_fd_sc_hd__o221a_1 _36415_ (.A1(_05616_),
    .A2(_05619_),
    .B1(_07357_),
    .B2(_07358_),
    .C1(_07325_),
    .X(_08641_));
 sky130_fd_sc_hd__a21o_1 _36416_ (.A1(_05598_),
    .A2(_04098_),
    .B1(_04089_),
    .X(_08642_));
 sky130_fd_sc_hd__o21ai_1 _36417_ (.A1(_07343_),
    .A2(_07345_),
    .B1(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36418_ (.A(_24627_),
    .X(_08644_));
 sky130_fd_sc_hd__buf_1 _36419_ (.A(_24629_),
    .X(_08645_));
 sky130_fd_sc_hd__o21bai_1 _36420_ (.A1(_08644_),
    .A2(_08645_),
    .B1_N(_04098_),
    .Y(_08647_));
 sky130_fd_sc_hd__or3b_1 _36421_ (.A(_08644_),
    .B(_24629_),
    .C_N(_21418_),
    .X(_08648_));
 sky130_fd_sc_hd__a21o_1 _36422_ (.A1(_04089_),
    .A2(_07343_),
    .B1(_07341_),
    .X(_08649_));
 sky130_fd_sc_hd__a21oi_1 _36423_ (.A1(_08647_),
    .A2(_08648_),
    .B1(_08649_),
    .Y(_08650_));
 sky130_fd_sc_hd__and3_1 _36424_ (.A(_08649_),
    .B(_08647_),
    .C(_08648_),
    .X(_08651_));
 sky130_fd_sc_hd__buf_1 _36425_ (.A(_07329_),
    .X(_08652_));
 sky130_fd_sc_hd__nand3b_1 _36426_ (.A_N(_08652_),
    .B(_05605_),
    .C(_04094_),
    .Y(_08653_));
 sky130_fd_sc_hd__nor2_1 _36427_ (.A(_07329_),
    .B(\delay_line[21][15] ),
    .Y(_08654_));
 sky130_fd_sc_hd__and2_1 _36428_ (.A(\delay_line[21][14] ),
    .B(\delay_line[21][15] ),
    .X(_08655_));
 sky130_fd_sc_hd__buf_1 _36429_ (.A(\delay_line[21][15] ),
    .X(_08656_));
 sky130_fd_sc_hd__a2bb2o_2 _36430_ (.A1_N(_08654_),
    .A2_N(_08655_),
    .B1(_05605_),
    .B2(_08656_),
    .X(_08658_));
 sky130_fd_sc_hd__nand2_2 _36431_ (.A(_05600_),
    .B(_07329_),
    .Y(_08659_));
 sky130_fd_sc_hd__or2_1 _36432_ (.A(_08656_),
    .B(_08659_),
    .X(_08660_));
 sky130_fd_sc_hd__a21oi_1 _36433_ (.A1(_08658_),
    .A2(_08660_),
    .B1(_02550_),
    .Y(_08661_));
 sky130_fd_sc_hd__and3_1 _36434_ (.A(_08658_),
    .B(_08660_),
    .C(_02550_),
    .X(_08662_));
 sky130_fd_sc_hd__a211o_1 _36435_ (.A1(_07335_),
    .A2(_08653_),
    .B1(_08661_),
    .C1(_08662_),
    .X(_08663_));
 sky130_fd_sc_hd__o211ai_1 _36436_ (.A1(_08662_),
    .A2(_08661_),
    .B1(_08653_),
    .C1(_07335_),
    .Y(_08664_));
 sky130_fd_sc_hd__and4bb_1 _36437_ (.A_N(_08650_),
    .B_N(_08651_),
    .C(_08663_),
    .D(_08664_),
    .X(_08665_));
 sky130_fd_sc_hd__clkbuf_2 _36438_ (.A(_08665_),
    .X(_08666_));
 sky130_fd_sc_hd__a2bb2oi_1 _36439_ (.A1_N(_08650_),
    .A2_N(_08651_),
    .B1(_08663_),
    .B2(_08664_),
    .Y(_08667_));
 sky130_fd_sc_hd__a221oi_2 _36440_ (.A1(_05609_),
    .A2(_05604_),
    .B1(_07334_),
    .B2(_07335_),
    .C1(_07337_),
    .Y(_08669_));
 sky130_fd_sc_hd__o21a_1 _36441_ (.A1(_07348_),
    .A2(_08669_),
    .B1(_07353_),
    .X(_08670_));
 sky130_fd_sc_hd__o21ai_1 _36442_ (.A1(_08666_),
    .A2(_08667_),
    .B1(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__or3_1 _36443_ (.A(_08670_),
    .B(_08666_),
    .C(_08667_),
    .X(_08672_));
 sky130_fd_sc_hd__nand3_1 _36444_ (.A(_08643_),
    .B(_08671_),
    .C(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__a21o_1 _36445_ (.A1(_08671_),
    .A2(_08672_),
    .B1(_08643_),
    .X(_08674_));
 sky130_fd_sc_hd__or4bb_1 _36446_ (.A(_07359_),
    .B(_08641_),
    .C_N(_08673_),
    .D_N(_08674_),
    .X(_08675_));
 sky130_fd_sc_hd__a2bb2o_1 _36447_ (.A1_N(_07359_),
    .A2_N(_08641_),
    .B1(_08673_),
    .B2(_08674_),
    .X(_08676_));
 sky130_fd_sc_hd__o221a_1 _36448_ (.A1(_18351_),
    .A2(_07324_),
    .B1(_21410_),
    .B2(_05614_),
    .C1(_05598_),
    .X(_08677_));
 sky130_fd_sc_hd__and3_1 _36449_ (.A(_08675_),
    .B(_08676_),
    .C(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__a21oi_1 _36450_ (.A1(_08675_),
    .A2(_08676_),
    .B1(_08677_),
    .Y(_08680_));
 sky130_fd_sc_hd__nor2_1 _36451_ (.A(_08678_),
    .B(_08680_),
    .Y(_08681_));
 sky130_fd_sc_hd__o21a_1 _36452_ (.A1(_07363_),
    .A2(_07365_),
    .B1(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__a311o_1 _36453_ (.A1(_18351_),
    .A2(_05597_),
    .A3(_07364_),
    .B1(_07363_),
    .C1(_08681_),
    .X(_08683_));
 sky130_fd_sc_hd__or2b_2 _36454_ (.A(_08682_),
    .B_N(_08683_),
    .X(_08684_));
 sky130_fd_sc_hd__o21bai_4 _36455_ (.A1(_07369_),
    .A2(_07373_),
    .B1_N(_07368_),
    .Y(_08685_));
 sky130_fd_sc_hd__xor2_4 _36456_ (.A(_08684_),
    .B(_08685_),
    .X(_08686_));
 sky130_fd_sc_hd__clkbuf_2 _36457_ (.A(_07378_),
    .X(_08687_));
 sky130_fd_sc_hd__o21ai_1 _36458_ (.A1(_08687_),
    .A2(_07375_),
    .B1(_07394_),
    .Y(_08688_));
 sky130_fd_sc_hd__a21o_1 _36459_ (.A1(_07376_),
    .A2(_07378_),
    .B1(_22931_),
    .X(_08689_));
 sky130_fd_sc_hd__inv_2 _36460_ (.A(_22925_),
    .Y(_08691_));
 sky130_fd_sc_hd__or3b_1 _36461_ (.A(_08691_),
    .B(_21362_),
    .C_N(_07378_),
    .X(_08692_));
 sky130_fd_sc_hd__or2_1 _36462_ (.A(\delay_line[18][11] ),
    .B(net372),
    .X(_08693_));
 sky130_fd_sc_hd__nand2_1 _36463_ (.A(_02635_),
    .B(net372),
    .Y(_08694_));
 sky130_fd_sc_hd__clkbuf_2 _36464_ (.A(_00712_),
    .X(_08695_));
 sky130_fd_sc_hd__nand4_2 _36465_ (.A(_08693_),
    .B(_08694_),
    .C(_08695_),
    .D(_07381_),
    .Y(_08696_));
 sky130_fd_sc_hd__a22o_1 _36466_ (.A1(_00712_),
    .A2(_07381_),
    .B1(_08693_),
    .B2(_08694_),
    .X(_08697_));
 sky130_fd_sc_hd__nand4_2 _36467_ (.A(_08689_),
    .B(_08692_),
    .C(_08696_),
    .D(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__a22o_1 _36468_ (.A1(_08689_),
    .A2(_08692_),
    .B1(_08696_),
    .B2(_08697_),
    .X(_08699_));
 sky130_fd_sc_hd__nand2_1 _36469_ (.A(_07385_),
    .B(_07387_),
    .Y(_08700_));
 sky130_fd_sc_hd__a21oi_1 _36470_ (.A1(_08698_),
    .A2(_08699_),
    .B1(_08700_),
    .Y(_08702_));
 sky130_fd_sc_hd__and3_1 _36471_ (.A(_08700_),
    .B(_08698_),
    .C(_08699_),
    .X(_08703_));
 sky130_fd_sc_hd__nor2_1 _36472_ (.A(_08702_),
    .B(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__xnor2_1 _36473_ (.A(_08688_),
    .B(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__nor3_1 _36474_ (.A(_07391_),
    .B(_07392_),
    .C(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__o21ai_1 _36475_ (.A1(_07391_),
    .A2(_07392_),
    .B1(_08705_),
    .Y(_08707_));
 sky130_fd_sc_hd__or2b_1 _36476_ (.A(_08706_),
    .B_N(_08707_),
    .X(_08708_));
 sky130_fd_sc_hd__xor2_2 _36477_ (.A(_07395_),
    .B(_08708_),
    .X(_08709_));
 sky130_fd_sc_hd__a21oi_1 _36478_ (.A1(_05663_),
    .A2(_07399_),
    .B1(_07398_),
    .Y(_08710_));
 sky130_fd_sc_hd__xnor2_2 _36479_ (.A(_08709_),
    .B(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__a21boi_1 _36480_ (.A1(_05674_),
    .A2(_05672_),
    .B1_N(_05671_),
    .Y(_08713_));
 sky130_fd_sc_hd__or2b_1 _36481_ (.A(_07401_),
    .B_N(_07400_),
    .X(_08714_));
 sky130_fd_sc_hd__o21ai_2 _36482_ (.A1(_08713_),
    .A2(_07402_),
    .B1(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__xnor2_1 _36483_ (.A(_08711_),
    .B(_08715_),
    .Y(_08716_));
 sky130_fd_sc_hd__nor2_1 _36484_ (.A(_20575_),
    .B(_07406_),
    .Y(_08717_));
 sky130_fd_sc_hd__a2111o_1 _36485_ (.A1(_21376_),
    .A2(_07410_),
    .B1(_08717_),
    .C1(_07449_),
    .D1(_19400_),
    .X(_08718_));
 sky130_fd_sc_hd__buf_1 _36486_ (.A(_20561_),
    .X(_08719_));
 sky130_fd_sc_hd__o221a_1 _36487_ (.A1(_20574_),
    .A2(_08719_),
    .B1(_05680_),
    .B2(_22953_),
    .C1(_07406_),
    .X(_08720_));
 sky130_fd_sc_hd__a21boi_2 _36488_ (.A1(_07412_),
    .A2(_07441_),
    .B1_N(_07442_),
    .Y(_08721_));
 sky130_fd_sc_hd__nor2_1 _36489_ (.A(_07433_),
    .B(_07431_),
    .Y(_08722_));
 sky130_fd_sc_hd__o2bb2a_1 _36490_ (.A1_N(_07409_),
    .A2_N(_05681_),
    .B1(_07430_),
    .B2(_08722_),
    .X(_08724_));
 sky130_fd_sc_hd__a21oi_1 _36491_ (.A1(_07422_),
    .A2(_07424_),
    .B1(_07428_),
    .Y(_08725_));
 sky130_fd_sc_hd__o21ai_1 _36492_ (.A1(_24656_),
    .A2(_24657_),
    .B1(_22944_),
    .Y(_08726_));
 sky130_fd_sc_hd__or3_1 _36493_ (.A(_24657_),
    .B(_21378_),
    .C(_24656_),
    .X(_08727_));
 sky130_fd_sc_hd__a221oi_1 _36494_ (.A1(_04055_),
    .A2(_07427_),
    .B1(_08726_),
    .B2(_08727_),
    .C1(_07432_),
    .Y(_08728_));
 sky130_fd_sc_hd__inv_2 _36495_ (.A(_08728_),
    .Y(_08729_));
 sky130_fd_sc_hd__o211ai_2 _36496_ (.A1(_07431_),
    .A2(_07432_),
    .B1(_08726_),
    .C1(_08727_),
    .Y(_08730_));
 sky130_fd_sc_hd__nand2_1 _36497_ (.A(_07421_),
    .B(_24660_),
    .Y(_08731_));
 sky130_fd_sc_hd__nor2_1 _36498_ (.A(_07414_),
    .B(\delay_line[19][15] ),
    .Y(_08732_));
 sky130_fd_sc_hd__and2_1 _36499_ (.A(\delay_line[19][14] ),
    .B(\delay_line[19][15] ),
    .X(_08733_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36500_ (.A(\delay_line[19][15] ),
    .X(_08735_));
 sky130_fd_sc_hd__a2bb2o_2 _36501_ (.A1_N(_08732_),
    .A2_N(_08733_),
    .B1(_07418_),
    .B2(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__or3b_1 _36502_ (.A(_05692_),
    .B(\delay_line[19][15] ),
    .C_N(_07414_),
    .X(_08737_));
 sky130_fd_sc_hd__and3_1 _36503_ (.A(_08736_),
    .B(_08737_),
    .C(_00662_),
    .X(_08738_));
 sky130_fd_sc_hd__a21oi_1 _36504_ (.A1(_08736_),
    .A2(_08737_),
    .B1(_00662_),
    .Y(_08739_));
 sky130_fd_sc_hd__a211o_1 _36505_ (.A1(_07417_),
    .A2(_08731_),
    .B1(_08738_),
    .C1(_08739_),
    .X(_08740_));
 sky130_fd_sc_hd__clkbuf_2 _36506_ (.A(_07417_),
    .X(_08741_));
 sky130_fd_sc_hd__o211ai_2 _36507_ (.A1(_08738_),
    .A2(_08739_),
    .B1(_08741_),
    .C1(_08731_),
    .Y(_08742_));
 sky130_fd_sc_hd__and4_1 _36508_ (.A(_08729_),
    .B(_08730_),
    .C(_08740_),
    .D(_08742_),
    .X(_08743_));
 sky130_fd_sc_hd__a22oi_2 _36509_ (.A1(_08729_),
    .A2(_08730_),
    .B1(_08740_),
    .B2(_08742_),
    .Y(_08744_));
 sky130_fd_sc_hd__o221a_1 _36510_ (.A1(_07436_),
    .A2(_08725_),
    .B1(_08743_),
    .B2(_08744_),
    .C1(_07438_),
    .X(_08746_));
 sky130_fd_sc_hd__o21a_1 _36511_ (.A1(_07436_),
    .A2(_08725_),
    .B1(_07438_),
    .X(_08747_));
 sky130_fd_sc_hd__nor3_1 _36512_ (.A(_08747_),
    .B(_08743_),
    .C(_08744_),
    .Y(_08748_));
 sky130_fd_sc_hd__nor3_1 _36513_ (.A(_08724_),
    .B(_08746_),
    .C(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__o21ai_1 _36514_ (.A1(_08746_),
    .A2(_08748_),
    .B1(_08724_),
    .Y(_08750_));
 sky130_fd_sc_hd__and2b_1 _36515_ (.A_N(_08749_),
    .B(_08750_),
    .X(_08751_));
 sky130_fd_sc_hd__xnor2_1 _36516_ (.A(_08721_),
    .B(_08751_),
    .Y(_08752_));
 sky130_fd_sc_hd__xor2_1 _36517_ (.A(_08720_),
    .B(_08752_),
    .X(_08753_));
 sky130_fd_sc_hd__a21oi_1 _36518_ (.A1(_07447_),
    .A2(_08718_),
    .B1(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__and3_1 _36519_ (.A(_07447_),
    .B(_08718_),
    .C(_08753_),
    .X(_08755_));
 sky130_fd_sc_hd__nor2_1 _36520_ (.A(_08754_),
    .B(_08755_),
    .Y(_08757_));
 sky130_fd_sc_hd__o21a_1 _36521_ (.A1(_07453_),
    .A2(_07456_),
    .B1(_08757_),
    .X(_08758_));
 sky130_fd_sc_hd__or3_1 _36522_ (.A(_07453_),
    .B(_07456_),
    .C(_08757_),
    .X(_08759_));
 sky130_fd_sc_hd__or3b_4 _36523_ (.A(_08716_),
    .B(_08758_),
    .C_N(_08759_),
    .X(_08760_));
 sky130_fd_sc_hd__inv_2 _36524_ (.A(_08758_),
    .Y(_08761_));
 sky130_fd_sc_hd__a21bo_1 _36525_ (.A1(_08759_),
    .A2(_08761_),
    .B1_N(_08716_),
    .X(_08762_));
 sky130_fd_sc_hd__and2_2 _36526_ (.A(_08760_),
    .B(_08762_),
    .X(_08763_));
 sky130_fd_sc_hd__xor2_4 _36527_ (.A(_08686_),
    .B(_08763_),
    .X(_08764_));
 sky130_fd_sc_hd__o21a_1 _36528_ (.A1(_08639_),
    .A2(_08640_),
    .B1(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__nor3_1 _36529_ (.A(_08640_),
    .B(_08764_),
    .C(_08639_),
    .Y(_08766_));
 sky130_fd_sc_hd__a21o_1 _36530_ (.A1(_07318_),
    .A2(_07319_),
    .B1(_07462_),
    .X(_08768_));
 sky130_fd_sc_hd__o21a_1 _36531_ (.A1(_07318_),
    .A2(_07319_),
    .B1(_08768_),
    .X(_08769_));
 sky130_fd_sc_hd__o21ai_1 _36532_ (.A1(_08765_),
    .A2(_08766_),
    .B1(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__or3_4 _36533_ (.A(_08769_),
    .B(_08765_),
    .C(_08766_),
    .X(_08771_));
 sky130_fd_sc_hd__nand2_4 _36534_ (.A(_08770_),
    .B(_08771_),
    .Y(_08772_));
 sky130_fd_sc_hd__xor2_1 _36535_ (.A(_08524_),
    .B(_08772_),
    .X(_08773_));
 sky130_fd_sc_hd__nor2_1 _36536_ (.A(_08396_),
    .B(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__nand2_1 _36537_ (.A(_08773_),
    .B(_08396_),
    .Y(_08775_));
 sky130_fd_sc_hd__and2b_1 _36538_ (.A_N(_08774_),
    .B(_08775_),
    .X(_08776_));
 sky130_fd_sc_hd__o21ai_4 _36539_ (.A1(_06988_),
    .A2(_07065_),
    .B1(_07067_),
    .Y(_08777_));
 sky130_fd_sc_hd__a21o_1 _36540_ (.A1(_05725_),
    .A2(_05729_),
    .B1(_07196_),
    .X(_08779_));
 sky130_fd_sc_hd__or2_1 _36541_ (.A(_07033_),
    .B(_07060_),
    .X(_08780_));
 sky130_fd_sc_hd__o21a_1 _36542_ (.A1(_05576_),
    .A2(_05581_),
    .B1(_07010_),
    .X(_08781_));
 sky130_fd_sc_hd__o211ai_2 _36543_ (.A1(_05569_),
    .A2(_05571_),
    .B1(_07003_),
    .C1(_07004_),
    .Y(_08782_));
 sky130_fd_sc_hd__a21o_1 _36544_ (.A1(_06989_),
    .A2(_06995_),
    .B1(_04267_),
    .X(_08783_));
 sky130_fd_sc_hd__clkbuf_2 _36545_ (.A(_06989_),
    .X(_08784_));
 sky130_fd_sc_hd__nand3_2 _36546_ (.A(_04267_),
    .B(_08784_),
    .C(_06995_),
    .Y(_08785_));
 sky130_fd_sc_hd__a31o_1 _36547_ (.A1(_06999_),
    .A2(_06989_),
    .A3(_06992_),
    .B1(_06998_),
    .X(_08786_));
 sky130_fd_sc_hd__a21oi_1 _36548_ (.A1(_08783_),
    .A2(_08785_),
    .B1(_08786_),
    .Y(_08787_));
 sky130_fd_sc_hd__and3_1 _36549_ (.A(_08783_),
    .B(_08785_),
    .C(_08786_),
    .X(_08788_));
 sky130_fd_sc_hd__nor3_1 _36550_ (.A(_08787_),
    .B(_01028_),
    .C(_08788_),
    .Y(_08790_));
 sky130_fd_sc_hd__o21a_1 _36551_ (.A1(_08788_),
    .A2(_08787_),
    .B1(_01028_),
    .X(_08791_));
 sky130_fd_sc_hd__o211a_1 _36552_ (.A1(_08790_),
    .A2(_08791_),
    .B1(_07001_),
    .C1(_07004_),
    .X(_08792_));
 sky130_fd_sc_hd__a211o_1 _36553_ (.A1(_07001_),
    .A2(_07004_),
    .B1(_08790_),
    .C1(_08791_),
    .X(_08793_));
 sky130_fd_sc_hd__or2b_1 _36554_ (.A(_08792_),
    .B_N(_08793_),
    .X(_08794_));
 sky130_fd_sc_hd__xor2_1 _36555_ (.A(_08782_),
    .B(_08794_),
    .X(_08795_));
 sky130_fd_sc_hd__or3_1 _36556_ (.A(net167),
    .B(_08781_),
    .C(_08795_),
    .X(_08796_));
 sky130_fd_sc_hd__o21ai_1 _36557_ (.A1(net167),
    .A2(_08781_),
    .B1(_08795_),
    .Y(_08797_));
 sky130_fd_sc_hd__nand2_2 _36558_ (.A(_08796_),
    .B(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__inv_2 _36559_ (.A(_07028_),
    .Y(_08799_));
 sky130_fd_sc_hd__nand2_1 _36560_ (.A(_07032_),
    .B(_07031_),
    .Y(_08801_));
 sky130_fd_sc_hd__clkbuf_2 _36561_ (.A(\delay_line[26][15] ),
    .X(_08802_));
 sky130_fd_sc_hd__inv_2 _36562_ (.A(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__nand2_1 _36563_ (.A(_24337_),
    .B(_00994_),
    .Y(_08804_));
 sky130_fd_sc_hd__nor2_1 _36564_ (.A(_00994_),
    .B(\delay_line[26][11] ),
    .Y(_08805_));
 sky130_fd_sc_hd__and2_1 _36565_ (.A(_00994_),
    .B(\delay_line[26][11] ),
    .X(_08806_));
 sky130_fd_sc_hd__or3b_2 _36566_ (.A(_08805_),
    .B(_08806_),
    .C_N(_21228_),
    .X(_08807_));
 sky130_fd_sc_hd__o21bai_1 _36567_ (.A1(_08805_),
    .A2(_08806_),
    .B1_N(_21228_),
    .Y(_08808_));
 sky130_fd_sc_hd__nand2_1 _36568_ (.A(_08807_),
    .B(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__a21oi_2 _36569_ (.A1(_08804_),
    .A2(_07018_),
    .B1(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__and3_1 _36570_ (.A(_08804_),
    .B(_07018_),
    .C(_08809_),
    .X(_08812_));
 sky130_fd_sc_hd__nor2_1 _36571_ (.A(_08810_),
    .B(_08812_),
    .Y(_08813_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36572_ (.A(_07022_),
    .X(_08814_));
 sky130_fd_sc_hd__a21oi_1 _36573_ (.A1(_05538_),
    .A2(_07024_),
    .B1(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__xor2_1 _36574_ (.A(_08813_),
    .B(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__xor2_1 _36575_ (.A(_08803_),
    .B(_08816_),
    .X(_08817_));
 sky130_fd_sc_hd__or3b_1 _36576_ (.A(_05538_),
    .B(_05539_),
    .C_N(_04298_),
    .X(_08818_));
 sky130_fd_sc_hd__o32a_1 _36577_ (.A1(_08814_),
    .A2(_07023_),
    .A3(_08818_),
    .B1(_07015_),
    .B2(_07026_),
    .X(_08819_));
 sky130_fd_sc_hd__and2b_1 _36578_ (.A_N(_08817_),
    .B(_08819_),
    .X(_08820_));
 sky130_fd_sc_hd__and2b_1 _36579_ (.A_N(_08819_),
    .B(_08817_),
    .X(_08821_));
 sky130_fd_sc_hd__or2_1 _36580_ (.A(_08820_),
    .B(_08821_),
    .X(_08823_));
 sky130_fd_sc_hd__and3_1 _36581_ (.A(_08799_),
    .B(_08801_),
    .C(_08823_),
    .X(_08824_));
 sky130_fd_sc_hd__a21oi_2 _36582_ (.A1(_08799_),
    .A2(_08801_),
    .B1(_08823_),
    .Y(_08825_));
 sky130_fd_sc_hd__o31a_1 _36583_ (.A1(_02223_),
    .A2(_05508_),
    .A3(_07035_),
    .B1(_05501_),
    .X(_08826_));
 sky130_fd_sc_hd__or3_1 _36584_ (.A(net329),
    .B(_05496_),
    .C(_04315_),
    .X(_08827_));
 sky130_fd_sc_hd__o2bb2a_1 _36585_ (.A1_N(_08826_),
    .A2_N(_08827_),
    .B1(_07034_),
    .B2(_05501_),
    .X(_08828_));
 sky130_fd_sc_hd__or2_1 _36586_ (.A(_24365_),
    .B(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__nand2_1 _36587_ (.A(_24365_),
    .B(_08828_),
    .Y(_08830_));
 sky130_fd_sc_hd__a2bb2o_1 _36588_ (.A1_N(_23157_),
    .A2_N(_07042_),
    .B1(_05497_),
    .B2(_07040_),
    .X(_08831_));
 sky130_fd_sc_hd__a21oi_1 _36589_ (.A1(_08829_),
    .A2(_08830_),
    .B1(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__nand3_1 _36590_ (.A(_08831_),
    .B(_08829_),
    .C(_08830_),
    .Y(_08834_));
 sky130_fd_sc_hd__inv_2 _36591_ (.A(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__nor3_1 _36592_ (.A(_23162_),
    .B(_08832_),
    .C(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__o32a_1 _36593_ (.A1(_21238_),
    .A2(_23152_),
    .A3(_23155_),
    .B1(_08832_),
    .B2(_08835_),
    .X(_08837_));
 sky130_fd_sc_hd__nor2_1 _36594_ (.A(_08836_),
    .B(_08837_),
    .Y(_08838_));
 sky130_fd_sc_hd__o21a_1 _36595_ (.A1(_07048_),
    .A2(_07049_),
    .B1(_08838_),
    .X(_08839_));
 sky130_fd_sc_hd__o221a_1 _36596_ (.A1(_05505_),
    .A2(_07046_),
    .B1(_08836_),
    .B2(_08837_),
    .C1(_07047_),
    .X(_08840_));
 sky130_fd_sc_hd__nor2_1 _36597_ (.A(_08839_),
    .B(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__and2_1 _36598_ (.A(_07055_),
    .B(_08841_),
    .X(_08842_));
 sky130_fd_sc_hd__nor2_1 _36599_ (.A(_07055_),
    .B(_08841_),
    .Y(_08843_));
 sky130_fd_sc_hd__nor2_1 _36600_ (.A(_08842_),
    .B(_08843_),
    .Y(_08845_));
 sky130_fd_sc_hd__o21bai_2 _36601_ (.A1(_07057_),
    .A2(_07059_),
    .B1_N(net128),
    .Y(_08846_));
 sky130_fd_sc_hd__or2_1 _36602_ (.A(_08845_),
    .B(_08846_),
    .X(_08847_));
 sky130_fd_sc_hd__nand2_1 _36603_ (.A(_08846_),
    .B(_08845_),
    .Y(_08848_));
 sky130_fd_sc_hd__a2bb2oi_1 _36604_ (.A1_N(_08824_),
    .A2_N(_08825_),
    .B1(_08847_),
    .B2(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__or4bb_1 _36605_ (.A(_08824_),
    .B(_08825_),
    .C_N(_08847_),
    .D_N(_08848_),
    .X(_08850_));
 sky130_fd_sc_hd__inv_2 _36606_ (.A(_08850_),
    .Y(_08851_));
 sky130_fd_sc_hd__nor3_1 _36607_ (.A(_08798_),
    .B(_08849_),
    .C(_08851_),
    .Y(_08852_));
 sky130_fd_sc_hd__o21a_1 _36608_ (.A1(_08851_),
    .A2(_08849_),
    .B1(_08798_),
    .X(_08853_));
 sky130_fd_sc_hd__a211oi_1 _36609_ (.A1(_08780_),
    .A2(_07064_),
    .B1(_08852_),
    .C1(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__o221a_1 _36610_ (.A1(_07033_),
    .A2(_07060_),
    .B1(_08852_),
    .B2(_08853_),
    .C1(_07064_),
    .X(_08856_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36611_ (.A(_05415_),
    .X(_08857_));
 sky130_fd_sc_hd__buf_1 _36612_ (.A(\delay_line[31][15] ),
    .X(_08858_));
 sky130_fd_sc_hd__and2b_1 _36613_ (.A_N(_05409_),
    .B(_04351_),
    .X(_08859_));
 sky130_fd_sc_hd__o21ai_1 _36614_ (.A1(_08858_),
    .A2(_08859_),
    .B1(_05415_),
    .Y(_08860_));
 sky130_fd_sc_hd__o31a_1 _36615_ (.A1(_08857_),
    .A2(_08858_),
    .A3(_05413_),
    .B1(_08860_),
    .X(_08861_));
 sky130_fd_sc_hd__or2_1 _36616_ (.A(_00884_),
    .B(_05423_),
    .X(_08862_));
 sky130_fd_sc_hd__nor2_1 _36617_ (.A(_20313_),
    .B(_06957_),
    .Y(_08863_));
 sky130_fd_sc_hd__buf_1 _36618_ (.A(_00884_),
    .X(_08864_));
 sky130_fd_sc_hd__nand2_1 _36619_ (.A(_05423_),
    .B(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__and3_1 _36620_ (.A(_08862_),
    .B(_08863_),
    .C(_08865_),
    .X(_08867_));
 sky130_fd_sc_hd__a22o_1 _36621_ (.A1(_23213_),
    .A2(_23212_),
    .B1(_08862_),
    .B2(_08865_),
    .X(_08868_));
 sky130_fd_sc_hd__inv_2 _36622_ (.A(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__nor3_1 _36623_ (.A(_08861_),
    .B(_08867_),
    .C(_08869_),
    .Y(_08870_));
 sky130_fd_sc_hd__o21a_1 _36624_ (.A1(_08867_),
    .A2(_08869_),
    .B1(_08861_),
    .X(_08871_));
 sky130_fd_sc_hd__a211o_1 _36625_ (.A1(_05419_),
    .A2(_06965_),
    .B1(_06960_),
    .C1(_06961_),
    .X(_08872_));
 sky130_fd_sc_hd__o221ai_2 _36626_ (.A1(_05419_),
    .A2(_06965_),
    .B1(net224),
    .B2(_08871_),
    .C1(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__a211o_1 _36627_ (.A1(_06966_),
    .A2(_08872_),
    .B1(net224),
    .C1(_08871_),
    .X(_08874_));
 sky130_fd_sc_hd__nand2_1 _36628_ (.A(_08873_),
    .B(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__xor2_1 _36629_ (.A(_06960_),
    .B(_08875_),
    .X(_08876_));
 sky130_fd_sc_hd__a21oi_2 _36630_ (.A1(_06972_),
    .A2(_06973_),
    .B1(_08876_),
    .Y(_08878_));
 sky130_fd_sc_hd__and3_1 _36631_ (.A(_06972_),
    .B(_06973_),
    .C(_08876_),
    .X(_08879_));
 sky130_fd_sc_hd__or2_1 _36632_ (.A(_08878_),
    .B(_08879_),
    .X(_08880_));
 sky130_fd_sc_hd__nor2_1 _36633_ (.A(_06978_),
    .B(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__and2_1 _36634_ (.A(_06978_),
    .B(_08880_),
    .X(_08882_));
 sky130_fd_sc_hd__or2_2 _36635_ (.A(_08881_),
    .B(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__a22oi_4 _36636_ (.A1(_06981_),
    .A2(_06979_),
    .B1(_06955_),
    .B2(_06980_),
    .Y(_08884_));
 sky130_fd_sc_hd__xor2_4 _36637_ (.A(_08883_),
    .B(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__and2b_1 _36638_ (.A_N(\delay_line[29][10] ),
    .B(\delay_line[29][14] ),
    .X(_08886_));
 sky130_fd_sc_hd__and2b_1 _36639_ (.A_N(\delay_line[29][14] ),
    .B(\delay_line[29][10] ),
    .X(_08887_));
 sky130_fd_sc_hd__or2_2 _36640_ (.A(_08886_),
    .B(_08887_),
    .X(_08889_));
 sky130_fd_sc_hd__a21bo_1 _36641_ (.A1(_05445_),
    .A2(_06944_),
    .B1_N(_06943_),
    .X(_08890_));
 sky130_fd_sc_hd__xnor2_4 _36642_ (.A(_08889_),
    .B(_08890_),
    .Y(_08891_));
 sky130_fd_sc_hd__a31o_2 _36643_ (.A1(_04408_),
    .A2(_05448_),
    .A3(_06945_),
    .B1(_06950_),
    .X(_08892_));
 sky130_fd_sc_hd__xnor2_4 _36644_ (.A(_08891_),
    .B(_08892_),
    .Y(_08893_));
 sky130_fd_sc_hd__nand4_1 _36645_ (.A(_06919_),
    .B(_06913_),
    .C(_06916_),
    .D(_06917_),
    .Y(_08894_));
 sky130_fd_sc_hd__buf_1 _36646_ (.A(_00932_),
    .X(_08895_));
 sky130_fd_sc_hd__inv_2 _36647_ (.A(_05457_),
    .Y(_08896_));
 sky130_fd_sc_hd__nor2_1 _36648_ (.A(_08895_),
    .B(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__nor2_1 _36649_ (.A(_02110_),
    .B(_05457_),
    .Y(_08898_));
 sky130_fd_sc_hd__o21ai_1 _36650_ (.A1(_08897_),
    .A2(_08898_),
    .B1(_06911_),
    .Y(_08900_));
 sky130_fd_sc_hd__or3_1 _36651_ (.A(_06911_),
    .B(_08897_),
    .C(_08898_),
    .X(_08901_));
 sky130_fd_sc_hd__buf_1 _36652_ (.A(_04383_),
    .X(_08902_));
 sky130_fd_sc_hd__a21boi_1 _36653_ (.A1(_06924_),
    .A2(_08902_),
    .B1_N(_04384_),
    .Y(_08903_));
 sky130_fd_sc_hd__or3b_1 _36654_ (.A(_04384_),
    .B(_02101_),
    .C_N(_06924_),
    .X(_08904_));
 sky130_fd_sc_hd__and4bb_1 _36655_ (.A_N(_02089_),
    .B_N(_08903_),
    .C(_08904_),
    .D(_05476_),
    .X(_08905_));
 sky130_fd_sc_hd__and3_1 _36656_ (.A(_04399_),
    .B(_06924_),
    .C(_04383_),
    .X(_08906_));
 sky130_fd_sc_hd__o2bb2a_1 _36657_ (.A1_N(_05476_),
    .A2_N(_20339_),
    .B1(_08906_),
    .B2(_08903_),
    .X(_08907_));
 sky130_fd_sc_hd__a211oi_2 _36658_ (.A1(_08900_),
    .A2(_08901_),
    .B1(_08905_),
    .C1(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__o211a_1 _36659_ (.A1(_08905_),
    .A2(_08907_),
    .B1(_08900_),
    .C1(_08901_),
    .X(_08909_));
 sky130_fd_sc_hd__a211o_1 _36660_ (.A1(_06919_),
    .A2(_08894_),
    .B1(_08908_),
    .C1(_08909_),
    .X(_08911_));
 sky130_fd_sc_hd__o211ai_1 _36661_ (.A1(_08908_),
    .A2(_08909_),
    .B1(_06919_),
    .C1(_08894_),
    .Y(_08912_));
 sky130_fd_sc_hd__and2b_1 _36662_ (.A_N(_06914_),
    .B(_06916_),
    .X(_08913_));
 sky130_fd_sc_hd__and3_1 _36663_ (.A(_08911_),
    .B(_08912_),
    .C(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__a21oi_1 _36664_ (.A1(_08911_),
    .A2(_08912_),
    .B1(_08913_),
    .Y(_08915_));
 sky130_fd_sc_hd__or2_1 _36665_ (.A(_08914_),
    .B(_08915_),
    .X(_08916_));
 sky130_fd_sc_hd__or3_1 _36666_ (.A(_06922_),
    .B(_06928_),
    .C(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__o21ai_1 _36667_ (.A1(_06922_),
    .A2(_06928_),
    .B1(_08916_),
    .Y(_08918_));
 sky130_fd_sc_hd__nand2_1 _36668_ (.A(_08917_),
    .B(_08918_),
    .Y(_08919_));
 sky130_fd_sc_hd__nor2_1 _36669_ (.A(_06932_),
    .B(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__and2_1 _36670_ (.A(_06932_),
    .B(_08919_),
    .X(_08922_));
 sky130_fd_sc_hd__nor2_2 _36671_ (.A(_08920_),
    .B(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__a21oi_1 _36672_ (.A1(_05484_),
    .A2(_05483_),
    .B1(_06933_),
    .Y(_08924_));
 sky130_fd_sc_hd__o22ai_4 _36673_ (.A1(_05479_),
    .A2(_08924_),
    .B1(_06934_),
    .B2(_06936_),
    .Y(_08925_));
 sky130_fd_sc_hd__xor2_4 _36674_ (.A(_08923_),
    .B(_08925_),
    .X(_08926_));
 sky130_fd_sc_hd__xnor2_4 _36675_ (.A(_08893_),
    .B(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__xnor2_4 _36676_ (.A(_08885_),
    .B(_08927_),
    .Y(_08928_));
 sky130_fd_sc_hd__o21ai_1 _36677_ (.A1(_08854_),
    .A2(_08856_),
    .B1(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__or3_1 _36678_ (.A(_08854_),
    .B(_08856_),
    .C(_08928_),
    .X(_08930_));
 sky130_fd_sc_hd__nand2_2 _36679_ (.A(_08929_),
    .B(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__a21oi_1 _36680_ (.A1(_08779_),
    .A2(_07201_),
    .B1(_08931_),
    .Y(_08933_));
 sky130_fd_sc_hd__and3_1 _36681_ (.A(_08779_),
    .B(_07201_),
    .C(_08931_),
    .X(_08934_));
 sky130_fd_sc_hd__nor2_1 _36682_ (.A(_08933_),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__xor2_1 _36683_ (.A(_08777_),
    .B(_08935_),
    .X(_08936_));
 sky130_fd_sc_hd__inv_2 _36684_ (.A(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__xnor2_1 _36685_ (.A(_08776_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__xnor2_1 _36686_ (.A(_08395_),
    .B(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__a21o_1 _36687_ (.A1(_08392_),
    .A2(_08394_),
    .B1(_08939_),
    .X(_08940_));
 sky130_fd_sc_hd__nand3_2 _36688_ (.A(_08392_),
    .B(_08394_),
    .C(_08939_),
    .Y(_08941_));
 sky130_fd_sc_hd__nand2_2 _36689_ (.A(_08940_),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__xor2_2 _36690_ (.A(_08190_),
    .B(_08942_),
    .X(_08944_));
 sky130_fd_sc_hd__nand2_2 _36691_ (.A(_08189_),
    .B(_08944_),
    .Y(_08945_));
 sky130_fd_sc_hd__and3_1 _36692_ (.A(_08185_),
    .B(_08174_),
    .C(_08180_),
    .X(_08946_));
 sky130_fd_sc_hd__o21bai_1 _36693_ (.A1(_08187_),
    .A2(_08946_),
    .B1_N(_08944_),
    .Y(_08947_));
 sky130_fd_sc_hd__o21a_1 _36694_ (.A1(_08188_),
    .A2(_08945_),
    .B1(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__o21ai_2 _36695_ (.A1(_07487_),
    .A2(_07484_),
    .B1(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__clkbuf_2 _36696_ (.A(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__nor2_1 _36697_ (.A(_08188_),
    .B(_08945_),
    .Y(_08951_));
 sky130_fd_sc_hd__a21o_1 _36698_ (.A1(_08175_),
    .A2(_08181_),
    .B1(_08186_),
    .X(_08952_));
 sky130_fd_sc_hd__a21oi_2 _36699_ (.A1(_08952_),
    .A2(_08189_),
    .B1(_08944_),
    .Y(_08953_));
 sky130_fd_sc_hd__o211ai_4 _36700_ (.A1(_08951_),
    .A2(_08953_),
    .B1(_07486_),
    .C1(_07586_),
    .Y(_08955_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36701_ (.A(_07497_),
    .X(_08956_));
 sky130_fd_sc_hd__buf_1 _36702_ (.A(_08956_),
    .X(_08957_));
 sky130_fd_sc_hd__nand2_2 _36703_ (.A(_23569_),
    .B(_01422_),
    .Y(_08958_));
 sky130_fd_sc_hd__buf_1 _36704_ (.A(_07507_),
    .X(_08959_));
 sky130_fd_sc_hd__and2b_2 _36705_ (.A_N(_08959_),
    .B(_08956_),
    .X(_08960_));
 sky130_fd_sc_hd__buf_2 _36706_ (.A(_07509_),
    .X(_08961_));
 sky130_fd_sc_hd__nor2_1 _36707_ (.A(_07508_),
    .B(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__a211oi_2 _36708_ (.A1(_08958_),
    .A2(_08962_),
    .B1(_07510_),
    .C1(_08960_),
    .Y(_08963_));
 sky130_fd_sc_hd__a221o_2 _36709_ (.A1(_07502_),
    .A2(_08957_),
    .B1(_08958_),
    .B2(_08960_),
    .C1(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__buf_1 _36710_ (.A(_08959_),
    .X(_08966_));
 sky130_fd_sc_hd__buf_2 _36711_ (.A(_08966_),
    .X(_08967_));
 sky130_fd_sc_hd__and3b_1 _36712_ (.A_N(_08967_),
    .B(_08958_),
    .C(_08956_),
    .X(_08968_));
 sky130_fd_sc_hd__clkbuf_4 _36713_ (.A(_04552_),
    .X(_08969_));
 sky130_fd_sc_hd__o21ai_4 _36714_ (.A1(_08968_),
    .A2(_08963_),
    .B1(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__nor2_1 _36715_ (.A(_03011_),
    .B(_23691_),
    .Y(_08971_));
 sky130_fd_sc_hd__and2_1 _36716_ (.A(_23691_),
    .B(_03011_),
    .X(_08972_));
 sky130_fd_sc_hd__buf_1 _36717_ (.A(_01444_),
    .X(_08973_));
 sky130_fd_sc_hd__o21a_1 _36718_ (.A1(_08973_),
    .A2(_07539_),
    .B1(_01443_),
    .X(_08974_));
 sky130_fd_sc_hd__buf_1 _36719_ (.A(_03037_),
    .X(_08975_));
 sky130_fd_sc_hd__o21ba_2 _36720_ (.A1(_03033_),
    .A2(_08974_),
    .B1_N(_08975_),
    .X(_08977_));
 sky130_fd_sc_hd__clkbuf_2 _36721_ (.A(_07539_),
    .X(_08978_));
 sky130_fd_sc_hd__a21o_1 _36722_ (.A1(_08973_),
    .A2(_08978_),
    .B1(_08974_),
    .X(_08979_));
 sky130_fd_sc_hd__and2b_1 _36723_ (.A_N(_08979_),
    .B(_08975_),
    .X(_08980_));
 sky130_fd_sc_hd__or3_1 _36724_ (.A(_03012_),
    .B(_08977_),
    .C(_08980_),
    .X(_08981_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36725_ (.A(_03012_),
    .X(_08982_));
 sky130_fd_sc_hd__o21ai_1 _36726_ (.A1(_08977_),
    .A2(_08980_),
    .B1(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__nor3_1 _36727_ (.A(_07520_),
    .B(_07517_),
    .C(_07518_),
    .Y(_08984_));
 sky130_fd_sc_hd__a211oi_1 _36728_ (.A1(_08981_),
    .A2(_08983_),
    .B1(_07517_),
    .C1(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__o211a_1 _36729_ (.A1(_07517_),
    .A2(_08984_),
    .B1(_08981_),
    .C1(_08983_),
    .X(_08986_));
 sky130_fd_sc_hd__o22a_1 _36730_ (.A1(_08971_),
    .A2(_08972_),
    .B1(_08985_),
    .B2(_08986_),
    .X(_08988_));
 sky130_fd_sc_hd__nor4_1 _36731_ (.A(_08971_),
    .B(_08972_),
    .C(_08985_),
    .D(_08986_),
    .Y(_08989_));
 sky130_fd_sc_hd__o221a_2 _36732_ (.A1(_07523_),
    .A2(_07515_),
    .B1(_08988_),
    .B2(_08989_),
    .C1(_07524_),
    .X(_08990_));
 sky130_fd_sc_hd__o21a_1 _36733_ (.A1(_07515_),
    .A2(_07523_),
    .B1(_07524_),
    .X(_08991_));
 sky130_fd_sc_hd__or2_1 _36734_ (.A(_08989_),
    .B(_08988_),
    .X(_08992_));
 sky130_fd_sc_hd__nor2_2 _36735_ (.A(_08991_),
    .B(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__a211oi_4 _36736_ (.A1(_08964_),
    .A2(_08970_),
    .B1(_08990_),
    .C1(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__a21bo_1 _36737_ (.A1(_07534_),
    .A2(_07557_),
    .B1_N(_07556_),
    .X(_08995_));
 sky130_fd_sc_hd__nor4_1 _36738_ (.A(_00435_),
    .B(_07546_),
    .C(_05133_),
    .D(_07551_),
    .Y(_08996_));
 sky130_fd_sc_hd__or2_1 _36739_ (.A(_06650_),
    .B(_06652_),
    .X(_08997_));
 sky130_fd_sc_hd__buf_1 _36740_ (.A(\delay_line[20][15] ),
    .X(_08999_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36741_ (.A(_04529_),
    .X(_09000_));
 sky130_fd_sc_hd__o21ba_1 _36742_ (.A1(_04528_),
    .A2(_09000_),
    .B1_N(_08973_),
    .X(_09001_));
 sky130_fd_sc_hd__o21ai_4 _36743_ (.A1(_04526_),
    .A2(_04525_),
    .B1(_03030_),
    .Y(_09002_));
 sky130_fd_sc_hd__a21oi_1 _36744_ (.A1(_07539_),
    .A2(_07540_),
    .B1(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__clkbuf_2 _36745_ (.A(_09003_),
    .X(_09004_));
 sky130_fd_sc_hd__o2bb2a_1 _36746_ (.A1_N(_07540_),
    .A2_N(_08999_),
    .B1(_09001_),
    .B2(_09004_),
    .X(_09005_));
 sky130_fd_sc_hd__buf_2 _36747_ (.A(_07540_),
    .X(_09006_));
 sky130_fd_sc_hd__nor2_1 _36748_ (.A(_09001_),
    .B(_09003_),
    .Y(_09007_));
 sky130_fd_sc_hd__and3_1 _36749_ (.A(_09006_),
    .B(_08999_),
    .C(_09007_),
    .X(_09008_));
 sky130_fd_sc_hd__or4_1 _36750_ (.A(_06633_),
    .B(_09005_),
    .C(_06635_),
    .D(_09008_),
    .X(_09010_));
 sky130_fd_sc_hd__o22ai_2 _36751_ (.A1(_06635_),
    .A2(_06633_),
    .B1(_09005_),
    .B2(_09008_),
    .Y(_09011_));
 sky130_fd_sc_hd__clkbuf_4 _36752_ (.A(_07538_),
    .X(_09012_));
 sky130_fd_sc_hd__a211oi_2 _36753_ (.A1(_09010_),
    .A2(_09011_),
    .B1(_09012_),
    .C1(_07551_),
    .Y(_09013_));
 sky130_fd_sc_hd__o211a_1 _36754_ (.A1(_09012_),
    .A2(_07551_),
    .B1(_09010_),
    .C1(_09011_),
    .X(_09014_));
 sky130_fd_sc_hd__a211o_1 _36755_ (.A1(_06642_),
    .A2(_08997_),
    .B1(_09013_),
    .C1(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__o221ai_2 _36756_ (.A1(_06650_),
    .A2(_06652_),
    .B1(_09013_),
    .B2(_09014_),
    .C1(_06643_),
    .Y(_09016_));
 sky130_fd_sc_hd__o211a_1 _36757_ (.A1(net197),
    .A2(_07554_),
    .B1(_09015_),
    .C1(_09016_),
    .X(_09017_));
 sky130_fd_sc_hd__a211oi_1 _36758_ (.A1(_09015_),
    .A2(_09016_),
    .B1(net197),
    .C1(_07554_),
    .Y(_09018_));
 sky130_fd_sc_hd__nor2_1 _36759_ (.A(_09017_),
    .B(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__xnor2_1 _36760_ (.A(_08995_),
    .B(_09019_),
    .Y(_09021_));
 sky130_fd_sc_hd__o211ai_4 _36761_ (.A1(_08990_),
    .A2(_08993_),
    .B1(_08964_),
    .C1(_08970_),
    .Y(_09022_));
 sky130_fd_sc_hd__inv_2 _36762_ (.A(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__nor3_2 _36763_ (.A(_08994_),
    .B(_09021_),
    .C(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__o21a_1 _36764_ (.A1(_09023_),
    .A2(_08994_),
    .B1(_09021_),
    .X(_09025_));
 sky130_fd_sc_hd__o21ai_1 _36765_ (.A1(_07491_),
    .A2(_07489_),
    .B1(_06662_),
    .Y(_09026_));
 sky130_fd_sc_hd__o211ai_4 _36766_ (.A1(_09024_),
    .A2(_09025_),
    .B1(_06659_),
    .C1(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__a21oi_1 _36767_ (.A1(_06660_),
    .A2(_06661_),
    .B1(_06077_),
    .Y(_09028_));
 sky130_fd_sc_hd__nor2_1 _36768_ (.A(_09024_),
    .B(_09025_),
    .Y(_09029_));
 sky130_fd_sc_hd__o21ai_2 _36769_ (.A1(_09028_),
    .A2(_06664_),
    .B1(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__nand2_1 _36770_ (.A(_09027_),
    .B(_09030_),
    .Y(_09032_));
 sky130_fd_sc_hd__nor2_1 _36771_ (.A(_07563_),
    .B(_07571_),
    .Y(_09033_));
 sky130_fd_sc_hd__nand2_1 _36772_ (.A(_09032_),
    .B(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__o211ai_2 _36773_ (.A1(_07563_),
    .A2(_07571_),
    .B1(_09027_),
    .C1(_09030_),
    .Y(_09035_));
 sky130_fd_sc_hd__nand4_1 _36774_ (.A(_08950_),
    .B(_08955_),
    .C(_09034_),
    .D(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__o21ai_1 _36775_ (.A1(_08188_),
    .A2(_08945_),
    .B1(_08947_),
    .Y(_09037_));
 sky130_fd_sc_hd__a21oi_1 _36776_ (.A1(_07486_),
    .A2(_07586_),
    .B1(_09037_),
    .Y(_09038_));
 sky130_fd_sc_hd__o211a_2 _36777_ (.A1(_08951_),
    .A2(_08953_),
    .B1(_07486_),
    .C1(_07586_),
    .X(_09039_));
 sky130_fd_sc_hd__nand2_1 _36778_ (.A(_09034_),
    .B(_09035_),
    .Y(_09040_));
 sky130_fd_sc_hd__o21ai_1 _36779_ (.A1(_09038_),
    .A2(_09039_),
    .B1(_09040_),
    .Y(_09041_));
 sky130_fd_sc_hd__nand3_1 _36780_ (.A(_07642_),
    .B(_09036_),
    .C(_09041_),
    .Y(_09043_));
 sky130_fd_sc_hd__a21oi_2 _36781_ (.A1(_07584_),
    .A2(_07578_),
    .B1(_07587_),
    .Y(_09044_));
 sky130_fd_sc_hd__clkbuf_2 _36782_ (.A(_09030_),
    .X(_09045_));
 sky130_fd_sc_hd__a21boi_2 _36783_ (.A1(_09027_),
    .A2(_09045_),
    .B1_N(_09033_),
    .Y(_09046_));
 sky130_fd_sc_hd__o211a_1 _36784_ (.A1(_07563_),
    .A2(_07571_),
    .B1(_09027_),
    .C1(_09030_),
    .X(_09047_));
 sky130_fd_sc_hd__nor2_1 _36785_ (.A(_09046_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__o21ai_2 _36786_ (.A1(_09038_),
    .A2(_09039_),
    .B1(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__o211ai_4 _36787_ (.A1(_09046_),
    .A2(_09047_),
    .B1(_08949_),
    .C1(_08955_),
    .Y(_09050_));
 sky130_fd_sc_hd__nand3_1 _36788_ (.A(_09044_),
    .B(_09049_),
    .C(_09050_),
    .Y(_09051_));
 sky130_fd_sc_hd__and2_1 _36789_ (.A(_07611_),
    .B(_07612_),
    .X(_09052_));
 sky130_fd_sc_hd__a211oi_1 _36790_ (.A1(_06033_),
    .A2(_06036_),
    .B1(_07609_),
    .C1(_07610_),
    .Y(_09054_));
 sky130_fd_sc_hd__o21ba_1 _36791_ (.A1(_06028_),
    .A2(_07605_),
    .B1_N(_07606_),
    .X(_09055_));
 sky130_fd_sc_hd__o2bb2a_1 _36792_ (.A1_N(_04573_),
    .A2_N(_04574_),
    .B1(_07498_),
    .B2(_04550_),
    .X(_09056_));
 sky130_fd_sc_hd__o21a_1 _36793_ (.A1(_20896_),
    .A2(_20967_),
    .B1(_25236_),
    .X(_09057_));
 sky130_fd_sc_hd__or3b_2 _36794_ (.A(_23604_),
    .B(_19812_),
    .C_N(_01409_),
    .X(_09058_));
 sky130_fd_sc_hd__nor2_1 _36795_ (.A(_23604_),
    .B(_19812_),
    .Y(_09059_));
 sky130_fd_sc_hd__or2_1 _36796_ (.A(_01409_),
    .B(_09059_),
    .X(_09060_));
 sky130_fd_sc_hd__o211ai_4 _36797_ (.A1(_18813_),
    .A2(_09057_),
    .B1(_09058_),
    .C1(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__a221o_1 _36798_ (.A1(_20896_),
    .A2(_20967_),
    .B1(_09058_),
    .B2(_09060_),
    .C1(_09057_),
    .X(_09062_));
 sky130_fd_sc_hd__and2_1 _36799_ (.A(_09061_),
    .B(_09062_),
    .X(_09063_));
 sky130_fd_sc_hd__or3b_4 _36800_ (.A(_07500_),
    .B(_09056_),
    .C_N(_09063_),
    .X(_09065_));
 sky130_fd_sc_hd__o21bai_1 _36801_ (.A1(_07500_),
    .A2(_09056_),
    .B1_N(_09063_),
    .Y(_09066_));
 sky130_fd_sc_hd__nand3_2 _36802_ (.A(_09065_),
    .B(_07603_),
    .C(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__a32o_1 _36803_ (.A1(_07600_),
    .A2(_07598_),
    .A3(_07599_),
    .B1(_09066_),
    .B2(_09065_),
    .X(_09068_));
 sky130_fd_sc_hd__nand2_1 _36804_ (.A(_09067_),
    .B(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__o21ba_1 _36805_ (.A1(_07506_),
    .A2(_07527_),
    .B1_N(_07530_),
    .X(_09070_));
 sky130_fd_sc_hd__xnor2_1 _36806_ (.A(_09069_),
    .B(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__or2_1 _36807_ (.A(_09055_),
    .B(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__nand2_1 _36808_ (.A(_09071_),
    .B(_09055_),
    .Y(_09073_));
 sky130_fd_sc_hd__and2_1 _36809_ (.A(_09072_),
    .B(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__nor3_2 _36810_ (.A(_07610_),
    .B(_09054_),
    .C(_09074_),
    .Y(_09076_));
 sky130_fd_sc_hd__o21a_2 _36811_ (.A1(_07610_),
    .A2(_09054_),
    .B1(_09074_),
    .X(_09077_));
 sky130_fd_sc_hd__a211o_2 _36812_ (.A1(_07570_),
    .A2(_07576_),
    .B1(_09076_),
    .C1(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__o211ai_2 _36813_ (.A1(_09076_),
    .A2(_09077_),
    .B1(_07570_),
    .C1(_07576_),
    .Y(_09079_));
 sky130_fd_sc_hd__a22oi_4 _36814_ (.A1(_09052_),
    .A2(_07615_),
    .B1(_09078_),
    .B2(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36815_ (.A(_09079_),
    .X(_09081_));
 sky130_fd_sc_hd__and4b_1 _36816_ (.A_N(_07614_),
    .B(_07615_),
    .C(_09078_),
    .D(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__o2bb2ai_2 _36817_ (.A1_N(_09043_),
    .A2_N(_09051_),
    .B1(_09080_),
    .B2(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__o211a_1 _36818_ (.A1(_06038_),
    .A2(_06043_),
    .B1(_09052_),
    .C1(_09078_),
    .X(_09084_));
 sky130_fd_sc_hd__a21oi_1 _36819_ (.A1(_09084_),
    .A2(_09081_),
    .B1(_09080_),
    .Y(_09085_));
 sky130_fd_sc_hd__nand3_1 _36820_ (.A(_09043_),
    .B(_09051_),
    .C(_09085_),
    .Y(_09087_));
 sky130_fd_sc_hd__o21ai_1 _36821_ (.A1(_07485_),
    .A2(_07495_),
    .B1(_07584_),
    .Y(_09088_));
 sky130_fd_sc_hd__a21oi_1 _36822_ (.A1(_09088_),
    .A2(_07578_),
    .B1(_06076_),
    .Y(_09089_));
 sky130_fd_sc_hd__a22oi_4 _36823_ (.A1(_09089_),
    .A2(_07593_),
    .B1(_07590_),
    .B2(_07622_),
    .Y(_09090_));
 sky130_fd_sc_hd__a21oi_1 _36824_ (.A1(_09083_),
    .A2(_09087_),
    .B1(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__a21oi_2 _36825_ (.A1(_09049_),
    .A2(_09050_),
    .B1(_09044_),
    .Y(_09092_));
 sky130_fd_sc_hd__a21o_1 _36826_ (.A1(_09084_),
    .A2(_09081_),
    .B1(_09080_),
    .X(_09093_));
 sky130_fd_sc_hd__a31o_1 _36827_ (.A1(_09044_),
    .A2(_09049_),
    .A3(_09050_),
    .B1(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__o211a_1 _36828_ (.A1(_09092_),
    .A2(_09094_),
    .B1(_09083_),
    .C1(_09090_),
    .X(_09095_));
 sky130_fd_sc_hd__a21oi_2 _36829_ (.A1(net95),
    .A2(_07619_),
    .B1(_07617_),
    .Y(_09096_));
 sky130_fd_sc_hd__o21ai_1 _36830_ (.A1(_09091_),
    .A2(_09095_),
    .B1(_09096_),
    .Y(_09098_));
 sky130_fd_sc_hd__inv_2 _36831_ (.A(_09096_),
    .Y(_09099_));
 sky130_fd_sc_hd__a21o_1 _36832_ (.A1(_09083_),
    .A2(_09087_),
    .B1(_09090_),
    .X(_09100_));
 sky130_fd_sc_hd__o211ai_2 _36833_ (.A1(_09092_),
    .A2(_09094_),
    .B1(_09083_),
    .C1(_09090_),
    .Y(_09101_));
 sky130_fd_sc_hd__nand3_1 _36834_ (.A(_09099_),
    .B(_09100_),
    .C(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__and2_1 _36835_ (.A(_06050_),
    .B(_06074_),
    .X(_09103_));
 sky130_fd_sc_hd__a31o_1 _36836_ (.A1(_07625_),
    .A2(_07627_),
    .A3(_07623_),
    .B1(_09103_),
    .X(_09104_));
 sky130_fd_sc_hd__nand2_1 _36837_ (.A(_07628_),
    .B(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__a21o_1 _36838_ (.A1(_09098_),
    .A2(_09102_),
    .B1(_09105_),
    .X(_09106_));
 sky130_fd_sc_hd__nand3_1 _36839_ (.A(_09105_),
    .B(_09098_),
    .C(_09102_),
    .Y(_09107_));
 sky130_fd_sc_hd__and2_2 _36840_ (.A(_09106_),
    .B(_09107_),
    .X(_09109_));
 sky130_fd_sc_hd__xnor2_4 _36841_ (.A(_07640_),
    .B(_09109_),
    .Y(_00010_));
 sky130_fd_sc_hd__inv_2 _36842_ (.A(_09081_),
    .Y(_09110_));
 sky130_fd_sc_hd__inv_2 _36843_ (.A(_09078_),
    .Y(_09111_));
 sky130_fd_sc_hd__a21oi_1 _36844_ (.A1(_09052_),
    .A2(_07615_),
    .B1(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__a21oi_1 _36845_ (.A1(_09051_),
    .A2(_09085_),
    .B1(_09092_),
    .Y(_09113_));
 sky130_fd_sc_hd__nand3_1 _36846_ (.A(_08955_),
    .B(_09034_),
    .C(_09035_),
    .Y(_09114_));
 sky130_fd_sc_hd__inv_2 _36847_ (.A(_08131_),
    .Y(_09115_));
 sky130_fd_sc_hd__and3_1 _36848_ (.A(_08110_),
    .B(_08111_),
    .C(_08113_),
    .X(_09116_));
 sky130_fd_sc_hd__a31o_1 _36849_ (.A1(_08040_),
    .A2(_08042_),
    .A3(_08095_),
    .B1(_08091_),
    .X(_09117_));
 sky130_fd_sc_hd__o2bb2ai_4 _36850_ (.A1_N(_07932_),
    .A2_N(_07923_),
    .B1(_07907_),
    .B2(_07903_),
    .Y(_09119_));
 sky130_fd_sc_hd__or3_1 _36851_ (.A(_06417_),
    .B(_06418_),
    .C(_06413_),
    .X(_09120_));
 sky130_fd_sc_hd__buf_1 _36852_ (.A(_06416_),
    .X(_09121_));
 sky130_fd_sc_hd__a21o_1 _36853_ (.A1(_03368_),
    .A2(_09121_),
    .B1(_06412_),
    .X(_09122_));
 sky130_fd_sc_hd__o21ai_1 _36854_ (.A1(_03368_),
    .A2(_09121_),
    .B1(_06412_),
    .Y(_09123_));
 sky130_fd_sc_hd__buf_1 _36855_ (.A(_03360_),
    .X(_09124_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36856_ (.A(_09124_),
    .X(_09125_));
 sky130_fd_sc_hd__nand3_1 _36857_ (.A(_09122_),
    .B(_09123_),
    .C(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__a21o_1 _36858_ (.A1(_09122_),
    .A2(_09123_),
    .B1(_09124_),
    .X(_09127_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36859_ (.A(_09121_),
    .X(_09128_));
 sky130_fd_sc_hd__nand4_1 _36860_ (.A(_23755_),
    .B(_09128_),
    .C(_01788_),
    .D(_01789_),
    .Y(_09130_));
 sky130_fd_sc_hd__a31o_1 _36861_ (.A1(_01788_),
    .A2(_25337_),
    .A3(_09121_),
    .B1(_23755_),
    .X(_09131_));
 sky130_fd_sc_hd__and4_1 _36862_ (.A(_09126_),
    .B(_09127_),
    .C(_09130_),
    .D(_09131_),
    .X(_09132_));
 sky130_fd_sc_hd__a22o_1 _36863_ (.A1(_09126_),
    .A2(_09127_),
    .B1(_09130_),
    .B2(_09131_),
    .X(_09133_));
 sky130_fd_sc_hd__or2b_1 _36864_ (.A(_09132_),
    .B_N(_09133_),
    .X(_09134_));
 sky130_fd_sc_hd__o211a_1 _36865_ (.A1(_09120_),
    .A2(_07676_),
    .B1(_09134_),
    .C1(_07682_),
    .X(_09135_));
 sky130_fd_sc_hd__o21ai_1 _36866_ (.A1(_07676_),
    .A2(_09120_),
    .B1(_07682_),
    .Y(_09136_));
 sky130_fd_sc_hd__and3b_1 _36867_ (.A_N(_09132_),
    .B(_09133_),
    .C(_09136_),
    .X(_09137_));
 sky130_fd_sc_hd__nor2_2 _36868_ (.A(_09135_),
    .B(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__clkbuf_2 _36869_ (.A(_06430_),
    .X(_09139_));
 sky130_fd_sc_hd__buf_1 _36870_ (.A(_01740_),
    .X(_09141_));
 sky130_fd_sc_hd__a21oi_1 _36871_ (.A1(_01739_),
    .A2(_09139_),
    .B1(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__and3_1 _36872_ (.A(_01739_),
    .B(_09141_),
    .C(_06430_),
    .X(_09143_));
 sky130_fd_sc_hd__o21ai_1 _36873_ (.A1(_03354_),
    .A2(_07672_),
    .B1(_07670_),
    .Y(_09144_));
 sky130_fd_sc_hd__or3_1 _36874_ (.A(_09142_),
    .B(_09143_),
    .C(_09144_),
    .X(_09145_));
 sky130_fd_sc_hd__o21ai_1 _36875_ (.A1(_09142_),
    .A2(_09143_),
    .B1(_09144_),
    .Y(_09146_));
 sky130_fd_sc_hd__nand2_2 _36876_ (.A(_09145_),
    .B(_09146_),
    .Y(_09147_));
 sky130_fd_sc_hd__clkbuf_2 _36877_ (.A(_09139_),
    .X(_09148_));
 sky130_fd_sc_hd__and3b_2 _36878_ (.A_N(_23954_),
    .B(_04642_),
    .C(_09148_),
    .X(_09149_));
 sky130_fd_sc_hd__xnor2_4 _36879_ (.A(_09147_),
    .B(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__xnor2_4 _36880_ (.A(_09138_),
    .B(_09150_),
    .Y(_09152_));
 sky130_fd_sc_hd__clkbuf_2 _36881_ (.A(_07694_),
    .X(_09153_));
 sky130_fd_sc_hd__clkbuf_2 _36882_ (.A(_09153_),
    .X(_09154_));
 sky130_fd_sc_hd__and3_2 _36883_ (.A(_03312_),
    .B(_06335_),
    .C(_09153_),
    .X(_09155_));
 sky130_fd_sc_hd__a21oi_2 _36884_ (.A1(_06335_),
    .A2(_09153_),
    .B1(_03312_),
    .Y(_09156_));
 sky130_fd_sc_hd__o211a_1 _36885_ (.A1(_09155_),
    .A2(_09156_),
    .B1(_07873_),
    .C1(_07877_),
    .X(_09157_));
 sky130_fd_sc_hd__a211oi_4 _36886_ (.A1(_07873_),
    .A2(_07877_),
    .B1(_09155_),
    .C1(_09156_),
    .Y(_09158_));
 sky130_fd_sc_hd__o221a_1 _36887_ (.A1(_07696_),
    .A2(_09154_),
    .B1(_09157_),
    .B2(_09158_),
    .C1(_07701_),
    .X(_09159_));
 sky130_fd_sc_hd__a211oi_4 _36888_ (.A1(_07702_),
    .A2(_07701_),
    .B1(_09158_),
    .C1(_09157_),
    .Y(_09160_));
 sky130_fd_sc_hd__o211ai_1 _36889_ (.A1(_09159_),
    .A2(_09160_),
    .B1(_07866_),
    .C1(_07880_),
    .Y(_09161_));
 sky130_fd_sc_hd__a211o_1 _36890_ (.A1(_07866_),
    .A2(_07880_),
    .B1(_09159_),
    .C1(_09160_),
    .X(_09163_));
 sky130_fd_sc_hd__nand2_1 _36891_ (.A(_09161_),
    .B(_09163_),
    .Y(_09164_));
 sky130_fd_sc_hd__nor2_1 _36892_ (.A(_07705_),
    .B(_07707_),
    .Y(_09165_));
 sky130_fd_sc_hd__xor2_1 _36893_ (.A(_09164_),
    .B(_09165_),
    .X(_09166_));
 sky130_fd_sc_hd__nand2_1 _36894_ (.A(_09166_),
    .B(_07714_),
    .Y(_09167_));
 sky130_fd_sc_hd__or2_1 _36895_ (.A(_07714_),
    .B(_09166_),
    .X(_09168_));
 sky130_fd_sc_hd__nand2_2 _36896_ (.A(_09167_),
    .B(_09168_),
    .Y(_09169_));
 sky130_fd_sc_hd__xnor2_4 _36897_ (.A(_09152_),
    .B(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__a21oi_4 _36898_ (.A1(_07858_),
    .A2(_07897_),
    .B1(_07900_),
    .Y(_09171_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36899_ (.A(_09171_),
    .X(_09172_));
 sky130_fd_sc_hd__and2_2 _36900_ (.A(_07718_),
    .B(_07719_),
    .X(_09174_));
 sky130_fd_sc_hd__o21ai_1 _36901_ (.A1(_09172_),
    .A2(_09170_),
    .B1(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__a21oi_2 _36902_ (.A1(_09170_),
    .A2(_09172_),
    .B1(_09175_),
    .Y(_09176_));
 sky130_fd_sc_hd__inv_2 _36903_ (.A(_09170_),
    .Y(_09177_));
 sky130_fd_sc_hd__a21oi_1 _36904_ (.A1(_09177_),
    .A2(_09172_),
    .B1(_09174_),
    .Y(_09178_));
 sky130_fd_sc_hd__o21a_1 _36905_ (.A1(_09177_),
    .A2(_09172_),
    .B1(_09178_),
    .X(_09179_));
 sky130_fd_sc_hd__inv_2 _36906_ (.A(_07902_),
    .Y(_09180_));
 sky130_fd_sc_hd__a21oi_1 _36907_ (.A1(_07844_),
    .A2(_07847_),
    .B1(_07727_),
    .Y(_09181_));
 sky130_fd_sc_hd__o22ai_2 _36908_ (.A1(_07911_),
    .A2(_07912_),
    .B1(_09180_),
    .B2(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__o21a_1 _36909_ (.A1(_07882_),
    .A2(_07896_),
    .B1(_07894_),
    .X(_09183_));
 sky130_fd_sc_hd__inv_2 _36910_ (.A(_09183_),
    .Y(_09185_));
 sky130_fd_sc_hd__nand2_1 _36911_ (.A(_06341_),
    .B(\delay_line[9][15] ),
    .Y(_09186_));
 sky130_fd_sc_hd__nand2_1 _36912_ (.A(_06330_),
    .B(_23771_),
    .Y(_09187_));
 sky130_fd_sc_hd__a22o_1 _36913_ (.A1(\delay_line[10][10] ),
    .A2(_25375_),
    .B1(_09186_),
    .B2(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__nand4_1 _36914_ (.A(_09186_),
    .B(_09187_),
    .C(\delay_line[10][10] ),
    .D(_25375_),
    .Y(_09189_));
 sky130_fd_sc_hd__and3_1 _36915_ (.A(_09188_),
    .B(_07871_),
    .C(_09189_),
    .X(_09190_));
 sky130_fd_sc_hd__o2bb2a_1 _36916_ (.A1_N(_09189_),
    .A2_N(_09188_),
    .B1(_22458_),
    .B2(_07870_),
    .X(_09191_));
 sky130_fd_sc_hd__or2_1 _36917_ (.A(\delay_line[10][11] ),
    .B(\delay_line[10][12] ),
    .X(_09192_));
 sky130_fd_sc_hd__nand2_1 _36918_ (.A(_25370_),
    .B(_03281_),
    .Y(_09193_));
 sky130_fd_sc_hd__a21o_1 _36919_ (.A1(_09192_),
    .A2(_09193_),
    .B1(_04856_),
    .X(_09194_));
 sky130_fd_sc_hd__nand3_2 _36920_ (.A(_09192_),
    .B(_09193_),
    .C(_06364_),
    .Y(_09196_));
 sky130_fd_sc_hd__and3b_1 _36921_ (.A_N(_07862_),
    .B(_09194_),
    .C(_09196_),
    .X(_09197_));
 sky130_fd_sc_hd__a32oi_1 _36922_ (.A1(_07863_),
    .A2(_07859_),
    .A3(_07860_),
    .B1(_09194_),
    .B2(_09196_),
    .Y(_09198_));
 sky130_fd_sc_hd__or4_2 _36923_ (.A(_09190_),
    .B(_09191_),
    .C(_09197_),
    .D(_09198_),
    .X(_09199_));
 sky130_fd_sc_hd__o22ai_1 _36924_ (.A1(_09190_),
    .A2(_09191_),
    .B1(_09197_),
    .B2(_09198_),
    .Y(_09200_));
 sky130_fd_sc_hd__nand2_1 _36925_ (.A(_09199_),
    .B(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__buf_1 _36926_ (.A(_06353_),
    .X(_09202_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _36927_ (.A(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__and2b_1 _36928_ (.A_N(_00121_),
    .B(_09202_),
    .X(_09204_));
 sky130_fd_sc_hd__a31o_1 _36929_ (.A1(_00121_),
    .A2(_04796_),
    .A3(net399),
    .B1(_09204_),
    .X(_09205_));
 sky130_fd_sc_hd__a21oi_1 _36930_ (.A1(_07730_),
    .A2(_07884_),
    .B1(_09205_),
    .Y(_09207_));
 sky130_fd_sc_hd__a21oi_1 _36931_ (.A1(_07884_),
    .A2(_09205_),
    .B1(_09207_),
    .Y(_09208_));
 sky130_fd_sc_hd__a31o_1 _36932_ (.A1(_25373_),
    .A2(_01529_),
    .A3(_09203_),
    .B1(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__or3_1 _36933_ (.A(_07891_),
    .B(_06355_),
    .C(_09207_),
    .X(_09210_));
 sky130_fd_sc_hd__o211a_1 _36934_ (.A1(_07886_),
    .A2(_07890_),
    .B1(_09209_),
    .C1(_09210_),
    .X(_09211_));
 sky130_fd_sc_hd__a221oi_1 _36935_ (.A1(_06356_),
    .A2(_07889_),
    .B1(_09209_),
    .B2(_09210_),
    .C1(_07886_),
    .Y(_09212_));
 sky130_fd_sc_hd__nor2_1 _36936_ (.A(_09211_),
    .B(_09212_),
    .Y(_09213_));
 sky130_fd_sc_hd__xnor2_1 _36937_ (.A(_09201_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__or3_1 _36938_ (.A(_07737_),
    .B(_07845_),
    .C(_09214_),
    .X(_09215_));
 sky130_fd_sc_hd__o21ai_1 _36939_ (.A1(_07737_),
    .A2(_07845_),
    .B1(_09214_),
    .Y(_09216_));
 sky130_fd_sc_hd__nand2_1 _36940_ (.A(_09215_),
    .B(_09216_),
    .Y(_09218_));
 sky130_fd_sc_hd__nor2_1 _36941_ (.A(_09185_),
    .B(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__and2_1 _36942_ (.A(_09185_),
    .B(_09218_),
    .X(_09220_));
 sky130_fd_sc_hd__o2bb2ai_2 _36943_ (.A1_N(_07910_),
    .A2_N(_07842_),
    .B1(_07851_),
    .B2(_07850_),
    .Y(_09221_));
 sky130_fd_sc_hd__and2_1 _36944_ (.A(_03131_),
    .B(_07729_),
    .X(_09222_));
 sky130_fd_sc_hd__nor2_1 _36945_ (.A(_07729_),
    .B(_03131_),
    .Y(_09223_));
 sky130_fd_sc_hd__o21ai_2 _36946_ (.A1(_09222_),
    .A2(_09223_),
    .B1(_00108_),
    .Y(_09224_));
 sky130_fd_sc_hd__or3_1 _36947_ (.A(_00092_),
    .B(_09222_),
    .C(_09223_),
    .X(_09225_));
 sky130_fd_sc_hd__nand2_1 _36948_ (.A(_09224_),
    .B(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__a31o_1 _36949_ (.A1(_00108_),
    .A2(_04771_),
    .A3(_07826_),
    .B1(_07825_),
    .X(_09227_));
 sky130_fd_sc_hd__xnor2_2 _36950_ (.A(_09226_),
    .B(_09227_),
    .Y(_09229_));
 sky130_fd_sc_hd__and2_1 _36951_ (.A(_09229_),
    .B(_07734_),
    .X(_09230_));
 sky130_fd_sc_hd__nor2_1 _36952_ (.A(_07734_),
    .B(_09229_),
    .Y(_09231_));
 sky130_fd_sc_hd__a21boi_1 _36953_ (.A1(_07820_),
    .A2(_07822_),
    .B1_N(_07829_),
    .Y(_09232_));
 sky130_fd_sc_hd__inv_2 _36954_ (.A(\delay_line[4][13] ),
    .Y(_09233_));
 sky130_fd_sc_hd__or2_1 _36955_ (.A(_06225_),
    .B(_09233_),
    .X(_09234_));
 sky130_fd_sc_hd__or3b_2 _36956_ (.A(_04701_),
    .B(_07765_),
    .C_N(_07771_),
    .X(_09235_));
 sky130_fd_sc_hd__xnor2_2 _36957_ (.A(net433),
    .B(net432),
    .Y(_09236_));
 sky130_fd_sc_hd__and3_2 _36958_ (.A(_09234_),
    .B(_09235_),
    .C(_09236_),
    .X(_09237_));
 sky130_fd_sc_hd__inv_2 _36959_ (.A(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__a21oi_4 _36960_ (.A1(_09234_),
    .A2(_09235_),
    .B1(_09236_),
    .Y(_09240_));
 sky130_fd_sc_hd__inv_2 _36961_ (.A(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__inv_2 _36962_ (.A(_07774_),
    .Y(_09242_));
 sky130_fd_sc_hd__o211ai_4 _36963_ (.A1(_06230_),
    .A2(_06231_),
    .B1(_09242_),
    .C1(_06222_),
    .Y(_09243_));
 sky130_fd_sc_hd__o32a_4 _36964_ (.A1(_07767_),
    .A2(_06218_),
    .A3(_07774_),
    .B1(_07770_),
    .B2(_09233_),
    .X(_09244_));
 sky130_fd_sc_hd__a22oi_4 _36965_ (.A1(_09238_),
    .A2(_09241_),
    .B1(_09243_),
    .B2(_09244_),
    .Y(_09245_));
 sky130_fd_sc_hd__clkbuf_2 _36966_ (.A(_07751_),
    .X(_09246_));
 sky130_fd_sc_hd__xnor2_2 _36967_ (.A(net410),
    .B(net408),
    .Y(_09247_));
 sky130_fd_sc_hd__o21ai_1 _36968_ (.A1(_07746_),
    .A2(_07751_),
    .B1(_07749_),
    .Y(_09248_));
 sky130_fd_sc_hd__xnor2_1 _36969_ (.A(_09247_),
    .B(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__clkbuf_2 _36970_ (.A(_09249_),
    .X(_09251_));
 sky130_fd_sc_hd__o221ai_4 _36971_ (.A1(_09246_),
    .A2(_07748_),
    .B1(_07754_),
    .B2(_07759_),
    .C1(_09251_),
    .Y(_09252_));
 sky130_fd_sc_hd__nand2_1 _36972_ (.A(_07763_),
    .B(_07761_),
    .Y(_09253_));
 sky130_fd_sc_hd__or2_1 _36973_ (.A(_09246_),
    .B(_07748_),
    .X(_09254_));
 sky130_fd_sc_hd__a21o_1 _36974_ (.A1(_09253_),
    .A2(_09254_),
    .B1(_09251_),
    .X(_09255_));
 sky130_fd_sc_hd__nor2_2 _36975_ (.A(_09237_),
    .B(_09240_),
    .Y(_09256_));
 sky130_fd_sc_hd__nand3_4 _36976_ (.A(_09243_),
    .B(_09244_),
    .C(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__nand3_2 _36977_ (.A(_09252_),
    .B(_09255_),
    .C(_09257_),
    .Y(_09258_));
 sky130_fd_sc_hd__a31oi_2 _36978_ (.A1(_07781_),
    .A2(_07782_),
    .A3(_07783_),
    .B1(_07786_),
    .Y(_09259_));
 sky130_fd_sc_hd__o2bb2ai_1 _36979_ (.A1_N(_09244_),
    .A2_N(_09243_),
    .B1(_09240_),
    .B2(_09237_),
    .Y(_09260_));
 sky130_fd_sc_hd__a22o_1 _36980_ (.A1(_09252_),
    .A2(_09255_),
    .B1(_09260_),
    .B2(_09257_),
    .X(_09262_));
 sky130_fd_sc_hd__o221ai_4 _36981_ (.A1(_09245_),
    .A2(_09258_),
    .B1(_07798_),
    .B2(_09259_),
    .C1(_09262_),
    .Y(_09263_));
 sky130_fd_sc_hd__clkbuf_4 _36982_ (.A(_09260_),
    .X(_09264_));
 sky130_fd_sc_hd__o221a_1 _36983_ (.A1(_09246_),
    .A2(_07748_),
    .B1(_07754_),
    .B2(_07759_),
    .C1(_09251_),
    .X(_09265_));
 sky130_fd_sc_hd__a21oi_1 _36984_ (.A1(_09253_),
    .A2(_09254_),
    .B1(_09251_),
    .Y(_09266_));
 sky130_fd_sc_hd__nor2_2 _36985_ (.A(_09265_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__a21oi_4 _36986_ (.A1(_09264_),
    .A2(_09257_),
    .B1(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__nor2_1 _36987_ (.A(_09245_),
    .B(_09258_),
    .Y(_09269_));
 sky130_fd_sc_hd__a21oi_1 _36988_ (.A1(_07796_),
    .A2(_07784_),
    .B1(_07798_),
    .Y(_09270_));
 sky130_fd_sc_hd__o21ai_2 _36989_ (.A1(_09268_),
    .A2(_09269_),
    .B1(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__o21ai_1 _36990_ (.A1(_07798_),
    .A2(_07801_),
    .B1(_07796_),
    .Y(_09273_));
 sky130_fd_sc_hd__nand2_1 _36991_ (.A(_07803_),
    .B(_09273_),
    .Y(_09274_));
 sky130_fd_sc_hd__a21oi_1 _36992_ (.A1(_09263_),
    .A2(_09271_),
    .B1(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__clkbuf_2 _36993_ (.A(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__nand2_2 _36994_ (.A(_03198_),
    .B(_07805_),
    .Y(_09277_));
 sky130_fd_sc_hd__clkbuf_2 _36995_ (.A(_07809_),
    .X(_09278_));
 sky130_fd_sc_hd__nand2_1 _36996_ (.A(_04745_),
    .B(_09278_),
    .Y(_09279_));
 sky130_fd_sc_hd__and2_1 _36997_ (.A(_09277_),
    .B(_09279_),
    .X(_09280_));
 sky130_fd_sc_hd__or3_1 _36998_ (.A(_03198_),
    .B(_09278_),
    .C(_04751_),
    .X(_09281_));
 sky130_fd_sc_hd__o21ai_1 _36999_ (.A1(_07811_),
    .A2(_09280_),
    .B1(_09281_),
    .Y(_09282_));
 sky130_fd_sc_hd__a31o_1 _37000_ (.A1(_09274_),
    .A2(_09263_),
    .A3(_09271_),
    .B1(_09282_),
    .X(_09284_));
 sky130_fd_sc_hd__o21a_1 _37001_ (.A1(_07804_),
    .A2(_06268_),
    .B1(_07813_),
    .X(_09285_));
 sky130_fd_sc_hd__and3_1 _37002_ (.A(_09274_),
    .B(_09263_),
    .C(_09271_),
    .X(_09286_));
 sky130_fd_sc_hd__o21ai_1 _37003_ (.A1(_09276_),
    .A2(_09286_),
    .B1(_09282_),
    .Y(_09287_));
 sky130_fd_sc_hd__o221ai_4 _37004_ (.A1(_09276_),
    .A2(_09284_),
    .B1(_07792_),
    .B2(_09285_),
    .C1(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__o21a_1 _37005_ (.A1(_07811_),
    .A2(_09280_),
    .B1(_09281_),
    .X(_09289_));
 sky130_fd_sc_hd__o21ai_1 _37006_ (.A1(_09276_),
    .A2(_09286_),
    .B1(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__a21oi_1 _37007_ (.A1(_07833_),
    .A2(_07813_),
    .B1(_07792_),
    .Y(_09291_));
 sky130_fd_sc_hd__nand3_1 _37008_ (.A(_09274_),
    .B(_09263_),
    .C(_09271_),
    .Y(_09292_));
 sky130_fd_sc_hd__nand3b_1 _37009_ (.A_N(_09275_),
    .B(_09292_),
    .C(_09282_),
    .Y(_09293_));
 sky130_fd_sc_hd__nand3_1 _37010_ (.A(_09290_),
    .B(_09291_),
    .C(_09293_),
    .Y(_09295_));
 sky130_fd_sc_hd__or2_1 _37011_ (.A(_01549_),
    .B(_07805_),
    .X(_09296_));
 sky130_fd_sc_hd__nand2_1 _37012_ (.A(_01549_),
    .B(_07807_),
    .Y(_09297_));
 sky130_fd_sc_hd__a32o_1 _37013_ (.A1(_01630_),
    .A2(_04751_),
    .A3(_07807_),
    .B1(_09296_),
    .B2(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__o31a_1 _37014_ (.A1(_04762_),
    .A2(_03206_),
    .A3(_06280_),
    .B1(_09298_),
    .X(_09299_));
 sky130_fd_sc_hd__and3_1 _37015_ (.A(_00096_),
    .B(_06287_),
    .C(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__a21oi_1 _37016_ (.A1(_03221_),
    .A2(_06287_),
    .B1(_09299_),
    .Y(_09301_));
 sky130_fd_sc_hd__nor2_1 _37017_ (.A(_09300_),
    .B(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__nand3_2 _37018_ (.A(_09288_),
    .B(_09295_),
    .C(_09302_),
    .Y(_09303_));
 sky130_fd_sc_hd__a21o_1 _37019_ (.A1(_09288_),
    .A2(_09295_),
    .B1(_09302_),
    .X(_09304_));
 sky130_fd_sc_hd__o211ai_4 _37020_ (.A1(_07831_),
    .A2(_09232_),
    .B1(_09303_),
    .C1(_09304_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand2_1 _37021_ (.A(_09303_),
    .B(_09302_),
    .Y(_09307_));
 sky130_fd_sc_hd__o211ai_1 _37022_ (.A1(_09300_),
    .A2(_09301_),
    .B1(_09288_),
    .C1(_09295_),
    .Y(_09308_));
 sky130_fd_sc_hd__a21oi_1 _37023_ (.A1(_07823_),
    .A2(_07829_),
    .B1(_07831_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand3_2 _37024_ (.A(_09307_),
    .B(_09308_),
    .C(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__o211ai_4 _37025_ (.A1(_09230_),
    .A2(_09231_),
    .B1(_09306_),
    .C1(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__and4_1 _37026_ (.A(_07732_),
    .B(_09229_),
    .C(_07731_),
    .D(_06299_),
    .X(_09312_));
 sky130_fd_sc_hd__a31oi_2 _37027_ (.A1(_06299_),
    .A2(_07732_),
    .A3(_07731_),
    .B1(_09229_),
    .Y(_09313_));
 sky130_fd_sc_hd__o2bb2ai_2 _37028_ (.A1_N(_09306_),
    .A2_N(_09310_),
    .B1(_09312_),
    .B2(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__nand3_2 _37029_ (.A(_09221_),
    .B(_09311_),
    .C(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__o21ai_1 _37030_ (.A1(_07739_),
    .A2(_07740_),
    .B1(_07841_),
    .Y(_09317_));
 sky130_fd_sc_hd__o211ai_1 _37031_ (.A1(_09312_),
    .A2(_09313_),
    .B1(_09306_),
    .C1(_09310_),
    .Y(_09318_));
 sky130_fd_sc_hd__o2bb2ai_1 _37032_ (.A1_N(_09306_),
    .A2_N(_09310_),
    .B1(_09230_),
    .B2(_09231_),
    .Y(_09319_));
 sky130_fd_sc_hd__nand4_1 _37033_ (.A(_07837_),
    .B(_09317_),
    .C(_09318_),
    .D(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__clkbuf_2 _37034_ (.A(_09320_),
    .X(_09321_));
 sky130_fd_sc_hd__o211ai_2 _37035_ (.A1(_09219_),
    .A2(_09220_),
    .B1(_09315_),
    .C1(_09321_),
    .Y(_09322_));
 sky130_fd_sc_hd__nor2_1 _37036_ (.A(_09183_),
    .B(_09218_),
    .Y(_09323_));
 sky130_fd_sc_hd__o211a_1 _37037_ (.A1(_07882_),
    .A2(_07896_),
    .B1(_09218_),
    .C1(_07894_),
    .X(_09324_));
 sky130_fd_sc_hd__o2bb2ai_1 _37038_ (.A1_N(_09315_),
    .A2_N(_09320_),
    .B1(_09323_),
    .B2(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__nand3_4 _37039_ (.A(_09182_),
    .B(_09322_),
    .C(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__clkbuf_2 _37040_ (.A(_09326_),
    .X(_09328_));
 sky130_fd_sc_hd__a21boi_2 _37041_ (.A1(_07856_),
    .A2(_07902_),
    .B1_N(_07848_),
    .Y(_09329_));
 sky130_fd_sc_hd__o211ai_2 _37042_ (.A1(_09323_),
    .A2(_09324_),
    .B1(_09315_),
    .C1(_09321_),
    .Y(_09330_));
 sky130_fd_sc_hd__o2bb2ai_1 _37043_ (.A1_N(_09315_),
    .A2_N(_09321_),
    .B1(_09219_),
    .B2(_09220_),
    .Y(_09331_));
 sky130_fd_sc_hd__nand3_4 _37044_ (.A(_09329_),
    .B(_09330_),
    .C(_09331_),
    .Y(_09332_));
 sky130_fd_sc_hd__o211ai_4 _37045_ (.A1(_09176_),
    .A2(_09179_),
    .B1(_09328_),
    .C1(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__nand2_1 _37046_ (.A(_09326_),
    .B(_09332_),
    .Y(_09334_));
 sky130_fd_sc_hd__nor2_1 _37047_ (.A(_09176_),
    .B(_09179_),
    .Y(_09335_));
 sky130_fd_sc_hd__nand2_1 _37048_ (.A(_09334_),
    .B(_09335_),
    .Y(_09336_));
 sky130_fd_sc_hd__nand3_2 _37049_ (.A(_09119_),
    .B(_09333_),
    .C(_09336_),
    .Y(_09337_));
 sky130_fd_sc_hd__a2bb2oi_1 _37050_ (.A1_N(_06391_),
    .A2_N(_07905_),
    .B1(_07913_),
    .B2(_07917_),
    .Y(_09339_));
 sky130_fd_sc_hd__a21oi_2 _37051_ (.A1(_07923_),
    .A2(_07932_),
    .B1(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__nand3_1 _37052_ (.A(_09328_),
    .B(_09332_),
    .C(_09335_),
    .Y(_09341_));
 sky130_fd_sc_hd__o2bb2ai_1 _37053_ (.A1_N(_09328_),
    .A2_N(_09332_),
    .B1(_09176_),
    .B2(_09179_),
    .Y(_09342_));
 sky130_fd_sc_hd__nand3_1 _37054_ (.A(_09340_),
    .B(_09341_),
    .C(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__buf_6 _37055_ (.A(_09343_),
    .X(_09344_));
 sky130_fd_sc_hd__or2_1 _37056_ (.A(_07960_),
    .B(_07965_),
    .X(_09345_));
 sky130_fd_sc_hd__buf_1 _37057_ (.A(_07955_),
    .X(_09346_));
 sky130_fd_sc_hd__or4_2 _37058_ (.A(_06098_),
    .B(_06099_),
    .C(_06104_),
    .D(_07958_),
    .X(_09347_));
 sky130_fd_sc_hd__and2b_1 _37059_ (.A_N(_07683_),
    .B(_07685_),
    .X(_09348_));
 sky130_fd_sc_hd__o2111ai_2 _37060_ (.A1(_06429_),
    .A2(_06431_),
    .B1(_06433_),
    .C1(_07659_),
    .D1(_07658_),
    .Y(_09350_));
 sky130_fd_sc_hd__nor2_1 _37061_ (.A(_01745_),
    .B(_03338_),
    .Y(_09351_));
 sky130_fd_sc_hd__and2_1 _37062_ (.A(_01744_),
    .B(_03334_),
    .X(_09352_));
 sky130_fd_sc_hd__o21bai_1 _37063_ (.A1(_09351_),
    .A2(_09352_),
    .B1_N(_01747_),
    .Y(_09353_));
 sky130_fd_sc_hd__or3b_1 _37064_ (.A(_09351_),
    .B(_09352_),
    .C_N(_25297_),
    .X(_09354_));
 sky130_fd_sc_hd__clkbuf_2 _37065_ (.A(_06091_),
    .X(_09355_));
 sky130_fd_sc_hd__or2_1 _37066_ (.A(\delay_line[7][9] ),
    .B(_06090_),
    .X(_09356_));
 sky130_fd_sc_hd__nand2_1 _37067_ (.A(_06091_),
    .B(_22525_),
    .Y(_09357_));
 sky130_fd_sc_hd__a21bo_1 _37068_ (.A1(_07950_),
    .A2(_04973_),
    .B1_N(_07951_),
    .X(_09358_));
 sky130_fd_sc_hd__a21oi_2 _37069_ (.A1(_09356_),
    .A2(_09357_),
    .B1(_09358_),
    .Y(_09359_));
 sky130_fd_sc_hd__and3_1 _37070_ (.A(_09358_),
    .B(_09356_),
    .C(_09357_),
    .X(_09361_));
 sky130_fd_sc_hd__or4_1 _37071_ (.A(_03412_),
    .B(_09355_),
    .C(_09359_),
    .D(_09361_),
    .X(_09362_));
 sky130_fd_sc_hd__o21ai_1 _37072_ (.A1(_09359_),
    .A2(_09361_),
    .B1(_07940_),
    .Y(_09363_));
 sky130_fd_sc_hd__and4_1 _37073_ (.A(_09353_),
    .B(_09354_),
    .C(_09362_),
    .D(_09363_),
    .X(_09364_));
 sky130_fd_sc_hd__a22oi_2 _37074_ (.A1(_09353_),
    .A2(_09354_),
    .B1(_09362_),
    .B2(_09363_),
    .Y(_09365_));
 sky130_fd_sc_hd__a211o_1 _37075_ (.A1(_07659_),
    .A2(_09350_),
    .B1(_09364_),
    .C1(_09365_),
    .X(_09366_));
 sky130_fd_sc_hd__o211ai_2 _37076_ (.A1(_09364_),
    .A2(_09365_),
    .B1(_07659_),
    .C1(_09350_),
    .Y(_09367_));
 sky130_fd_sc_hd__nand3_1 _37077_ (.A(_09366_),
    .B(_09367_),
    .C(_09346_),
    .Y(_09368_));
 sky130_fd_sc_hd__a21o_1 _37078_ (.A1(_09366_),
    .A2(_09367_),
    .B1(_09346_),
    .X(_09369_));
 sky130_fd_sc_hd__nand2_1 _37079_ (.A(_09368_),
    .B(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__nand2_1 _37080_ (.A(_09348_),
    .B(_09370_),
    .Y(_09372_));
 sky130_fd_sc_hd__or2_1 _37081_ (.A(_09370_),
    .B(_09348_),
    .X(_09373_));
 sky130_fd_sc_hd__nand2_1 _37082_ (.A(_09372_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__o311a_1 _37083_ (.A1(_07939_),
    .A2(_09346_),
    .A3(_07956_),
    .B1(_09347_),
    .C1(_09374_),
    .X(_09375_));
 sky130_fd_sc_hd__or3_1 _37084_ (.A(_07939_),
    .B(_09346_),
    .C(_07956_),
    .X(_09376_));
 sky130_fd_sc_hd__a21oi_2 _37085_ (.A1(_09376_),
    .A2(_09347_),
    .B1(_09374_),
    .Y(_09377_));
 sky130_fd_sc_hd__a211oi_2 _37086_ (.A1(_07961_),
    .A2(_09345_),
    .B1(_09375_),
    .C1(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__o221ai_4 _37087_ (.A1(_07960_),
    .A2(_07965_),
    .B1(_09377_),
    .B2(_09375_),
    .C1(_07961_),
    .Y(_09379_));
 sky130_fd_sc_hd__inv_2 _37088_ (.A(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__a21oi_1 _37089_ (.A1(_01863_),
    .A2(_07996_),
    .B1(_07972_),
    .Y(_09381_));
 sky130_fd_sc_hd__and3_1 _37090_ (.A(_01863_),
    .B(_07996_),
    .C(_07972_),
    .X(_09383_));
 sky130_fd_sc_hd__nor2_1 _37091_ (.A(_09381_),
    .B(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__xor2_1 _37092_ (.A(_08000_),
    .B(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__a21bo_1 _37093_ (.A1(_07977_),
    .A2(_07976_),
    .B1_N(_07974_),
    .X(_09386_));
 sky130_fd_sc_hd__xor2_1 _37094_ (.A(_09385_),
    .B(_09386_),
    .X(_09387_));
 sky130_fd_sc_hd__a311oi_1 _37095_ (.A1(_08001_),
    .A2(_07995_),
    .A3(_08000_),
    .B1(net250),
    .C1(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__o21a_1 _37096_ (.A1(net250),
    .A2(_08002_),
    .B1(_09387_),
    .X(_09389_));
 sky130_fd_sc_hd__nor2_1 _37097_ (.A(_09388_),
    .B(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__clkbuf_2 _37098_ (.A(_06151_),
    .X(_09391_));
 sky130_fd_sc_hd__a41o_1 _37099_ (.A1(_09391_),
    .A2(_06146_),
    .A3(_06149_),
    .A4(_07980_),
    .B1(_07983_),
    .X(_09392_));
 sky130_fd_sc_hd__nor2_1 _37100_ (.A(_09390_),
    .B(_09392_),
    .Y(_09394_));
 sky130_fd_sc_hd__and4_1 _37101_ (.A(_06146_),
    .B(_07980_),
    .C(_06149_),
    .D(_06151_),
    .X(_09395_));
 sky130_fd_sc_hd__o21a_1 _37102_ (.A1(_09395_),
    .A2(_07983_),
    .B1(_09390_),
    .X(_09396_));
 sky130_fd_sc_hd__or2_2 _37103_ (.A(_09394_),
    .B(_09396_),
    .X(_09397_));
 sky130_fd_sc_hd__o31a_2 _37104_ (.A1(_08013_),
    .A2(_08014_),
    .A3(_08016_),
    .B1(_08018_),
    .X(_09398_));
 sky130_fd_sc_hd__buf_1 _37105_ (.A(\delay_line[5][15] ),
    .X(_09399_));
 sky130_fd_sc_hd__nor2_1 _37106_ (.A(_01872_),
    .B(_06147_),
    .Y(_09400_));
 sky130_fd_sc_hd__and2_1 _37107_ (.A(_06147_),
    .B(_01872_),
    .X(_09401_));
 sky130_fd_sc_hd__nor2_1 _37108_ (.A(_09400_),
    .B(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__nor2_1 _37109_ (.A(_09399_),
    .B(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__and2_1 _37110_ (.A(_09399_),
    .B(_09402_),
    .X(_09405_));
 sky130_fd_sc_hd__or2b_1 _37111_ (.A(_24062_),
    .B_N(_09399_),
    .X(_09406_));
 sky130_fd_sc_hd__or2b_1 _37112_ (.A(_09399_),
    .B_N(_24062_),
    .X(_09407_));
 sky130_fd_sc_hd__nand3_1 _37113_ (.A(_07991_),
    .B(_09406_),
    .C(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__a21o_1 _37114_ (.A1(_09406_),
    .A2(_09407_),
    .B1(_07991_),
    .X(_09409_));
 sky130_fd_sc_hd__or4bb_1 _37115_ (.A(_09403_),
    .B(_09405_),
    .C_N(_09408_),
    .D_N(_09409_),
    .X(_09410_));
 sky130_fd_sc_hd__a2bb2o_1 _37116_ (.A1_N(_09403_),
    .A2_N(_09405_),
    .B1(_09408_),
    .B2(_09409_),
    .X(_09411_));
 sky130_fd_sc_hd__and2_1 _37117_ (.A(_09410_),
    .B(_09411_),
    .X(_09412_));
 sky130_fd_sc_hd__a21boi_2 _37118_ (.A1(_08011_),
    .A2(_08012_),
    .B1_N(_08009_),
    .Y(_09413_));
 sky130_fd_sc_hd__o21ai_2 _37119_ (.A1(_08010_),
    .A2(_06097_),
    .B1(_04928_),
    .Y(_09414_));
 sky130_fd_sc_hd__o21a_1 _37120_ (.A1(net426),
    .A2(_04978_),
    .B1(_07946_),
    .X(_09416_));
 sky130_fd_sc_hd__nor3_1 _37121_ (.A(net426),
    .B(_04978_),
    .C(_07946_),
    .Y(_09417_));
 sky130_fd_sc_hd__nand3b_1 _37122_ (.A_N(_06089_),
    .B(_07944_),
    .C(_07945_),
    .Y(_09418_));
 sky130_fd_sc_hd__o211ai_1 _37123_ (.A1(_09416_),
    .A2(_09417_),
    .B1(_07945_),
    .C1(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__a211o_1 _37124_ (.A1(_07945_),
    .A2(_09418_),
    .B1(_09416_),
    .C1(_09417_),
    .X(_09420_));
 sky130_fd_sc_hd__nand2_2 _37125_ (.A(_09419_),
    .B(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__xor2_2 _37126_ (.A(_09414_),
    .B(_09421_),
    .X(_09422_));
 sky130_fd_sc_hd__xor2_2 _37127_ (.A(_09413_),
    .B(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__xor2_2 _37128_ (.A(_09412_),
    .B(_09423_),
    .X(_09424_));
 sky130_fd_sc_hd__xnor2_2 _37129_ (.A(_09398_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__xor2_2 _37130_ (.A(_09397_),
    .B(_09425_),
    .X(_09427_));
 sky130_fd_sc_hd__o21bai_1 _37131_ (.A1(_09378_),
    .A2(_09380_),
    .B1_N(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand3b_1 _37132_ (.A_N(_09378_),
    .B(_09379_),
    .C(_09427_),
    .Y(_09429_));
 sky130_fd_sc_hd__a211oi_1 _37133_ (.A1(_09428_),
    .A2(_09429_),
    .B1(_07721_),
    .C1(_07725_),
    .Y(_09430_));
 sky130_fd_sc_hd__o211ai_2 _37134_ (.A1(_07721_),
    .A2(_07725_),
    .B1(_09428_),
    .C1(_09429_),
    .Y(_09431_));
 sky130_fd_sc_hd__nand2b_1 _37135_ (.A_N(_09430_),
    .B(_09431_),
    .Y(_09432_));
 sky130_fd_sc_hd__xor2_1 _37136_ (.A(_07962_),
    .B(_07965_),
    .X(_09433_));
 sky130_fd_sc_hd__a21oi_2 _37137_ (.A1(_07937_),
    .A2(_09433_),
    .B1(_08024_),
    .Y(_09434_));
 sky130_fd_sc_hd__and2_1 _37138_ (.A(_09432_),
    .B(_09434_),
    .X(_09435_));
 sky130_fd_sc_hd__or2_1 _37139_ (.A(_09434_),
    .B(_09432_),
    .X(_09436_));
 sky130_fd_sc_hd__and2b_1 _37140_ (.A_N(_09435_),
    .B(_09436_),
    .X(_09438_));
 sky130_fd_sc_hd__buf_1 _37141_ (.A(_09438_),
    .X(_09439_));
 sky130_fd_sc_hd__a21boi_2 _37142_ (.A1(_09337_),
    .A2(_09344_),
    .B1_N(_09439_),
    .Y(_09440_));
 sky130_fd_sc_hd__nand2_1 _37143_ (.A(_07928_),
    .B(_08031_),
    .Y(_09441_));
 sky130_fd_sc_hd__inv_2 _37144_ (.A(_09436_),
    .Y(_09442_));
 sky130_fd_sc_hd__o211ai_1 _37145_ (.A1(_09435_),
    .A2(_09442_),
    .B1(_09344_),
    .C1(_09337_),
    .Y(_09443_));
 sky130_fd_sc_hd__nand3_2 _37146_ (.A(_07934_),
    .B(_09441_),
    .C(_09443_),
    .Y(_09444_));
 sky130_fd_sc_hd__and3_2 _37147_ (.A(_07929_),
    .B(_07930_),
    .C(_07933_),
    .X(_09445_));
 sky130_fd_sc_hd__a31oi_4 _37148_ (.A1(_07652_),
    .A2(_07919_),
    .A3(_07926_),
    .B1(_08039_),
    .Y(_09446_));
 sky130_fd_sc_hd__nand3_1 _37149_ (.A(_09337_),
    .B(_09344_),
    .C(_09439_),
    .Y(_09447_));
 sky130_fd_sc_hd__a21o_1 _37150_ (.A1(_09337_),
    .A2(_09344_),
    .B1(_09439_),
    .X(_09449_));
 sky130_fd_sc_hd__o211ai_4 _37151_ (.A1(_09445_),
    .A2(_09446_),
    .B1(_09447_),
    .C1(_09449_),
    .Y(_09450_));
 sky130_fd_sc_hd__xor2_1 _37152_ (.A(_08076_),
    .B(_08077_),
    .X(_09451_));
 sky130_fd_sc_hd__a21o_1 _37153_ (.A1(_06121_),
    .A2(_06189_),
    .B1(_08027_),
    .X(_09452_));
 sky130_fd_sc_hd__a21boi_2 _37154_ (.A1(_08075_),
    .A2(_08077_),
    .B1_N(_08073_),
    .Y(_09453_));
 sky130_fd_sc_hd__o31a_1 _37155_ (.A1(_08050_),
    .A2(net199),
    .A3(_08060_),
    .B1(_08065_),
    .X(_09454_));
 sky130_fd_sc_hd__clkbuf_2 _37156_ (.A(_06510_),
    .X(_09455_));
 sky130_fd_sc_hd__or3_1 _37157_ (.A(_08047_),
    .B(_04908_),
    .C(_05024_),
    .X(_09456_));
 sky130_fd_sc_hd__o21ai_1 _37158_ (.A1(_08047_),
    .A2(_08046_),
    .B1(_04908_),
    .Y(_09457_));
 sky130_fd_sc_hd__and4bb_1 _37159_ (.A_N(_08051_),
    .B_N(_08058_),
    .C(_09456_),
    .D(_09457_),
    .X(_09458_));
 sky130_fd_sc_hd__a2bb2oi_2 _37160_ (.A1_N(_08051_),
    .A2_N(_08058_),
    .B1(_09456_),
    .B2(_09457_),
    .Y(_09460_));
 sky130_fd_sc_hd__o2111ai_2 _37161_ (.A1(_09455_),
    .A2(_05023_),
    .B1(_01494_),
    .C1(_08047_),
    .D1(_08054_),
    .Y(_09461_));
 sky130_fd_sc_hd__o221ai_1 _37162_ (.A1(_09455_),
    .A2(_05023_),
    .B1(_09458_),
    .B2(_09460_),
    .C1(_09461_),
    .Y(_09462_));
 sky130_fd_sc_hd__a211o_1 _37163_ (.A1(_08055_),
    .A2(_09461_),
    .B1(_09458_),
    .C1(_09460_),
    .X(_09463_));
 sky130_fd_sc_hd__nand2_1 _37164_ (.A(_09462_),
    .B(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__a21oi_1 _37165_ (.A1(_07988_),
    .A2(_07968_),
    .B1(_07987_),
    .Y(_09465_));
 sky130_fd_sc_hd__xnor2_1 _37166_ (.A(_09464_),
    .B(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__xor2_1 _37167_ (.A(_09454_),
    .B(_09466_),
    .X(_09467_));
 sky130_fd_sc_hd__nand2_1 _37168_ (.A(_07989_),
    .B(_08022_),
    .Y(_09468_));
 sky130_fd_sc_hd__o21ai_2 _37169_ (.A1(_07990_),
    .A2(_08021_),
    .B1(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__nand2_1 _37170_ (.A(_09467_),
    .B(_09469_),
    .Y(_09471_));
 sky130_fd_sc_hd__or2_1 _37171_ (.A(_09469_),
    .B(_09467_),
    .X(_09472_));
 sky130_fd_sc_hd__nand2_1 _37172_ (.A(_09471_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__nor2_1 _37173_ (.A(_08067_),
    .B(_08071_),
    .Y(_09474_));
 sky130_fd_sc_hd__xnor2_2 _37174_ (.A(_09473_),
    .B(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__xnor2_1 _37175_ (.A(_09453_),
    .B(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__a21oi_2 _37176_ (.A1(_08028_),
    .A2(_09452_),
    .B1(_09476_),
    .Y(_09477_));
 sky130_fd_sc_hd__nand3_1 _37177_ (.A(_08028_),
    .B(_09476_),
    .C(_09452_),
    .Y(_09478_));
 sky130_fd_sc_hd__nand2b_1 _37178_ (.A_N(_09477_),
    .B(_09478_),
    .Y(_09479_));
 sky130_fd_sc_hd__o21a_1 _37179_ (.A1(_08045_),
    .A2(_09451_),
    .B1(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__nor3_1 _37180_ (.A(_08045_),
    .B(_09451_),
    .C(_09479_),
    .Y(_09482_));
 sky130_fd_sc_hd__nor2_1 _37181_ (.A(_09480_),
    .B(net89),
    .Y(_09483_));
 sky130_fd_sc_hd__o211ai_1 _37182_ (.A1(_09440_),
    .A2(_09444_),
    .B1(_09450_),
    .C1(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__o21ai_1 _37183_ (.A1(_09440_),
    .A2(_09444_),
    .B1(_09450_),
    .Y(_09485_));
 sky130_fd_sc_hd__nor2_1 _37184_ (.A(_08045_),
    .B(_09451_),
    .Y(_09486_));
 sky130_fd_sc_hd__xor2_1 _37185_ (.A(_09486_),
    .B(_09479_),
    .X(_09487_));
 sky130_fd_sc_hd__nand2_1 _37186_ (.A(_09485_),
    .B(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__nand4_2 _37187_ (.A(_08036_),
    .B(_09117_),
    .C(_09484_),
    .D(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__a31oi_2 _37188_ (.A1(_08040_),
    .A2(_08042_),
    .A3(_08095_),
    .B1(_08091_),
    .Y(_09490_));
 sky130_fd_sc_hd__o221ai_4 _37189_ (.A1(_09440_),
    .A2(_09444_),
    .B1(_09480_),
    .B2(_09482_),
    .C1(_09450_),
    .Y(_09491_));
 sky130_fd_sc_hd__nand2_1 _37190_ (.A(_09485_),
    .B(_09483_),
    .Y(_09493_));
 sky130_fd_sc_hd__o211ai_4 _37191_ (.A1(_08097_),
    .A2(_09490_),
    .B1(_09491_),
    .C1(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__or2_1 _37192_ (.A(_06538_),
    .B(_06539_),
    .X(_09495_));
 sky130_fd_sc_hd__o21ba_1 _37193_ (.A1(_06504_),
    .A2(_09495_),
    .B1_N(_08082_),
    .X(_09496_));
 sky130_fd_sc_hd__nor2_1 _37194_ (.A(_08083_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__a21oi_2 _37195_ (.A1(_09489_),
    .A2(_09494_),
    .B1(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__a21o_1 _37196_ (.A1(_08086_),
    .A2(_08043_),
    .B1(_08097_),
    .X(_09499_));
 sky130_fd_sc_hd__a21oi_2 _37197_ (.A1(_09491_),
    .A2(_09493_),
    .B1(_09499_),
    .Y(_09500_));
 sky130_fd_sc_hd__nand2_1 _37198_ (.A(_09494_),
    .B(_09497_),
    .Y(_09501_));
 sky130_fd_sc_hd__nor2_1 _37199_ (.A(_09500_),
    .B(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__nor2_1 _37200_ (.A(_08104_),
    .B(_08112_),
    .Y(_09504_));
 sky130_fd_sc_hd__o21ai_4 _37201_ (.A1(_09498_),
    .A2(_09502_),
    .B1(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__o2bb2ai_1 _37202_ (.A1_N(_09489_),
    .A2_N(_09494_),
    .B1(_09496_),
    .B2(_08083_),
    .Y(_09506_));
 sky130_fd_sc_hd__o221ai_2 _37203_ (.A1(_09500_),
    .A2(_09501_),
    .B1(_08104_),
    .B2(_08112_),
    .C1(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__clkbuf_2 _37204_ (.A(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__nand2_1 _37205_ (.A(_09505_),
    .B(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__o21bai_1 _37206_ (.A1(_09116_),
    .A2(_08121_),
    .B1_N(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37207_ (.A(_09509_),
    .X(_09511_));
 sky130_fd_sc_hd__o211ai_2 _37208_ (.A1(_08106_),
    .A2(_08108_),
    .B1(_09511_),
    .C1(_08130_),
    .Y(_09512_));
 sky130_fd_sc_hd__a41o_2 _37209_ (.A1(_08212_),
    .A2(_08213_),
    .A3(_08221_),
    .A4(_08222_),
    .B1(_08225_),
    .X(_09513_));
 sky130_fd_sc_hd__a21oi_2 _37210_ (.A1(_09510_),
    .A2(_09512_),
    .B1(_09513_),
    .Y(_09515_));
 sky130_fd_sc_hd__a21oi_1 _37211_ (.A1(_07650_),
    .A2(_08101_),
    .B1(_08108_),
    .Y(_09516_));
 sky130_fd_sc_hd__a22oi_2 _37212_ (.A1(_08113_),
    .A2(_09516_),
    .B1(_08127_),
    .B2(_08128_),
    .Y(_09517_));
 sky130_fd_sc_hd__inv_2 _37213_ (.A(_09513_),
    .Y(_09518_));
 sky130_fd_sc_hd__o21bai_2 _37214_ (.A1(_09511_),
    .A2(_09517_),
    .B1_N(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__a21oi_1 _37215_ (.A1(_09511_),
    .A2(_09517_),
    .B1(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37216_ (.A(_06586_),
    .X(_09521_));
 sky130_fd_sc_hd__o21bai_4 _37217_ (.A1(_09515_),
    .A2(_09520_),
    .B1_N(_09521_),
    .Y(_09522_));
 sky130_fd_sc_hd__clkbuf_2 _37218_ (.A(_08114_),
    .X(_09523_));
 sky130_fd_sc_hd__and3_1 _37219_ (.A(_09523_),
    .B(_08130_),
    .C(_09511_),
    .X(_09524_));
 sky130_fd_sc_hd__buf_2 _37220_ (.A(_09521_),
    .X(_09526_));
 sky130_fd_sc_hd__a21o_1 _37221_ (.A1(_09510_),
    .A2(_09512_),
    .B1(_09513_),
    .X(_09527_));
 sky130_fd_sc_hd__o211ai_4 _37222_ (.A1(_09524_),
    .A2(_09519_),
    .B1(_09526_),
    .C1(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__o32a_1 _37223_ (.A1(_08225_),
    .A2(_08227_),
    .A3(_08276_),
    .B1(_08273_),
    .B2(_08230_),
    .X(_09529_));
 sky130_fd_sc_hd__a21boi_2 _37224_ (.A1(_09522_),
    .A2(_09528_),
    .B1_N(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__o211a_2 _37225_ (.A1(_08274_),
    .A2(_08277_),
    .B1(_09522_),
    .C1(_09528_),
    .X(_09531_));
 sky130_fd_sc_hd__o22ai_2 _37226_ (.A1(_09115_),
    .A2(_08141_),
    .B1(_09530_),
    .B2(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__nand2_1 _37227_ (.A(_09522_),
    .B(_09528_),
    .Y(_09533_));
 sky130_fd_sc_hd__nand2_1 _37228_ (.A(_09533_),
    .B(_09529_),
    .Y(_09534_));
 sky130_fd_sc_hd__o211ai_2 _37229_ (.A1(_08274_),
    .A2(_08277_),
    .B1(_09522_),
    .C1(_09528_),
    .Y(_09535_));
 sky130_fd_sc_hd__a21o_1 _37230_ (.A1(_08133_),
    .A2(_08123_),
    .B1(_09115_),
    .X(_09537_));
 sky130_fd_sc_hd__inv_2 _37231_ (.A(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__nand3_1 _37232_ (.A(_09534_),
    .B(_09535_),
    .C(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__o32a_1 _37233_ (.A1(_08142_),
    .A2(_08137_),
    .A3(_08141_),
    .B1(_08153_),
    .B2(_08145_),
    .X(_09540_));
 sky130_fd_sc_hd__nand3b_2 _37234_ (.A_N(_24250_),
    .B(_24286_),
    .C(_22782_),
    .Y(_09541_));
 sky130_fd_sc_hd__o21ai_2 _37235_ (.A1(_20266_),
    .A2(_22094_),
    .B1(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__xor2_4 _37236_ (.A(_03564_),
    .B(_06586_),
    .X(_09543_));
 sky130_fd_sc_hd__a21oi_1 _37237_ (.A1(_02017_),
    .A2(_06607_),
    .B1(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__and3_1 _37238_ (.A(_09543_),
    .B(_06588_),
    .C(_02017_),
    .X(_09545_));
 sky130_fd_sc_hd__nor3_1 _37239_ (.A(_09542_),
    .B(_09544_),
    .C(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__o21a_1 _37240_ (.A1(_09544_),
    .A2(_09545_),
    .B1(_09542_),
    .X(_09548_));
 sky130_fd_sc_hd__nor2_1 _37241_ (.A(_09546_),
    .B(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__inv_2 _37242_ (.A(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__a31o_1 _37243_ (.A1(_09532_),
    .A2(_09539_),
    .A3(_09540_),
    .B1(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__a31o_1 _37244_ (.A1(_06614_),
    .A2(_08144_),
    .A3(_08143_),
    .B1(_08152_),
    .X(_09552_));
 sky130_fd_sc_hd__o21bai_1 _37245_ (.A1(_09530_),
    .A2(_09531_),
    .B1_N(_09537_),
    .Y(_09553_));
 sky130_fd_sc_hd__o211ai_2 _37246_ (.A1(_09115_),
    .A2(_08141_),
    .B1(_09534_),
    .C1(_09535_),
    .Y(_09554_));
 sky130_fd_sc_hd__and3_1 _37247_ (.A(_09552_),
    .B(_09553_),
    .C(_09554_),
    .X(_09555_));
 sky130_fd_sc_hd__a21oi_4 _37248_ (.A1(_08391_),
    .A2(_08191_),
    .B1(_08390_),
    .Y(_09556_));
 sky130_fd_sc_hd__inv_2 _37249_ (.A(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__nand3_1 _37250_ (.A(_09552_),
    .B(_09553_),
    .C(_09554_),
    .Y(_09559_));
 sky130_fd_sc_hd__nand3_2 _37251_ (.A(_09532_),
    .B(_09539_),
    .C(_09540_),
    .Y(_09560_));
 sky130_fd_sc_hd__a21o_1 _37252_ (.A1(_09559_),
    .A2(_09560_),
    .B1(_09549_),
    .X(_09561_));
 sky130_fd_sc_hd__o211ai_4 _37253_ (.A1(_09551_),
    .A2(_09555_),
    .B1(_09557_),
    .C1(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__nand2_1 _37254_ (.A(_09559_),
    .B(_09560_),
    .Y(_09563_));
 sky130_fd_sc_hd__nand2_1 _37255_ (.A(_09563_),
    .B(_09549_),
    .Y(_09564_));
 sky130_fd_sc_hd__nand3_2 _37256_ (.A(_09559_),
    .B(_09560_),
    .C(_09550_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand3_2 _37257_ (.A(_09564_),
    .B(_09556_),
    .C(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__a21o_1 _37258_ (.A1(_08156_),
    .A2(_08169_),
    .B1(_08177_),
    .X(_09567_));
 sky130_fd_sc_hd__a21oi_2 _37259_ (.A1(_09562_),
    .A2(_09566_),
    .B1(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__clkbuf_2 _37260_ (.A(_09568_),
    .X(_09570_));
 sky130_fd_sc_hd__or2b_1 _37261_ (.A(_08395_),
    .B_N(_08938_),
    .X(_09571_));
 sky130_fd_sc_hd__and2_1 _37262_ (.A(_09571_),
    .B(_08941_),
    .X(_09572_));
 sky130_fd_sc_hd__and3b_1 _37263_ (.A_N(_08351_),
    .B(_08376_),
    .C(_08352_),
    .X(_09573_));
 sky130_fd_sc_hd__a21o_2 _37264_ (.A1(_08318_),
    .A2(_08377_),
    .B1(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__or2b_1 _37265_ (.A(_08893_),
    .B_N(_08926_),
    .X(_09575_));
 sky130_fd_sc_hd__a21boi_4 _37266_ (.A1(_08885_),
    .A2(_08927_),
    .B1_N(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__nor2_1 _37267_ (.A(_06867_),
    .B(_06868_),
    .Y(_09577_));
 sky130_fd_sc_hd__nand2_1 _37268_ (.A(_06869_),
    .B(_06870_),
    .Y(_09578_));
 sky130_fd_sc_hd__and3_1 _37269_ (.A(_09577_),
    .B(_08374_),
    .C(_09578_),
    .X(_09579_));
 sky130_fd_sc_hd__a21oi_1 _37270_ (.A1(_06882_),
    .A2(_06874_),
    .B1(_08356_),
    .Y(_09581_));
 sky130_fd_sc_hd__buf_1 _37271_ (.A(_05196_),
    .X(_09582_));
 sky130_fd_sc_hd__o21ai_1 _37272_ (.A1(_03812_),
    .A2(_06847_),
    .B1(_05196_),
    .Y(_09583_));
 sky130_fd_sc_hd__o21ai_1 _37273_ (.A1(_09582_),
    .A2(_06846_),
    .B1(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__nand2_1 _37274_ (.A(_02805_),
    .B(_05207_),
    .Y(_09585_));
 sky130_fd_sc_hd__clkbuf_2 _37275_ (.A(_05204_),
    .X(_09586_));
 sky130_fd_sc_hd__nand2_1 _37276_ (.A(_09586_),
    .B(_01115_),
    .Y(_09587_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37277_ (.A(_02795_),
    .X(_09588_));
 sky130_fd_sc_hd__nand4_2 _37278_ (.A(_05211_),
    .B(_09585_),
    .C(_09587_),
    .D(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__a22o_1 _37279_ (.A1(_05211_),
    .A2(_09588_),
    .B1(_09585_),
    .B2(_09587_),
    .X(_09590_));
 sky130_fd_sc_hd__nand2_1 _37280_ (.A(_09589_),
    .B(_09590_),
    .Y(_09592_));
 sky130_fd_sc_hd__or2_1 _37281_ (.A(_09584_),
    .B(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__nand2_1 _37282_ (.A(_09584_),
    .B(_09592_),
    .Y(_09594_));
 sky130_fd_sc_hd__o21bai_1 _37283_ (.A1(_08359_),
    .A2(_08362_),
    .B1_N(_08363_),
    .Y(_09595_));
 sky130_fd_sc_hd__a21oi_1 _37284_ (.A1(_09593_),
    .A2(_09594_),
    .B1(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__and3_1 _37285_ (.A(_09595_),
    .B(_09593_),
    .C(_09594_),
    .X(_09597_));
 sky130_fd_sc_hd__nor4_1 _37286_ (.A(_24971_),
    .B(_08358_),
    .C(_09596_),
    .D(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__o32a_1 _37287_ (.A1(_21126_),
    .A2(_02805_),
    .A3(_08358_),
    .B1(_09596_),
    .B2(_09597_),
    .X(_09599_));
 sky130_fd_sc_hd__nor2_1 _37288_ (.A(net155),
    .B(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__a32oi_4 _37289_ (.A1(_08364_),
    .A2(_08365_),
    .A3(_08367_),
    .B1(_08370_),
    .B2(_06842_),
    .Y(_09601_));
 sky130_fd_sc_hd__xor2_1 _37290_ (.A(_09600_),
    .B(_09601_),
    .X(_09603_));
 sky130_fd_sc_hd__o21ai_1 _37291_ (.A1(_08375_),
    .A2(_09581_),
    .B1(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__a21o_1 _37292_ (.A1(_09577_),
    .A2(_09578_),
    .B1(_08374_),
    .X(_09605_));
 sky130_fd_sc_hd__a21oi_1 _37293_ (.A1(_08357_),
    .A2(_09605_),
    .B1(_09579_),
    .Y(_09606_));
 sky130_fd_sc_hd__o22a_1 _37294_ (.A1(_09579_),
    .A2(_09604_),
    .B1(_09603_),
    .B2(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__o21ai_1 _37295_ (.A1(_08372_),
    .A2(_08373_),
    .B1(_09607_),
    .Y(_09608_));
 sky130_fd_sc_hd__or3_1 _37296_ (.A(_08372_),
    .B(_08373_),
    .C(_09607_),
    .X(_09609_));
 sky130_fd_sc_hd__inv_2 _37297_ (.A(net309),
    .Y(_09610_));
 sky130_fd_sc_hd__nor2_1 _37298_ (.A(_08330_),
    .B(_08332_),
    .Y(_09611_));
 sky130_fd_sc_hd__nor2_1 _37299_ (.A(_03774_),
    .B(net311),
    .Y(_09612_));
 sky130_fd_sc_hd__and2_1 _37300_ (.A(_03774_),
    .B(net311),
    .X(_09614_));
 sky130_fd_sc_hd__or2_1 _37301_ (.A(_09612_),
    .B(_09614_),
    .X(_09615_));
 sky130_fd_sc_hd__o21ba_1 _37302_ (.A1(_09610_),
    .A2(_09611_),
    .B1_N(_09615_),
    .X(_09616_));
 sky130_fd_sc_hd__clkbuf_2 _37303_ (.A(net309),
    .X(_09617_));
 sky130_fd_sc_hd__o221a_1 _37304_ (.A1(_08330_),
    .A2(_08332_),
    .B1(_09612_),
    .B2(_09614_),
    .C1(_09617_),
    .X(_09618_));
 sky130_fd_sc_hd__clkbuf_2 _37305_ (.A(_03774_),
    .X(_09619_));
 sky130_fd_sc_hd__nand2_1 _37306_ (.A(_08320_),
    .B(_06817_),
    .Y(_09620_));
 sky130_fd_sc_hd__a21o_1 _37307_ (.A1(_02838_),
    .A2(_06817_),
    .B1(_05252_),
    .X(_09621_));
 sky130_fd_sc_hd__o21ai_1 _37308_ (.A1(_09619_),
    .A2(_09620_),
    .B1(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__a21o_1 _37309_ (.A1(_23357_),
    .A2(_08321_),
    .B1(_09622_),
    .X(_09623_));
 sky130_fd_sc_hd__or3b_1 _37310_ (.A(_05237_),
    .B(_06812_),
    .C_N(_09622_),
    .X(_09625_));
 sky130_fd_sc_hd__o211a_1 _37311_ (.A1(_09616_),
    .A2(_09618_),
    .B1(_09623_),
    .C1(_09625_),
    .X(_09626_));
 sky130_fd_sc_hd__a211oi_1 _37312_ (.A1(_09623_),
    .A2(_09625_),
    .B1(_09616_),
    .C1(_09618_),
    .Y(_09627_));
 sky130_fd_sc_hd__nand4_1 _37313_ (.A(_08328_),
    .B(_08329_),
    .C(_08333_),
    .D(_08334_),
    .Y(_09628_));
 sky130_fd_sc_hd__o31a_1 _37314_ (.A1(_09610_),
    .A2(_06818_),
    .A3(_09611_),
    .B1(_09628_),
    .X(_09629_));
 sky130_fd_sc_hd__o21ai_1 _37315_ (.A1(_09626_),
    .A2(_09627_),
    .B1(_09629_),
    .Y(_09630_));
 sky130_fd_sc_hd__or3_1 _37316_ (.A(_09629_),
    .B(_09626_),
    .C(_09627_),
    .X(_09631_));
 sky130_fd_sc_hd__and2_1 _37317_ (.A(_09630_),
    .B(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__clkbuf_2 _37318_ (.A(_06817_),
    .X(_09633_));
 sky130_fd_sc_hd__a31o_1 _37319_ (.A1(_05237_),
    .A2(_08322_),
    .A3(_09633_),
    .B1(net249),
    .X(_09634_));
 sky130_fd_sc_hd__nand2_1 _37320_ (.A(_09632_),
    .B(_09634_),
    .Y(_09636_));
 sky130_fd_sc_hd__a311o_1 _37321_ (.A1(_05237_),
    .A2(_08322_),
    .A3(_09633_),
    .B1(net249),
    .C1(_09632_),
    .X(_09637_));
 sky130_fd_sc_hd__a21bo_1 _37322_ (.A1(_08323_),
    .A2(_08339_),
    .B1_N(_08340_),
    .X(_09638_));
 sky130_fd_sc_hd__and3_1 _37323_ (.A(_09636_),
    .B(_09637_),
    .C(_09638_),
    .X(_09639_));
 sky130_fd_sc_hd__a21oi_1 _37324_ (.A1(_09636_),
    .A2(_09637_),
    .B1(_09638_),
    .Y(_09640_));
 sky130_fd_sc_hd__nor2_1 _37325_ (.A(_09639_),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__and3_1 _37326_ (.A(_09641_),
    .B(_08319_),
    .C(_08343_),
    .X(_09642_));
 sky130_fd_sc_hd__o2bb2a_1 _37327_ (.A1_N(_08343_),
    .A2_N(_08319_),
    .B1(_09640_),
    .B2(_09639_),
    .X(_09643_));
 sky130_fd_sc_hd__or2_1 _37328_ (.A(_09642_),
    .B(_09643_),
    .X(_09644_));
 sky130_fd_sc_hd__o21ba_1 _37329_ (.A1(_08345_),
    .A2(_08351_),
    .B1_N(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__or3b_1 _37330_ (.A(_08345_),
    .B(_08351_),
    .C_N(_09644_),
    .X(_09647_));
 sky130_fd_sc_hd__or2b_1 _37331_ (.A(_09645_),
    .B_N(_09647_),
    .X(_09648_));
 sky130_fd_sc_hd__a21oi_2 _37332_ (.A1(_09608_),
    .A2(_09609_),
    .B1(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21bo_1 _37333_ (.A1(_08284_),
    .A2(_06786_),
    .B1_N(_05160_),
    .X(_09650_));
 sky130_fd_sc_hd__or3b_1 _37334_ (.A(_08290_),
    .B(_05160_),
    .C_N(_08284_),
    .X(_09651_));
 sky130_fd_sc_hd__o2bb2a_1 _37335_ (.A1_N(_08291_),
    .A2_N(_06779_),
    .B1(_08290_),
    .B2(_08296_),
    .X(_09652_));
 sky130_fd_sc_hd__a21oi_1 _37336_ (.A1(_08292_),
    .A2(_08299_),
    .B1(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__o31a_1 _37337_ (.A1(_08288_),
    .A2(_08289_),
    .A3(_08297_),
    .B1(_09652_),
    .X(_09654_));
 sky130_fd_sc_hd__o2bb2a_1 _37338_ (.A1_N(_09650_),
    .A2_N(_09651_),
    .B1(_09653_),
    .B2(_09654_),
    .X(_09655_));
 sky130_fd_sc_hd__inv_2 _37339_ (.A(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__nand2_1 _37340_ (.A(_09650_),
    .B(_09651_),
    .Y(_09658_));
 sky130_fd_sc_hd__or3_1 _37341_ (.A(_09654_),
    .B(_09658_),
    .C(_09653_),
    .X(_09659_));
 sky130_fd_sc_hd__a32o_1 _37342_ (.A1(_08298_),
    .A2(_08299_),
    .A3(_08300_),
    .B1(_08303_),
    .B2(_08306_),
    .X(_09660_));
 sky130_fd_sc_hd__and3_1 _37343_ (.A(_09656_),
    .B(_09659_),
    .C(_09660_),
    .X(_09661_));
 sky130_fd_sc_hd__a21o_1 _37344_ (.A1(_09656_),
    .A2(_09659_),
    .B1(_09660_),
    .X(_09662_));
 sky130_fd_sc_hd__and2b_1 _37345_ (.A_N(_09661_),
    .B(_09662_),
    .X(_09663_));
 sky130_fd_sc_hd__xor2_1 _37346_ (.A(_08285_),
    .B(_09663_),
    .X(_09664_));
 sky130_fd_sc_hd__a211oi_1 _37347_ (.A1(_06772_),
    .A2(_08311_),
    .B1(_09664_),
    .C1(_08308_),
    .Y(_09665_));
 sky130_fd_sc_hd__o21a_1 _37348_ (.A1(_08308_),
    .A2(_08312_),
    .B1(_09664_),
    .X(_09666_));
 sky130_fd_sc_hd__or2_1 _37349_ (.A(_09665_),
    .B(_09666_),
    .X(_09667_));
 sky130_fd_sc_hd__nand2_1 _37350_ (.A(_08313_),
    .B(_09667_),
    .Y(_09669_));
 sky130_fd_sc_hd__inv_2 _37351_ (.A(_08313_),
    .Y(_09670_));
 sky130_fd_sc_hd__o21ba_1 _37352_ (.A1(_09670_),
    .A2(_08315_),
    .B1_N(_09667_),
    .X(_09671_));
 sky130_fd_sc_hd__o21bai_1 _37353_ (.A1(_08315_),
    .A2(_09669_),
    .B1_N(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__and3_1 _37354_ (.A(_09608_),
    .B(_09609_),
    .C(_09648_),
    .X(_09673_));
 sky130_fd_sc_hd__nor3_1 _37355_ (.A(_09649_),
    .B(_09672_),
    .C(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__o21ai_1 _37356_ (.A1(_09673_),
    .A2(_09649_),
    .B1(_09672_),
    .Y(_09675_));
 sky130_fd_sc_hd__inv_2 _37357_ (.A(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__nor3_1 _37358_ (.A(_09576_),
    .B(_09674_),
    .C(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__o21ai_1 _37359_ (.A1(_09674_),
    .A2(_09676_),
    .B1(_09576_),
    .Y(_09678_));
 sky130_fd_sc_hd__and2b_1 _37360_ (.A_N(_09677_),
    .B(_09678_),
    .X(_09680_));
 sky130_fd_sc_hd__xnor2_4 _37361_ (.A(_09574_),
    .B(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__nand2_1 _37362_ (.A(_08378_),
    .B(_08280_),
    .Y(_09682_));
 sky130_fd_sc_hd__o21a_2 _37363_ (.A1(_08380_),
    .A2(_08379_),
    .B1(_09682_),
    .X(_09683_));
 sky130_fd_sc_hd__nand2_1 _37364_ (.A(_09681_),
    .B(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__or2_1 _37365_ (.A(_09683_),
    .B(_09681_),
    .X(_09685_));
 sky130_fd_sc_hd__a21o_2 _37366_ (.A1(_08237_),
    .A2(_08232_),
    .B1(_08231_),
    .X(_09686_));
 sky130_fd_sc_hd__nor2b_1 _37367_ (.A(_06670_),
    .B_N(net295),
    .Y(_09687_));
 sky130_fd_sc_hd__and2b_1 _37368_ (.A_N(net295),
    .B(_06670_),
    .X(_09688_));
 sky130_fd_sc_hd__nor2_1 _37369_ (.A(_09687_),
    .B(_09688_),
    .Y(_09689_));
 sky130_fd_sc_hd__inv_2 _37370_ (.A(\delay_line[36][13] ),
    .Y(_09691_));
 sky130_fd_sc_hd__nand2_1 _37371_ (.A(_08240_),
    .B(_08242_),
    .Y(_09692_));
 sky130_fd_sc_hd__o21ai_1 _37372_ (.A1(_06669_),
    .A2(_09691_),
    .B1(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__xor2_1 _37373_ (.A(_09689_),
    .B(_09693_),
    .X(_09694_));
 sky130_fd_sc_hd__a2bb2o_1 _37374_ (.A1_N(_08245_),
    .A2_N(_08246_),
    .B1(\delay_line[36][13] ),
    .B2(_08241_),
    .X(_09695_));
 sky130_fd_sc_hd__xor2_1 _37375_ (.A(_09694_),
    .B(_09695_),
    .X(_09696_));
 sky130_fd_sc_hd__nand2_1 _37376_ (.A(_08253_),
    .B(_03702_),
    .Y(_09697_));
 sky130_fd_sc_hd__or2_1 _37377_ (.A(_03702_),
    .B(_08253_),
    .X(_09698_));
 sky130_fd_sc_hd__and4bb_1 _37378_ (.A_N(_08248_),
    .B_N(_08249_),
    .C(_08251_),
    .D(_05319_),
    .X(_09699_));
 sky130_fd_sc_hd__a211oi_1 _37379_ (.A1(_09697_),
    .A2(_09698_),
    .B1(_09699_),
    .C1(_08257_),
    .Y(_09700_));
 sky130_fd_sc_hd__o211a_1 _37380_ (.A1(_09699_),
    .A2(_08257_),
    .B1(_09697_),
    .C1(_09698_),
    .X(_09702_));
 sky130_fd_sc_hd__or4_1 _37381_ (.A(_08262_),
    .B(_08265_),
    .C(_09700_),
    .D(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__o22ai_1 _37382_ (.A1(_08262_),
    .A2(_08265_),
    .B1(_09700_),
    .B2(_09702_),
    .Y(_09704_));
 sky130_fd_sc_hd__nand2_1 _37383_ (.A(_09703_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__or2_1 _37384_ (.A(_09696_),
    .B(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__nand2_1 _37385_ (.A(_09705_),
    .B(_09696_),
    .Y(_09707_));
 sky130_fd_sc_hd__nand2_1 _37386_ (.A(_09706_),
    .B(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__xor2_2 _37387_ (.A(_09686_),
    .B(_09708_),
    .X(_09709_));
 sky130_fd_sc_hd__o22a_1 _37388_ (.A1(_08247_),
    .A2(_08266_),
    .B1(_08269_),
    .B2(_08238_),
    .X(_09710_));
 sky130_fd_sc_hd__nand2_1 _37389_ (.A(_09709_),
    .B(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__a21o_1 _37390_ (.A1(_08267_),
    .A2(_08270_),
    .B1(_09709_),
    .X(_09713_));
 sky130_fd_sc_hd__a21bo_1 _37391_ (.A1(_03663_),
    .A2(_08193_),
    .B1_N(_08192_),
    .X(_09714_));
 sky130_fd_sc_hd__xnor2_4 _37392_ (.A(_05342_),
    .B(_09714_),
    .Y(_09715_));
 sky130_fd_sc_hd__a211oi_1 _37393_ (.A1(_06758_),
    .A2(_08197_),
    .B1(_08194_),
    .C1(_08196_),
    .Y(_09716_));
 sky130_fd_sc_hd__a21oi_2 _37394_ (.A1(_08198_),
    .A2(_08200_),
    .B1(_09716_),
    .Y(_09717_));
 sky130_fd_sc_hd__xor2_4 _37395_ (.A(_09715_),
    .B(_09717_),
    .X(_09718_));
 sky130_fd_sc_hd__nand2_1 _37396_ (.A(_05383_),
    .B(_06719_),
    .Y(_09719_));
 sky130_fd_sc_hd__o21a_1 _37397_ (.A1(_08205_),
    .A2(_09719_),
    .B1(_08213_),
    .X(_09720_));
 sky130_fd_sc_hd__buf_2 _37398_ (.A(\delay_line[38][15] ),
    .X(_09721_));
 sky130_fd_sc_hd__or3b_1 _37399_ (.A(_08204_),
    .B(_06717_),
    .C_N(_09721_),
    .X(_09722_));
 sky130_fd_sc_hd__nand2_1 _37400_ (.A(_09722_),
    .B(_05379_),
    .Y(_09724_));
 sky130_fd_sc_hd__or4b_1 _37401_ (.A(_08204_),
    .B(_06717_),
    .C(_05379_),
    .D_N(_09721_),
    .X(_09725_));
 sky130_fd_sc_hd__and3_1 _37402_ (.A(_09720_),
    .B(_09724_),
    .C(_09725_),
    .X(_09726_));
 sky130_fd_sc_hd__a21oi_1 _37403_ (.A1(_09725_),
    .A2(_09724_),
    .B1(_09720_),
    .Y(_09727_));
 sky130_fd_sc_hd__or2_2 _37404_ (.A(_09726_),
    .B(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__mux2_1 _37405_ (.A0(_05364_),
    .A1(_05363_),
    .S(_08215_),
    .X(_09729_));
 sky130_fd_sc_hd__o21ai_1 _37406_ (.A1(_06732_),
    .A2(_06737_),
    .B1(_08214_),
    .Y(_09730_));
 sky130_fd_sc_hd__o31a_1 _37407_ (.A1(_06732_),
    .A2(_06737_),
    .A3(_09729_),
    .B1(_09730_),
    .X(_09731_));
 sky130_fd_sc_hd__or3_1 _37408_ (.A(_08214_),
    .B(_06732_),
    .C(_06737_),
    .X(_09732_));
 sky130_fd_sc_hd__a211oi_1 _37409_ (.A1(_09730_),
    .A2(_09732_),
    .B1(_09729_),
    .C1(_08220_),
    .Y(_09733_));
 sky130_fd_sc_hd__a21o_2 _37410_ (.A1(_08221_),
    .A2(_09731_),
    .B1(_09733_),
    .X(_09735_));
 sky130_fd_sc_hd__xor2_2 _37411_ (.A(_09728_),
    .B(_09735_),
    .X(_09736_));
 sky130_fd_sc_hd__xnor2_4 _37412_ (.A(_09718_),
    .B(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__a21oi_1 _37413_ (.A1(_09711_),
    .A2(_09713_),
    .B1(_09737_),
    .Y(_09738_));
 sky130_fd_sc_hd__and3_1 _37414_ (.A(_09737_),
    .B(_09711_),
    .C(_09713_),
    .X(_09739_));
 sky130_fd_sc_hd__nor2_2 _37415_ (.A(_09738_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__a21oi_1 _37416_ (.A1(_09684_),
    .A2(_09685_),
    .B1(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__and2_1 _37417_ (.A(_09681_),
    .B(_09683_),
    .X(_09742_));
 sky130_fd_sc_hd__and3b_1 _37418_ (.A_N(_09742_),
    .B(_09685_),
    .C(_09740_),
    .X(_09743_));
 sky130_fd_sc_hd__a21oi_1 _37419_ (.A1(_08935_),
    .A2(_08777_),
    .B1(_08933_),
    .Y(_09744_));
 sky130_fd_sc_hd__o21a_1 _37420_ (.A1(_09741_),
    .A2(_09743_),
    .B1(_09744_),
    .X(_09746_));
 sky130_fd_sc_hd__inv_2 _37421_ (.A(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__or3_2 _37422_ (.A(_09744_),
    .B(_09741_),
    .C(_09743_),
    .X(_09748_));
 sky130_fd_sc_hd__and2_1 _37423_ (.A(_08384_),
    .B(_08386_),
    .X(_09749_));
 sky130_fd_sc_hd__a21boi_1 _37424_ (.A1(_09747_),
    .A2(_09748_),
    .B1_N(_09749_),
    .Y(_09750_));
 sky130_fd_sc_hd__nor3b_2 _37425_ (.A(_09749_),
    .B(_09746_),
    .C_N(_09748_),
    .Y(_09751_));
 sky130_fd_sc_hd__o21bai_4 _37426_ (.A1(_08764_),
    .A2(_08640_),
    .B1_N(_08639_),
    .Y(_09752_));
 sky130_fd_sc_hd__buf_1 _37427_ (.A(_08687_),
    .X(_09753_));
 sky130_fd_sc_hd__and3b_1 _37428_ (.A_N(_09753_),
    .B(_07394_),
    .C(_21354_),
    .X(_09754_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37429_ (.A(_22931_),
    .X(_09755_));
 sky130_fd_sc_hd__o21ai_2 _37430_ (.A1(_09755_),
    .A2(_07376_),
    .B1(_08687_),
    .Y(_09757_));
 sky130_fd_sc_hd__buf_1 _37431_ (.A(net372),
    .X(_09758_));
 sky130_fd_sc_hd__nand2_1 _37432_ (.A(_04013_),
    .B(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__inv_2 _37433_ (.A(\delay_line[18][12] ),
    .Y(_09760_));
 sky130_fd_sc_hd__inv_2 _37434_ (.A(\delay_line[18][15] ),
    .Y(_09761_));
 sky130_fd_sc_hd__nand2_1 _37435_ (.A(_09760_),
    .B(_09761_),
    .Y(_09762_));
 sky130_fd_sc_hd__a22o_1 _37436_ (.A1(_02635_),
    .A2(_09758_),
    .B1(_09759_),
    .B2(_09762_),
    .X(_09763_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37437_ (.A(_04013_),
    .X(_09764_));
 sky130_fd_sc_hd__or3b_1 _37438_ (.A(_09764_),
    .B(_09761_),
    .C_N(_02635_),
    .X(_09765_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37439_ (.A(_08691_),
    .X(_09766_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37440_ (.A(\delay_line[18][9] ),
    .X(_09768_));
 sky130_fd_sc_hd__or2_1 _37441_ (.A(_21363_),
    .B(_09768_),
    .X(_09769_));
 sky130_fd_sc_hd__o21ai_1 _37442_ (.A1(_07378_),
    .A2(_09766_),
    .B1(_09768_),
    .Y(_09770_));
 sky130_fd_sc_hd__o21a_1 _37443_ (.A1(_09766_),
    .A2(_09769_),
    .B1(_09770_),
    .X(_09771_));
 sky130_fd_sc_hd__a21oi_1 _37444_ (.A1(_09763_),
    .A2(_09765_),
    .B1(_09771_),
    .Y(_09772_));
 sky130_fd_sc_hd__and3_1 _37445_ (.A(_09771_),
    .B(_09763_),
    .C(_09765_),
    .X(_09773_));
 sky130_fd_sc_hd__nand2_1 _37446_ (.A(_08696_),
    .B(_08698_),
    .Y(_09774_));
 sky130_fd_sc_hd__or3_1 _37447_ (.A(_09772_),
    .B(_09773_),
    .C(_09774_),
    .X(_09775_));
 sky130_fd_sc_hd__o21ai_1 _37448_ (.A1(_09772_),
    .A2(_09773_),
    .B1(_09774_),
    .Y(_09776_));
 sky130_fd_sc_hd__nand2_1 _37449_ (.A(_09775_),
    .B(_09776_),
    .Y(_09777_));
 sky130_fd_sc_hd__xor2_2 _37450_ (.A(_09757_),
    .B(_09777_),
    .X(_09779_));
 sky130_fd_sc_hd__o211a_1 _37451_ (.A1(_08687_),
    .A2(_07375_),
    .B1(_07394_),
    .C1(_08704_),
    .X(_09780_));
 sky130_fd_sc_hd__a31o_1 _37452_ (.A1(_08700_),
    .A2(_08698_),
    .A3(_08699_),
    .B1(_09780_),
    .X(_09781_));
 sky130_fd_sc_hd__nor2_1 _37453_ (.A(_09779_),
    .B(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__o21ai_1 _37454_ (.A1(_08703_),
    .A2(_09780_),
    .B1(_09779_),
    .Y(_09783_));
 sky130_fd_sc_hd__and2b_1 _37455_ (.A_N(_09782_),
    .B(_09783_),
    .X(_09784_));
 sky130_fd_sc_hd__nor2_2 _37456_ (.A(_09754_),
    .B(_09784_),
    .Y(_09785_));
 sky130_fd_sc_hd__o41a_1 _37457_ (.A1(_18389_),
    .A2(_07375_),
    .A3(_07394_),
    .A4(_08706_),
    .B1(_08707_),
    .X(_09786_));
 sky130_fd_sc_hd__a21o_1 _37458_ (.A1(_09754_),
    .A2(_09784_),
    .B1(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__o211a_1 _37459_ (.A1(_08703_),
    .A2(_09779_),
    .B1(_09754_),
    .C1(_09783_),
    .X(_09788_));
 sky130_fd_sc_hd__o21ai_1 _37460_ (.A1(_09785_),
    .A2(_09788_),
    .B1(_09786_),
    .Y(_09790_));
 sky130_fd_sc_hd__o21ai_4 _37461_ (.A1(_09785_),
    .A2(_09787_),
    .B1(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__and2b_1 _37462_ (.A_N(_08710_),
    .B(_08709_),
    .X(_09792_));
 sky130_fd_sc_hd__a21oi_4 _37463_ (.A1(_08715_),
    .A2(_08711_),
    .B1(_09792_),
    .Y(_09793_));
 sky130_fd_sc_hd__xnor2_4 _37464_ (.A(_09791_),
    .B(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__o21ai_1 _37465_ (.A1(_20574_),
    .A2(_08719_),
    .B1(_07406_),
    .Y(_09795_));
 sky130_fd_sc_hd__o32a_1 _37466_ (.A1(_07408_),
    .A2(_09795_),
    .A3(_08752_),
    .B1(_08751_),
    .B2(_08721_),
    .X(_09796_));
 sky130_fd_sc_hd__clkbuf_2 _37467_ (.A(_08735_),
    .X(_09797_));
 sky130_fd_sc_hd__nand2_2 _37468_ (.A(_07418_),
    .B(_07416_),
    .Y(_09798_));
 sky130_fd_sc_hd__buf_1 _37469_ (.A(_02586_),
    .X(_09799_));
 sky130_fd_sc_hd__a21oi_2 _37470_ (.A1(_07416_),
    .A2(_09797_),
    .B1(_09799_),
    .Y(_09801_));
 sky130_fd_sc_hd__and3_1 _37471_ (.A(_02586_),
    .B(_07416_),
    .C(_08735_),
    .X(_09802_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37472_ (.A(_00662_),
    .X(_09803_));
 sky130_fd_sc_hd__o211ai_2 _37473_ (.A1(_08735_),
    .A2(_09798_),
    .B1(_09803_),
    .C1(_08736_),
    .Y(_09804_));
 sky130_fd_sc_hd__o221ai_4 _37474_ (.A1(_09797_),
    .A2(_09798_),
    .B1(_09801_),
    .B2(_09802_),
    .C1(_09804_),
    .Y(_09805_));
 sky130_fd_sc_hd__a211o_1 _37475_ (.A1(_08737_),
    .A2(_09804_),
    .B1(_09801_),
    .C1(_09802_),
    .X(_09806_));
 sky130_fd_sc_hd__nor2_1 _37476_ (.A(_00653_),
    .B(_00654_),
    .Y(_09807_));
 sky130_fd_sc_hd__a21oi_1 _37477_ (.A1(_24661_),
    .A2(_21382_),
    .B1(_07433_),
    .Y(_09808_));
 sky130_fd_sc_hd__and3_1 _37478_ (.A(_00663_),
    .B(_00659_),
    .C(_09808_),
    .X(_09809_));
 sky130_fd_sc_hd__o21ba_1 _37479_ (.A1(_09807_),
    .A2(_09808_),
    .B1_N(_09809_),
    .X(_09810_));
 sky130_fd_sc_hd__and3_1 _37480_ (.A(_09805_),
    .B(_09806_),
    .C(_09810_),
    .X(_09812_));
 sky130_fd_sc_hd__a21oi_1 _37481_ (.A1(_09805_),
    .A2(_09806_),
    .B1(_09810_),
    .Y(_09813_));
 sky130_fd_sc_hd__a211oi_1 _37482_ (.A1(_08741_),
    .A2(_08731_),
    .B1(_08738_),
    .C1(_08739_),
    .Y(_09814_));
 sky130_fd_sc_hd__nor2_1 _37483_ (.A(_09814_),
    .B(_08743_),
    .Y(_09815_));
 sky130_fd_sc_hd__o21ai_1 _37484_ (.A1(_09812_),
    .A2(_09813_),
    .B1(_09815_),
    .Y(_09816_));
 sky130_fd_sc_hd__or3_1 _37485_ (.A(_09815_),
    .B(_09812_),
    .C(_09813_),
    .X(_09817_));
 sky130_fd_sc_hd__o21a_1 _37486_ (.A1(_07409_),
    .A2(_07433_),
    .B1(_24658_),
    .X(_09818_));
 sky130_fd_sc_hd__nor2_1 _37487_ (.A(_24656_),
    .B(_24657_),
    .Y(_09819_));
 sky130_fd_sc_hd__o22a_1 _37488_ (.A1(_04055_),
    .A2(_07432_),
    .B1(_09818_),
    .B2(_09819_),
    .X(_09820_));
 sky130_fd_sc_hd__a21o_1 _37489_ (.A1(_09816_),
    .A2(_09817_),
    .B1(_09820_),
    .X(_09821_));
 sky130_fd_sc_hd__nand3_1 _37490_ (.A(_09817_),
    .B(_09820_),
    .C(_09816_),
    .Y(_09823_));
 sky130_fd_sc_hd__o21ai_1 _37491_ (.A1(_08743_),
    .A2(_08744_),
    .B1(_08747_),
    .Y(_09824_));
 sky130_fd_sc_hd__a21o_1 _37492_ (.A1(_09824_),
    .A2(_08724_),
    .B1(_08748_),
    .X(_09825_));
 sky130_fd_sc_hd__and3_1 _37493_ (.A(_09821_),
    .B(_09823_),
    .C(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__o22a_1 _37494_ (.A1(_07406_),
    .A2(_04055_),
    .B1(_07433_),
    .B2(_07431_),
    .X(_09827_));
 sky130_fd_sc_hd__a21o_1 _37495_ (.A1(_09821_),
    .A2(_09823_),
    .B1(_09825_),
    .X(_09828_));
 sky130_fd_sc_hd__and4b_1 _37496_ (.A_N(_09826_),
    .B(_09827_),
    .C(_08719_),
    .D(_09828_),
    .X(_09829_));
 sky130_fd_sc_hd__inv_2 _37497_ (.A(_09828_),
    .Y(_09830_));
 sky130_fd_sc_hd__o2bb2a_1 _37498_ (.A1_N(_08719_),
    .A2_N(_09827_),
    .B1(_09830_),
    .B2(_09826_),
    .X(_09831_));
 sky130_fd_sc_hd__or2_1 _37499_ (.A(_09829_),
    .B(_09831_),
    .X(_09832_));
 sky130_fd_sc_hd__nor2_1 _37500_ (.A(_09796_),
    .B(_09832_),
    .Y(_09834_));
 sky130_fd_sc_hd__nand2_1 _37501_ (.A(_09832_),
    .B(_09796_),
    .Y(_09835_));
 sky130_fd_sc_hd__or2b_1 _37502_ (.A(_09834_),
    .B_N(_09835_),
    .X(_09836_));
 sky130_fd_sc_hd__and2b_1 _37503_ (.A_N(_08754_),
    .B(_09836_),
    .X(_09837_));
 sky130_fd_sc_hd__o21bai_1 _37504_ (.A1(_07454_),
    .A2(_07455_),
    .B1_N(_07453_),
    .Y(_09838_));
 sky130_fd_sc_hd__a21oi_1 _37505_ (.A1(_09838_),
    .A2(_08757_),
    .B1(_08754_),
    .Y(_09839_));
 sky130_fd_sc_hd__nor2_1 _37506_ (.A(_09836_),
    .B(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__a21o_2 _37507_ (.A1(_09837_),
    .A2(_08761_),
    .B1(_09840_),
    .X(_09841_));
 sky130_fd_sc_hd__xor2_4 _37508_ (.A(_09794_),
    .B(_09841_),
    .X(_09842_));
 sky130_fd_sc_hd__inv_2 _37509_ (.A(_08676_),
    .Y(_09843_));
 sky130_fd_sc_hd__clkbuf_2 _37510_ (.A(_08656_),
    .X(_09845_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37511_ (.A(_04106_),
    .X(_09846_));
 sky130_fd_sc_hd__a21oi_2 _37512_ (.A1(_08652_),
    .A2(_09845_),
    .B1(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__and3_1 _37513_ (.A(_04106_),
    .B(_08652_),
    .C(_08656_),
    .X(_09848_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37514_ (.A(_02550_),
    .X(_09849_));
 sky130_fd_sc_hd__o211ai_2 _37515_ (.A1(_08656_),
    .A2(_08659_),
    .B1(_09849_),
    .C1(_08658_),
    .Y(_09850_));
 sky130_fd_sc_hd__o221ai_4 _37516_ (.A1(_09845_),
    .A2(_08659_),
    .B1(_09847_),
    .B2(_09848_),
    .C1(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__a211o_2 _37517_ (.A1(_08660_),
    .A2(_09850_),
    .B1(_09847_),
    .C1(_09848_),
    .X(_09852_));
 sky130_fd_sc_hd__clkbuf_2 _37518_ (.A(_00615_),
    .X(_09853_));
 sky130_fd_sc_hd__nor2_1 _37519_ (.A(_00614_),
    .B(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__mux2_1 _37520_ (.A0(_22992_),
    .A1(_24635_),
    .S(_21418_),
    .X(_09856_));
 sky130_fd_sc_hd__and3_1 _37521_ (.A(_00617_),
    .B(_09856_),
    .C(_00618_),
    .X(_09857_));
 sky130_fd_sc_hd__o21ba_1 _37522_ (.A1(_09854_),
    .A2(_09856_),
    .B1_N(_09857_),
    .X(_09858_));
 sky130_fd_sc_hd__nand3_4 _37523_ (.A(_09851_),
    .B(_09852_),
    .C(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__a21o_1 _37524_ (.A1(_09851_),
    .A2(_09852_),
    .B1(_09858_),
    .X(_09860_));
 sky130_fd_sc_hd__inv_2 _37525_ (.A(_08663_),
    .Y(_09861_));
 sky130_fd_sc_hd__a211o_1 _37526_ (.A1(_09859_),
    .A2(_09860_),
    .B1(_09861_),
    .C1(_08666_),
    .X(_09862_));
 sky130_fd_sc_hd__o211ai_4 _37527_ (.A1(_09861_),
    .A2(_08666_),
    .B1(_09859_),
    .C1(_09860_),
    .Y(_09863_));
 sky130_fd_sc_hd__or2_1 _37528_ (.A(_08644_),
    .B(_08645_),
    .X(_09864_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37529_ (.A(_05609_),
    .X(_09865_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37530_ (.A(_04098_),
    .X(_09867_));
 sky130_fd_sc_hd__a21oi_1 _37531_ (.A1(_07324_),
    .A2(_09865_),
    .B1(_09867_),
    .Y(_09868_));
 sky130_fd_sc_hd__a21oi_1 _37532_ (.A1(_09864_),
    .A2(_08649_),
    .B1(_09868_),
    .Y(_09869_));
 sky130_fd_sc_hd__a21oi_1 _37533_ (.A1(_09862_),
    .A2(_09863_),
    .B1(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__inv_2 _37534_ (.A(_09870_),
    .Y(_09871_));
 sky130_fd_sc_hd__nand3_1 _37535_ (.A(_09863_),
    .B(_09869_),
    .C(_09862_),
    .Y(_09872_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37536_ (.A(_09872_),
    .X(_09873_));
 sky130_fd_sc_hd__o221a_1 _37537_ (.A1(_07348_),
    .A2(_08669_),
    .B1(_08665_),
    .B2(_08667_),
    .C1(_07353_),
    .X(_09874_));
 sky130_fd_sc_hd__o32a_1 _37538_ (.A1(_08670_),
    .A2(_08666_),
    .A3(_08667_),
    .B1(_08643_),
    .B2(_09874_),
    .X(_09875_));
 sky130_fd_sc_hd__inv_2 _37539_ (.A(_09875_),
    .Y(_09876_));
 sky130_fd_sc_hd__a21oi_1 _37540_ (.A1(_09871_),
    .A2(_09873_),
    .B1(_09876_),
    .Y(_09878_));
 sky130_fd_sc_hd__and3_1 _37541_ (.A(_09871_),
    .B(_09872_),
    .C(_09876_),
    .X(_09879_));
 sky130_fd_sc_hd__nor2_1 _37542_ (.A(_09878_),
    .B(_09879_),
    .Y(_09880_));
 sky130_fd_sc_hd__o221a_2 _37543_ (.A1(_20513_),
    .A2(_05614_),
    .B1(_07340_),
    .B2(_07341_),
    .C1(_09880_),
    .X(_09881_));
 sky130_fd_sc_hd__o221a_1 _37544_ (.A1(_05598_),
    .A2(_09867_),
    .B1(_07340_),
    .B2(_07341_),
    .C1(_07324_),
    .X(_09882_));
 sky130_fd_sc_hd__nor2_1 _37545_ (.A(_09882_),
    .B(_09880_),
    .Y(_09883_));
 sky130_fd_sc_hd__nor2_1 _37546_ (.A(_09881_),
    .B(_09883_),
    .Y(_09884_));
 sky130_fd_sc_hd__o21a_1 _37547_ (.A1(_09843_),
    .A2(_08678_),
    .B1(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__a211oi_1 _37548_ (.A1(_08677_),
    .A2(_08675_),
    .B1(_09843_),
    .C1(_09884_),
    .Y(_09886_));
 sky130_fd_sc_hd__or2_1 _37549_ (.A(_09885_),
    .B(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__a21oi_1 _37550_ (.A1(_08683_),
    .A2(_08685_),
    .B1(_08682_),
    .Y(_09889_));
 sky130_fd_sc_hd__nor2_1 _37551_ (.A(_09887_),
    .B(_09889_),
    .Y(_09890_));
 sky130_fd_sc_hd__nor2_1 _37552_ (.A(_09885_),
    .B(_09886_),
    .Y(_09891_));
 sky130_fd_sc_hd__a21o_1 _37553_ (.A1(_08683_),
    .A2(_08685_),
    .B1(_08682_),
    .X(_09892_));
 sky130_fd_sc_hd__nor2_1 _37554_ (.A(_09891_),
    .B(_09892_),
    .Y(_09893_));
 sky130_fd_sc_hd__or2_2 _37555_ (.A(_09890_),
    .B(_09893_),
    .X(_09894_));
 sky130_fd_sc_hd__xor2_4 _37556_ (.A(_09842_),
    .B(_09894_),
    .X(_09895_));
 sky130_fd_sc_hd__a21oi_2 _37557_ (.A1(_08585_),
    .A2(_08586_),
    .B1(_08589_),
    .Y(_09896_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37558_ (.A(\delay_line[14][11] ),
    .X(_09897_));
 sky130_fd_sc_hd__a21oi_1 _37559_ (.A1(_08570_),
    .A2(_09897_),
    .B1(_07285_),
    .Y(_09898_));
 sky130_fd_sc_hd__and3_1 _37560_ (.A(_07285_),
    .B(_02405_),
    .C(_09897_),
    .X(_09900_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37561_ (.A(_08572_),
    .X(_09901_));
 sky130_fd_sc_hd__xor2_1 _37562_ (.A(_09897_),
    .B(\delay_line[14][12] ),
    .X(_09902_));
 sky130_fd_sc_hd__o21ai_1 _37563_ (.A1(_09901_),
    .A2(_08573_),
    .B1(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__or3_1 _37564_ (.A(_08572_),
    .B(_08573_),
    .C(_09902_),
    .X(_09904_));
 sky130_fd_sc_hd__o211a_1 _37565_ (.A1(_09898_),
    .A2(_09900_),
    .B1(_09903_),
    .C1(_09904_),
    .X(_09905_));
 sky130_fd_sc_hd__a211oi_2 _37566_ (.A1(_09903_),
    .A2(_09904_),
    .B1(_09898_),
    .C1(_09900_),
    .Y(_09906_));
 sky130_fd_sc_hd__o221a_1 _37567_ (.A1(_07291_),
    .A2(_08574_),
    .B1(_09905_),
    .B2(_09906_),
    .C1(_08578_),
    .X(_09907_));
 sky130_fd_sc_hd__a211oi_1 _37568_ (.A1(_08575_),
    .A2(_08578_),
    .B1(_09905_),
    .C1(_09906_),
    .Y(_09908_));
 sky130_fd_sc_hd__nor2_1 _37569_ (.A(_09907_),
    .B(_09908_),
    .Y(_09909_));
 sky130_fd_sc_hd__xor2_1 _37570_ (.A(_08567_),
    .B(_09909_),
    .X(_09911_));
 sky130_fd_sc_hd__a21o_1 _37571_ (.A1(_08578_),
    .A2(_08579_),
    .B1(_08581_),
    .X(_09912_));
 sky130_fd_sc_hd__a31o_1 _37572_ (.A1(_09912_),
    .A2(_05780_),
    .A3(_03922_),
    .B1(_08583_),
    .X(_09913_));
 sky130_fd_sc_hd__and2_1 _37573_ (.A(_09911_),
    .B(_09913_),
    .X(_09914_));
 sky130_fd_sc_hd__inv_2 _37574_ (.A(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__a311o_1 _37575_ (.A1(_03922_),
    .A2(_05780_),
    .A3(_09912_),
    .B1(_08583_),
    .C1(_09911_),
    .X(_09916_));
 sky130_fd_sc_hd__nand2_1 _37576_ (.A(_09915_),
    .B(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__xor2_2 _37577_ (.A(_09896_),
    .B(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__o22ai_1 _37578_ (.A1(_08622_),
    .A2(_08626_),
    .B1(_08629_),
    .B2(_08630_),
    .Y(_09919_));
 sky130_fd_sc_hd__nand2_1 _37579_ (.A(_08619_),
    .B(_08625_),
    .Y(_09920_));
 sky130_fd_sc_hd__buf_1 _37580_ (.A(_08594_),
    .X(_09922_));
 sky130_fd_sc_hd__or3b_1 _37581_ (.A(_05823_),
    .B(_08611_),
    .C_N(_09922_),
    .X(_09923_));
 sky130_fd_sc_hd__buf_1 _37582_ (.A(_05805_),
    .X(_09924_));
 sky130_fd_sc_hd__clkbuf_2 _37583_ (.A(_07249_),
    .X(_09925_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37584_ (.A(_03957_),
    .X(_09926_));
 sky130_fd_sc_hd__a21oi_2 _37585_ (.A1(_09924_),
    .A2(_09925_),
    .B1(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__and3_1 _37586_ (.A(_09926_),
    .B(_05805_),
    .C(_07249_),
    .X(_09928_));
 sky130_fd_sc_hd__o211a_1 _37587_ (.A1(_09927_),
    .A2(_09928_),
    .B1(_08600_),
    .C1(_08603_),
    .X(_09929_));
 sky130_fd_sc_hd__buf_1 _37588_ (.A(_24745_),
    .X(_09930_));
 sky130_fd_sc_hd__o21a_1 _37589_ (.A1(_24735_),
    .A2(_24741_),
    .B1(_05813_),
    .X(_09931_));
 sky130_fd_sc_hd__a21oi_1 _37590_ (.A1(_24740_),
    .A2(_09930_),
    .B1(_09931_),
    .Y(_09933_));
 sky130_fd_sc_hd__a221oi_4 _37591_ (.A1(_09925_),
    .A2(_05809_),
    .B1(_08600_),
    .B2(_08603_),
    .C1(_09927_),
    .Y(_09934_));
 sky130_fd_sc_hd__nor3_2 _37592_ (.A(_09929_),
    .B(_09933_),
    .C(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__o21a_1 _37593_ (.A1(_09929_),
    .A2(_09934_),
    .B1(_09933_),
    .X(_09936_));
 sky130_fd_sc_hd__a211o_1 _37594_ (.A1(_08605_),
    .A2(_08612_),
    .B1(_09935_),
    .C1(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__o211ai_2 _37595_ (.A1(_09935_),
    .A2(_09936_),
    .B1(_08605_),
    .C1(_08612_),
    .Y(_09938_));
 sky130_fd_sc_hd__a22oi_1 _37596_ (.A1(_09922_),
    .A2(_09923_),
    .B1(_09937_),
    .B2(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__and4_1 _37597_ (.A(_09937_),
    .B(_09922_),
    .C(_09923_),
    .D(_09938_),
    .X(_09940_));
 sky130_fd_sc_hd__a211o_1 _37598_ (.A1(_08616_),
    .A2(_08618_),
    .B1(_09939_),
    .C1(_09940_),
    .X(_09941_));
 sky130_fd_sc_hd__o211ai_1 _37599_ (.A1(_09939_),
    .A2(_09940_),
    .B1(_08616_),
    .C1(_08618_),
    .Y(_09942_));
 sky130_fd_sc_hd__and3_1 _37600_ (.A(_08595_),
    .B(_09941_),
    .C(_09942_),
    .X(_09944_));
 sky130_fd_sc_hd__a21oi_1 _37601_ (.A1(_09941_),
    .A2(_09942_),
    .B1(_08595_),
    .Y(_09945_));
 sky130_fd_sc_hd__nor2_1 _37602_ (.A(_09944_),
    .B(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__xnor2_1 _37603_ (.A(_09920_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__nand2_1 _37604_ (.A(_09919_),
    .B(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__or2_1 _37605_ (.A(_09947_),
    .B(_09919_),
    .X(_09949_));
 sky130_fd_sc_hd__and2_1 _37606_ (.A(_09948_),
    .B(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__and2_1 _37607_ (.A(_09918_),
    .B(_09950_),
    .X(_09951_));
 sky130_fd_sc_hd__nor2_1 _37608_ (.A(_09918_),
    .B(_09950_),
    .Y(_09952_));
 sky130_fd_sc_hd__a21oi_1 _37609_ (.A1(_07211_),
    .A2(_05754_),
    .B1(_05756_),
    .Y(_09953_));
 sky130_fd_sc_hd__and3_1 _37610_ (.A(_07211_),
    .B(_05754_),
    .C(_05756_),
    .X(_09955_));
 sky130_fd_sc_hd__nor2_1 _37611_ (.A(_09953_),
    .B(_09955_),
    .Y(_09956_));
 sky130_fd_sc_hd__nor3_1 _37612_ (.A(_08533_),
    .B(_08545_),
    .C(_08546_),
    .Y(_09957_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37613_ (.A(net379),
    .X(_09958_));
 sky130_fd_sc_hd__nand2_1 _37614_ (.A(_03880_),
    .B(_05745_),
    .Y(_09959_));
 sky130_fd_sc_hd__o21a_1 _37615_ (.A1(_08535_),
    .A2(_05745_),
    .B1(_02489_),
    .X(_09960_));
 sky130_fd_sc_hd__and2_1 _37616_ (.A(\delay_line[16][12] ),
    .B(\delay_line[16][13] ),
    .X(_09961_));
 sky130_fd_sc_hd__nor2_1 _37617_ (.A(_08535_),
    .B(_05745_),
    .Y(_09962_));
 sky130_fd_sc_hd__o21a_1 _37618_ (.A1(_09961_),
    .A2(_09962_),
    .B1(_07210_),
    .X(_09963_));
 sky130_fd_sc_hd__a21o_1 _37619_ (.A1(_09959_),
    .A2(_09960_),
    .B1(_09963_),
    .X(_09964_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37620_ (.A(_09964_),
    .X(_09966_));
 sky130_fd_sc_hd__a21oi_2 _37621_ (.A1(_09958_),
    .A2(_08543_),
    .B1(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__and3_1 _37622_ (.A(_09966_),
    .B(net379),
    .C(_08543_),
    .X(_09968_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37623_ (.A(_02494_),
    .X(_09969_));
 sky130_fd_sc_hd__buf_1 _37624_ (.A(_03885_),
    .X(_09970_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37625_ (.A(_00834_),
    .X(_09971_));
 sky130_fd_sc_hd__a21o_1 _37626_ (.A1(_09969_),
    .A2(_09970_),
    .B1(_09971_),
    .X(_09972_));
 sky130_fd_sc_hd__o221ai_4 _37627_ (.A1(_08540_),
    .A2(_02498_),
    .B1(_09967_),
    .B2(_09968_),
    .C1(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__a211o_1 _37628_ (.A1(_08537_),
    .A2(_09972_),
    .B1(_09968_),
    .C1(_09967_),
    .X(_09974_));
 sky130_fd_sc_hd__o211a_1 _37629_ (.A1(_08546_),
    .A2(_09957_),
    .B1(_09973_),
    .C1(_09974_),
    .X(_09975_));
 sky130_fd_sc_hd__a211oi_1 _37630_ (.A1(_09973_),
    .A2(_09974_),
    .B1(_08546_),
    .C1(_09957_),
    .Y(_09977_));
 sky130_fd_sc_hd__nor2_1 _37631_ (.A(_09975_),
    .B(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__xnor2_1 _37632_ (.A(_09956_),
    .B(_09978_),
    .Y(_09979_));
 sky130_fd_sc_hd__o31a_1 _37633_ (.A1(_08530_),
    .A2(_08531_),
    .A3(_08552_),
    .B1(_08553_),
    .X(_09980_));
 sky130_fd_sc_hd__xor2_1 _37634_ (.A(_09979_),
    .B(_09980_),
    .X(_09981_));
 sky130_fd_sc_hd__xnor2_1 _37635_ (.A(_08530_),
    .B(_09981_),
    .Y(_09982_));
 sky130_fd_sc_hd__and3_1 _37636_ (.A(_08557_),
    .B(_08560_),
    .C(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__a21oi_1 _37637_ (.A1(_08557_),
    .A2(_08560_),
    .B1(_09982_),
    .Y(_09984_));
 sky130_fd_sc_hd__nor2_1 _37638_ (.A(_09983_),
    .B(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__and3_1 _37639_ (.A(_08527_),
    .B(_08560_),
    .C(_08561_),
    .X(_09986_));
 sky130_fd_sc_hd__a21oi_2 _37640_ (.A1(_08564_),
    .A2(_08563_),
    .B1(_09986_),
    .Y(_09988_));
 sky130_fd_sc_hd__xor2_2 _37641_ (.A(_09985_),
    .B(_09988_),
    .X(_09989_));
 sky130_fd_sc_hd__o21a_1 _37642_ (.A1(_09951_),
    .A2(_09952_),
    .B1(_09989_),
    .X(_09990_));
 sky130_fd_sc_hd__o32a_1 _37643_ (.A1(_08589_),
    .A2(_08631_),
    .A3(_08592_),
    .B1(_08565_),
    .B2(_08634_),
    .X(_09991_));
 sky130_fd_sc_hd__o31ai_1 _37644_ (.A1(_09951_),
    .A2(_09952_),
    .A3(_09989_),
    .B1(_09991_),
    .Y(_09992_));
 sky130_fd_sc_hd__nor3_2 _37645_ (.A(_09989_),
    .B(_09952_),
    .C(_09951_),
    .Y(_09993_));
 sky130_fd_sc_hd__o21bai_1 _37646_ (.A1(_09993_),
    .A2(_09990_),
    .B1_N(_09991_),
    .Y(_09994_));
 sky130_fd_sc_hd__o21a_2 _37647_ (.A1(_09990_),
    .A2(_09992_),
    .B1(_09994_),
    .X(_09995_));
 sky130_fd_sc_hd__xor2_4 _37648_ (.A(_09895_),
    .B(_09995_),
    .X(_09996_));
 sky130_fd_sc_hd__xnor2_4 _37649_ (.A(_09752_),
    .B(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__or2b_4 _37650_ (.A(_08686_),
    .B_N(_08763_),
    .X(_09999_));
 sky130_fd_sc_hd__o21bai_1 _37651_ (.A1(_08443_),
    .A2(_08446_),
    .B1_N(_08442_),
    .Y(_10000_));
 sky130_fd_sc_hd__a31o_1 _37652_ (.A1(_08399_),
    .A2(_08403_),
    .A3(_08438_),
    .B1(_08435_),
    .X(_10001_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37653_ (.A(_08406_),
    .X(_10002_));
 sky130_fd_sc_hd__and3_1 _37654_ (.A(_08410_),
    .B(_08408_),
    .C(_08401_),
    .X(_10003_));
 sky130_fd_sc_hd__clkbuf_2 _37655_ (.A(_07088_),
    .X(_10004_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37656_ (.A(_05871_),
    .X(_10005_));
 sky130_fd_sc_hd__o21a_1 _37657_ (.A1(_24504_),
    .A2(_24508_),
    .B1(_10005_),
    .X(_10006_));
 sky130_fd_sc_hd__a21oi_1 _37658_ (.A1(_08410_),
    .A2(_10004_),
    .B1(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__buf_1 _37659_ (.A(_07081_),
    .X(_10008_));
 sky130_fd_sc_hd__buf_1 _37660_ (.A(_05862_),
    .X(_10010_));
 sky130_fd_sc_hd__a21oi_1 _37661_ (.A1(_08411_),
    .A2(_10008_),
    .B1(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__and3_1 _37662_ (.A(_10010_),
    .B(_08411_),
    .C(_10008_),
    .X(_10012_));
 sky130_fd_sc_hd__a211oi_2 _37663_ (.A1(_08418_),
    .A2(_08416_),
    .B1(_10011_),
    .C1(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__o221a_1 _37664_ (.A1(_08411_),
    .A2(_07082_),
    .B1(_10011_),
    .B2(_10012_),
    .C1(_08416_),
    .X(_10014_));
 sky130_fd_sc_hd__nor3_1 _37665_ (.A(_10007_),
    .B(_10013_),
    .C(_10014_),
    .Y(_10015_));
 sky130_fd_sc_hd__o21a_1 _37666_ (.A1(_10014_),
    .A2(_10013_),
    .B1(_10007_),
    .X(_10016_));
 sky130_fd_sc_hd__nor2_1 _37667_ (.A(_10015_),
    .B(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__o21a_1 _37668_ (.A1(_08421_),
    .A2(net179),
    .B1(_10017_),
    .X(_10018_));
 sky130_fd_sc_hd__a311oi_4 _37669_ (.A1(_08416_),
    .A2(_08419_),
    .A3(_08420_),
    .B1(net179),
    .C1(_10017_),
    .Y(_10019_));
 sky130_fd_sc_hd__o22ai_2 _37670_ (.A1(_10003_),
    .A2(_10002_),
    .B1(_10018_),
    .B2(_10019_),
    .Y(_10021_));
 sky130_fd_sc_hd__or4_1 _37671_ (.A(_08406_),
    .B(_10003_),
    .C(_10019_),
    .D(_10018_),
    .X(_10022_));
 sky130_fd_sc_hd__o211a_1 _37672_ (.A1(_08428_),
    .A2(_08431_),
    .B1(_10021_),
    .C1(_10022_),
    .X(_10023_));
 sky130_fd_sc_hd__a211oi_2 _37673_ (.A1(_10021_),
    .A2(_10022_),
    .B1(_08428_),
    .C1(_08431_),
    .Y(_10024_));
 sky130_fd_sc_hd__a311o_1 _37674_ (.A1(_08399_),
    .A2(_08402_),
    .A3(_10002_),
    .B1(_10023_),
    .C1(_10024_),
    .X(_10025_));
 sky130_fd_sc_hd__o2111ai_1 _37675_ (.A1(_10023_),
    .A2(_10024_),
    .B1(_08399_),
    .C1(_08402_),
    .D1(_10002_),
    .Y(_10026_));
 sky130_fd_sc_hd__nand2_1 _37676_ (.A(_10025_),
    .B(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__xor2_1 _37677_ (.A(_10001_),
    .B(_10027_),
    .X(_10028_));
 sky130_fd_sc_hd__and2_1 _37678_ (.A(_10000_),
    .B(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__nor2_1 _37679_ (.A(_10028_),
    .B(_10000_),
    .Y(_10030_));
 sky130_fd_sc_hd__or2_2 _37680_ (.A(_10029_),
    .B(_10030_),
    .X(_10032_));
 sky130_fd_sc_hd__buf_1 _37681_ (.A(_07115_),
    .X(_10033_));
 sky130_fd_sc_hd__buf_1 _37682_ (.A(_08450_),
    .X(_10034_));
 sky130_fd_sc_hd__or3b_1 _37683_ (.A(_07132_),
    .B(_10034_),
    .C_N(_10033_),
    .X(_10035_));
 sky130_fd_sc_hd__buf_1 _37684_ (.A(_08453_),
    .X(_10036_));
 sky130_fd_sc_hd__buf_1 _37685_ (.A(net350),
    .X(_10037_));
 sky130_fd_sc_hd__buf_1 _37686_ (.A(_10037_),
    .X(_10038_));
 sky130_fd_sc_hd__buf_1 _37687_ (.A(_04179_),
    .X(_10039_));
 sky130_fd_sc_hd__nand2_1 _37688_ (.A(_10039_),
    .B(_10038_),
    .Y(_10040_));
 sky130_fd_sc_hd__or2_1 _37689_ (.A(_04179_),
    .B(_10037_),
    .X(_10041_));
 sky130_fd_sc_hd__a22o_1 _37690_ (.A1(_10036_),
    .A2(_10038_),
    .B1(_10040_),
    .B2(_10041_),
    .X(_10043_));
 sky130_fd_sc_hd__inv_2 _37691_ (.A(\delay_line[22][15] ),
    .Y(_10044_));
 sky130_fd_sc_hd__clkbuf_2 _37692_ (.A(_10044_),
    .X(_10045_));
 sky130_fd_sc_hd__or3b_1 _37693_ (.A(_10039_),
    .B(_10045_),
    .C_N(_10036_),
    .X(_10046_));
 sky130_fd_sc_hd__clkbuf_2 _37694_ (.A(_00520_),
    .X(_10047_));
 sky130_fd_sc_hd__and2b_1 _37695_ (.A_N(_07115_),
    .B(_08450_),
    .X(_10048_));
 sky130_fd_sc_hd__xor2_1 _37696_ (.A(_10047_),
    .B(_10048_),
    .X(_10049_));
 sky130_fd_sc_hd__a21oi_1 _37697_ (.A1(_10043_),
    .A2(_10046_),
    .B1(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__and3_1 _37698_ (.A(_10049_),
    .B(_10043_),
    .C(_10046_),
    .X(_10051_));
 sky130_fd_sc_hd__nand2_1 _37699_ (.A(_08457_),
    .B(_08460_),
    .Y(_10052_));
 sky130_fd_sc_hd__or3_1 _37700_ (.A(_10050_),
    .B(_10051_),
    .C(_10052_),
    .X(_10054_));
 sky130_fd_sc_hd__o21ai_2 _37701_ (.A1(_10050_),
    .A2(_10051_),
    .B1(_10052_),
    .Y(_10055_));
 sky130_fd_sc_hd__a22o_1 _37702_ (.A1(_10033_),
    .A2(_10035_),
    .B1(_10054_),
    .B2(_10055_),
    .X(_10056_));
 sky130_fd_sc_hd__buf_1 _37703_ (.A(_10034_),
    .X(_10057_));
 sky130_fd_sc_hd__o2111ai_2 _37704_ (.A1(_07132_),
    .A2(_10057_),
    .B1(_10033_),
    .C1(_10055_),
    .D1(_10054_),
    .Y(_10058_));
 sky130_fd_sc_hd__and2_1 _37705_ (.A(_10056_),
    .B(_10058_),
    .X(_10059_));
 sky130_fd_sc_hd__a311o_1 _37706_ (.A1(_08462_),
    .A2(_08460_),
    .A3(_08461_),
    .B1(net198),
    .C1(_10059_),
    .X(_10060_));
 sky130_fd_sc_hd__o21ai_1 _37707_ (.A1(_08464_),
    .A2(net198),
    .B1(_10059_),
    .Y(_10061_));
 sky130_fd_sc_hd__and3_1 _37708_ (.A(_10060_),
    .B(_10061_),
    .C(_08449_),
    .X(_10062_));
 sky130_fd_sc_hd__a21oi_1 _37709_ (.A1(_10060_),
    .A2(_10061_),
    .B1(_08449_),
    .Y(_10063_));
 sky130_fd_sc_hd__a21boi_1 _37710_ (.A1(_08468_),
    .A2(_07114_),
    .B1_N(_08469_),
    .Y(_10065_));
 sky130_fd_sc_hd__o21ai_1 _37711_ (.A1(_10062_),
    .A2(_10063_),
    .B1(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__or3_1 _37712_ (.A(_10065_),
    .B(_10062_),
    .C(_10063_),
    .X(_10067_));
 sky130_fd_sc_hd__a21o_1 _37713_ (.A1(_07144_),
    .A2(_07142_),
    .B1(_07139_),
    .X(_10068_));
 sky130_fd_sc_hd__a21o_1 _37714_ (.A1(_10068_),
    .A2(_08475_),
    .B1(_08473_),
    .X(_10069_));
 sky130_fd_sc_hd__a21oi_1 _37715_ (.A1(_10066_),
    .A2(_10067_),
    .B1(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__and3_1 _37716_ (.A(_10066_),
    .B(_10067_),
    .C(_10069_),
    .X(_10071_));
 sky130_fd_sc_hd__a31o_1 _37717_ (.A1(_08504_),
    .A2(_08505_),
    .A3(_08507_),
    .B1(_08509_),
    .X(_10072_));
 sky130_fd_sc_hd__nor2_1 _37718_ (.A(_05961_),
    .B(_08491_),
    .Y(_10073_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37719_ (.A(_02322_),
    .X(_10074_));
 sky130_fd_sc_hd__o211a_1 _37720_ (.A1(_07167_),
    .A2(_10074_),
    .B1(_05961_),
    .C1(_07166_),
    .X(_10076_));
 sky130_fd_sc_hd__and2_1 _37721_ (.A(net341),
    .B(\delay_line[24][13] ),
    .X(_10077_));
 sky130_fd_sc_hd__nor2_1 _37722_ (.A(net341),
    .B(_05947_),
    .Y(_10078_));
 sky130_fd_sc_hd__nor2_1 _37723_ (.A(_10077_),
    .B(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__o21a_1 _37724_ (.A1(net341),
    .A2(_05947_),
    .B1(\delay_line[24][11] ),
    .X(_10080_));
 sky130_fd_sc_hd__nand2_1 _37725_ (.A(_04213_),
    .B(_05947_),
    .Y(_10081_));
 sky130_fd_sc_hd__a2bb2o_1 _37726_ (.A1_N(_07153_),
    .A2_N(_10079_),
    .B1(_10080_),
    .B2(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__buf_1 _37727_ (.A(_10082_),
    .X(_10083_));
 sky130_fd_sc_hd__a21oi_2 _37728_ (.A1(_08488_),
    .A2(_08487_),
    .B1(_10083_),
    .Y(_10084_));
 sky130_fd_sc_hd__and3_1 _37729_ (.A(_10083_),
    .B(_08488_),
    .C(_08487_),
    .X(_10085_));
 sky130_fd_sc_hd__buf_1 _37730_ (.A(_04214_),
    .X(_10087_));
 sky130_fd_sc_hd__a21o_1 _37731_ (.A1(_10074_),
    .A2(_10087_),
    .B1(_00560_),
    .X(_10088_));
 sky130_fd_sc_hd__o221ai_4 _37732_ (.A1(_08483_),
    .A2(_08484_),
    .B1(_10084_),
    .B2(_10085_),
    .C1(_10088_),
    .Y(_10089_));
 sky130_fd_sc_hd__a211o_1 _37733_ (.A1(_08479_),
    .A2(_10088_),
    .B1(_10085_),
    .C1(_10084_),
    .X(_10090_));
 sky130_fd_sc_hd__nand2_1 _37734_ (.A(_08490_),
    .B(_08495_),
    .Y(_10091_));
 sky130_fd_sc_hd__and3_1 _37735_ (.A(_10089_),
    .B(_10090_),
    .C(_10091_),
    .X(_10092_));
 sky130_fd_sc_hd__a21oi_1 _37736_ (.A1(_10089_),
    .A2(_10090_),
    .B1(_10091_),
    .Y(_10093_));
 sky130_fd_sc_hd__nor4_1 _37737_ (.A(_10073_),
    .B(_10076_),
    .C(_10092_),
    .D(_10093_),
    .Y(_10094_));
 sky130_fd_sc_hd__o22a_1 _37738_ (.A1(_10073_),
    .A2(_10076_),
    .B1(_10092_),
    .B2(_10093_),
    .X(_10095_));
 sky130_fd_sc_hd__o211a_1 _37739_ (.A1(_10094_),
    .A2(_10095_),
    .B1(_08499_),
    .C1(_08504_),
    .X(_10096_));
 sky130_fd_sc_hd__a211o_1 _37740_ (.A1(_08499_),
    .A2(_08504_),
    .B1(_10094_),
    .C1(_10095_),
    .X(_10098_));
 sky130_fd_sc_hd__inv_2 _37741_ (.A(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__or3b_2 _37742_ (.A(_10096_),
    .B(_10099_),
    .C_N(_08500_),
    .X(_10100_));
 sky130_fd_sc_hd__nand2_1 _37743_ (.A(_10072_),
    .B(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__a2bb2o_1 _37744_ (.A1_N(_10096_),
    .A2_N(_10099_),
    .B1(_04225_),
    .B2(_07169_),
    .X(_10102_));
 sky130_fd_sc_hd__inv_2 _37745_ (.A(_10102_),
    .Y(_10103_));
 sky130_fd_sc_hd__a21o_1 _37746_ (.A1(_10102_),
    .A2(_10100_),
    .B1(_10072_),
    .X(_10104_));
 sky130_fd_sc_hd__o21ai_2 _37747_ (.A1(_10101_),
    .A2(_10103_),
    .B1(_10104_),
    .Y(_10105_));
 sky130_fd_sc_hd__a21oi_2 _37748_ (.A1(_08516_),
    .A2(_08515_),
    .B1(_08513_),
    .Y(_10106_));
 sky130_fd_sc_hd__or2_1 _37749_ (.A(_10105_),
    .B(_10106_),
    .X(_10107_));
 sky130_fd_sc_hd__nand2_1 _37750_ (.A(_10106_),
    .B(_10105_),
    .Y(_10109_));
 sky130_fd_sc_hd__or4bb_1 _37751_ (.A(_10070_),
    .B(_10071_),
    .C_N(_10107_),
    .D_N(_10109_),
    .X(_10110_));
 sky130_fd_sc_hd__a2bb2o_1 _37752_ (.A1_N(_10070_),
    .A2_N(_10071_),
    .B1(_10107_),
    .B2(_10109_),
    .X(_10111_));
 sky130_fd_sc_hd__nand2_1 _37753_ (.A(_10110_),
    .B(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__xnor2_1 _37754_ (.A(_10032_),
    .B(_10112_),
    .Y(_10113_));
 sky130_fd_sc_hd__a21oi_1 _37755_ (.A1(_08760_),
    .A2(_09999_),
    .B1(_10113_),
    .Y(_10114_));
 sky130_fd_sc_hd__and3_1 _37756_ (.A(_08760_),
    .B(_09999_),
    .C(_10113_),
    .X(_10115_));
 sky130_fd_sc_hd__nor2_2 _37757_ (.A(_10114_),
    .B(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__nand3b_1 _37758_ (.A_N(_08476_),
    .B(_08517_),
    .C(_08477_),
    .Y(_10117_));
 sky130_fd_sc_hd__a21bo_2 _37759_ (.A1(_08447_),
    .A2(_08518_),
    .B1_N(_10117_),
    .X(_10118_));
 sky130_fd_sc_hd__xnor2_4 _37760_ (.A(_10116_),
    .B(_10118_),
    .Y(_10120_));
 sky130_fd_sc_hd__or2b_1 _37761_ (.A(_09997_),
    .B_N(_10120_),
    .X(_10121_));
 sky130_fd_sc_hd__or2b_1 _37762_ (.A(_10120_),
    .B_N(_09997_),
    .X(_10122_));
 sky130_fd_sc_hd__o21a_1 _37763_ (.A1(_08524_),
    .A2(_08772_),
    .B1(_08771_),
    .X(_10123_));
 sky130_fd_sc_hd__a21oi_1 _37764_ (.A1(_10121_),
    .A2(_10122_),
    .B1(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__o2111ai_1 _37765_ (.A1(_08524_),
    .A2(_08772_),
    .B1(_10121_),
    .C1(_10122_),
    .D1(_08771_),
    .Y(_10125_));
 sky130_fd_sc_hd__or2b_1 _37766_ (.A(_10124_),
    .B_N(_10125_),
    .X(_10126_));
 sky130_fd_sc_hd__o21bai_4 _37767_ (.A1(_08856_),
    .A2(_08928_),
    .B1_N(_08854_),
    .Y(_10127_));
 sky130_fd_sc_hd__o21ai_2 _37768_ (.A1(_08849_),
    .A2(_08798_),
    .B1(_08850_),
    .Y(_10128_));
 sky130_fd_sc_hd__a21o_1 _37769_ (.A1(_08846_),
    .A2(_08845_),
    .B1(_08842_),
    .X(_10129_));
 sky130_fd_sc_hd__o21a_1 _37770_ (.A1(_05508_),
    .A2(_05501_),
    .B1(net329),
    .X(_10131_));
 sky130_fd_sc_hd__and3_1 _37771_ (.A(_02214_),
    .B(_00969_),
    .C(_10131_),
    .X(_10132_));
 sky130_fd_sc_hd__a21oi_1 _37772_ (.A1(_02214_),
    .A2(_00969_),
    .B1(_10131_),
    .Y(_10133_));
 sky130_fd_sc_hd__a211oi_1 _37773_ (.A1(_08827_),
    .A2(_08829_),
    .B1(_10132_),
    .C1(_10133_),
    .Y(_10134_));
 sky130_fd_sc_hd__o221a_1 _37774_ (.A1(_05496_),
    .A2(_07036_),
    .B1(_10132_),
    .B2(_10133_),
    .C1(_08829_),
    .X(_10135_));
 sky130_fd_sc_hd__nor2_1 _37775_ (.A(_10134_),
    .B(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__xor2_1 _37776_ (.A(_24362_),
    .B(_10136_),
    .X(_10137_));
 sky130_fd_sc_hd__o21ba_1 _37777_ (.A1(_08835_),
    .A2(_08836_),
    .B1_N(_10137_),
    .X(_10138_));
 sky130_fd_sc_hd__o211a_1 _37778_ (.A1(_23162_),
    .A2(_08832_),
    .B1(_08834_),
    .C1(_10137_),
    .X(_10139_));
 sky130_fd_sc_hd__or2_1 _37779_ (.A(_10138_),
    .B(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__xnor2_1 _37780_ (.A(_08839_),
    .B(_10140_),
    .Y(_10142_));
 sky130_fd_sc_hd__xor2_1 _37781_ (.A(_10129_),
    .B(_10142_),
    .X(_10143_));
 sky130_fd_sc_hd__a2111o_1 _37782_ (.A1(_04292_),
    .A2(_04299_),
    .B1(_05537_),
    .C1(_08814_),
    .D1(_07023_),
    .X(_10144_));
 sky130_fd_sc_hd__o32a_1 _37783_ (.A1(_08810_),
    .A2(_08812_),
    .A3(_10144_),
    .B1(_08803_),
    .B2(_08816_),
    .X(_10145_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37784_ (.A(_02207_),
    .X(_10146_));
 sky130_fd_sc_hd__nand2_1 _37785_ (.A(_00995_),
    .B(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__nor2_1 _37786_ (.A(_02207_),
    .B(net336),
    .Y(_10148_));
 sky130_fd_sc_hd__and2_1 _37787_ (.A(_02207_),
    .B(net336),
    .X(_10149_));
 sky130_fd_sc_hd__nor3_1 _37788_ (.A(_23141_),
    .B(_10148_),
    .C(_10149_),
    .Y(_10150_));
 sky130_fd_sc_hd__o21a_1 _37789_ (.A1(_10148_),
    .A2(_10149_),
    .B1(_23141_),
    .X(_10151_));
 sky130_fd_sc_hd__or2_1 _37790_ (.A(_10150_),
    .B(_10151_),
    .X(_10153_));
 sky130_fd_sc_hd__a21oi_2 _37791_ (.A1(_10147_),
    .A2(_08807_),
    .B1(_10153_),
    .Y(_10154_));
 sky130_fd_sc_hd__and3_1 _37792_ (.A(_10147_),
    .B(_08807_),
    .C(_10153_),
    .X(_10155_));
 sky130_fd_sc_hd__nor2_1 _37793_ (.A(_10154_),
    .B(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__a21oi_1 _37794_ (.A1(_08814_),
    .A2(_08813_),
    .B1(_08810_),
    .Y(_10157_));
 sky130_fd_sc_hd__xnor2_1 _37795_ (.A(_10156_),
    .B(_10157_),
    .Y(_10158_));
 sky130_fd_sc_hd__xor2_1 _37796_ (.A(_08802_),
    .B(_10158_),
    .X(_10159_));
 sky130_fd_sc_hd__or2b_1 _37797_ (.A(_10145_),
    .B_N(_10159_),
    .X(_10160_));
 sky130_fd_sc_hd__or2b_1 _37798_ (.A(_10159_),
    .B_N(_10145_),
    .X(_10161_));
 sky130_fd_sc_hd__o211ai_2 _37799_ (.A1(_08821_),
    .A2(_08825_),
    .B1(_10160_),
    .C1(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__a211o_1 _37800_ (.A1(_10160_),
    .A2(_10161_),
    .B1(_08821_),
    .C1(_08825_),
    .X(_10164_));
 sky130_fd_sc_hd__nand3_1 _37801_ (.A(_10143_),
    .B(_10162_),
    .C(_10164_),
    .Y(_10165_));
 sky130_fd_sc_hd__a21o_1 _37802_ (.A1(_10164_),
    .A2(_10162_),
    .B1(_10143_),
    .X(_10166_));
 sky130_fd_sc_hd__o21a_1 _37803_ (.A1(_08782_),
    .A2(_08794_),
    .B1(_08797_),
    .X(_10167_));
 sky130_fd_sc_hd__buf_1 _37804_ (.A(_06995_),
    .X(_10168_));
 sky130_fd_sc_hd__nand2_1 _37805_ (.A(_04266_),
    .B(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__nand2_1 _37806_ (.A(_05559_),
    .B(_06992_),
    .Y(_10170_));
 sky130_fd_sc_hd__and2_1 _37807_ (.A(_10169_),
    .B(_10170_),
    .X(_10171_));
 sky130_fd_sc_hd__o221ai_4 _37808_ (.A1(_10169_),
    .A2(_08784_),
    .B1(_04266_),
    .B2(_06993_),
    .C1(_04267_),
    .Y(_10172_));
 sky130_fd_sc_hd__o21ai_1 _37809_ (.A1(_04267_),
    .A2(_10171_),
    .B1(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__nor2_1 _37810_ (.A(_08788_),
    .B(_08790_),
    .Y(_10175_));
 sky130_fd_sc_hd__xor2_1 _37811_ (.A(_10173_),
    .B(_10175_),
    .X(_10176_));
 sky130_fd_sc_hd__xor2_2 _37812_ (.A(_08793_),
    .B(_10176_),
    .X(_10177_));
 sky130_fd_sc_hd__xnor2_2 _37813_ (.A(_10167_),
    .B(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__a21oi_1 _37814_ (.A1(_10165_),
    .A2(_10166_),
    .B1(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__and3_1 _37815_ (.A(_10178_),
    .B(_10165_),
    .C(_10166_),
    .X(_10180_));
 sky130_fd_sc_hd__or2_2 _37816_ (.A(_10179_),
    .B(_10180_),
    .X(_10181_));
 sky130_fd_sc_hd__xnor2_1 _37817_ (.A(_10128_),
    .B(_10181_),
    .Y(_10182_));
 sky130_fd_sc_hd__nor2b_2 _37818_ (.A(_04409_),
    .B_N(\delay_line[29][15] ),
    .Y(_10183_));
 sky130_fd_sc_hd__and2b_1 _37819_ (.A_N(\delay_line[29][15] ),
    .B(_04409_),
    .X(_10184_));
 sky130_fd_sc_hd__nor2_2 _37820_ (.A(_10183_),
    .B(_10184_),
    .Y(_10186_));
 sky130_fd_sc_hd__o21ba_1 _37821_ (.A1(_06943_),
    .A2(_08887_),
    .B1_N(_08886_),
    .X(_10187_));
 sky130_fd_sc_hd__xor2_2 _37822_ (.A(_10186_),
    .B(_10187_),
    .X(_10188_));
 sky130_fd_sc_hd__nand2_1 _37823_ (.A(_05445_),
    .B(_06945_),
    .Y(_10189_));
 sky130_fd_sc_hd__o2bb2a_1 _37824_ (.A1_N(_08891_),
    .A2_N(_08892_),
    .B1(_10189_),
    .B2(_08889_),
    .X(_10190_));
 sky130_fd_sc_hd__nand2_1 _37825_ (.A(_10188_),
    .B(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__or2_1 _37826_ (.A(_10188_),
    .B(_10190_),
    .X(_10192_));
 sky130_fd_sc_hd__nand2_1 _37827_ (.A(_10191_),
    .B(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__o211a_1 _37828_ (.A1(_08908_),
    .A2(_08909_),
    .B1(_06919_),
    .C1(_08894_),
    .X(_10194_));
 sky130_fd_sc_hd__o21a_1 _37829_ (.A1(_08913_),
    .A2(_10194_),
    .B1(_08911_),
    .X(_10195_));
 sky130_fd_sc_hd__or4b_1 _37830_ (.A(_02089_),
    .B(_08903_),
    .C(_08906_),
    .D_N(_05477_),
    .X(_10197_));
 sky130_fd_sc_hd__o21a_1 _37831_ (.A1(_08895_),
    .A2(_08896_),
    .B1(_05455_),
    .X(_10198_));
 sky130_fd_sc_hd__buf_1 _37832_ (.A(_05457_),
    .X(_10199_));
 sky130_fd_sc_hd__and3_1 _37833_ (.A(_05476_),
    .B(_02110_),
    .C(_10199_),
    .X(_10200_));
 sky130_fd_sc_hd__or4b_1 _37834_ (.A(_04399_),
    .B(_10198_),
    .C(_10200_),
    .D_N(_06925_),
    .X(_10201_));
 sky130_fd_sc_hd__a2bb2o_1 _37835_ (.A1_N(_10198_),
    .A2_N(_10200_),
    .B1(_23246_),
    .B2(_06925_),
    .X(_10202_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37836_ (.A(_08897_),
    .X(_10203_));
 sky130_fd_sc_hd__buf_1 _37837_ (.A(_05459_),
    .X(_10204_));
 sky130_fd_sc_hd__nor2_1 _37838_ (.A(_08902_),
    .B(_10204_),
    .Y(_10205_));
 sky130_fd_sc_hd__inv_2 _37839_ (.A(_05459_),
    .Y(_10206_));
 sky130_fd_sc_hd__nor2_1 _37840_ (.A(_02101_),
    .B(_10206_),
    .Y(_10208_));
 sky130_fd_sc_hd__nor2_1 _37841_ (.A(_10205_),
    .B(_10208_),
    .Y(_10209_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37842_ (.A(_10209_),
    .X(_10210_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37843_ (.A(net319),
    .X(_10211_));
 sky130_fd_sc_hd__o211ai_2 _37844_ (.A1(_10203_),
    .A2(_08898_),
    .B1(_10210_),
    .C1(_10211_),
    .Y(_10212_));
 sky130_fd_sc_hd__or2_1 _37845_ (.A(_10203_),
    .B(_08898_),
    .X(_10213_));
 sky130_fd_sc_hd__a2bb2o_1 _37846_ (.A1_N(_10205_),
    .A2_N(_10208_),
    .B1(_10211_),
    .B2(_10213_),
    .X(_10214_));
 sky130_fd_sc_hd__and4_1 _37847_ (.A(_10201_),
    .B(_10202_),
    .C(_10212_),
    .D(_10214_),
    .X(_10215_));
 sky130_fd_sc_hd__a22oi_2 _37848_ (.A1(_10201_),
    .A2(_10202_),
    .B1(_10212_),
    .B2(_10214_),
    .Y(_10216_));
 sky130_fd_sc_hd__buf_1 _37849_ (.A(\delay_line[30][15] ),
    .X(_10217_));
 sky130_fd_sc_hd__a31o_1 _37850_ (.A1(_10217_),
    .A2(_06908_),
    .A3(_10213_),
    .B1(_08908_),
    .X(_10219_));
 sky130_fd_sc_hd__nor3b_2 _37851_ (.A(_10215_),
    .B(_10216_),
    .C_N(_10219_),
    .Y(_10220_));
 sky130_fd_sc_hd__o21ba_1 _37852_ (.A1(_10215_),
    .A2(_10216_),
    .B1_N(_10219_),
    .X(_10221_));
 sky130_fd_sc_hd__a211oi_1 _37853_ (.A1(_08904_),
    .A2(_10197_),
    .B1(_10220_),
    .C1(_10221_),
    .Y(_10222_));
 sky130_fd_sc_hd__buf_1 _37854_ (.A(_10222_),
    .X(_10223_));
 sky130_fd_sc_hd__o211a_1 _37855_ (.A1(_10220_),
    .A2(_10221_),
    .B1(_08904_),
    .C1(_10197_),
    .X(_10224_));
 sky130_fd_sc_hd__nor3_2 _37856_ (.A(_10195_),
    .B(_10223_),
    .C(_10224_),
    .Y(_10225_));
 sky130_fd_sc_hd__o221a_1 _37857_ (.A1(_08913_),
    .A2(_10194_),
    .B1(_10222_),
    .B2(_10224_),
    .C1(_08911_),
    .X(_10226_));
 sky130_fd_sc_hd__or3_1 _37858_ (.A(_10225_),
    .B(_10226_),
    .C(_08918_),
    .X(_10227_));
 sky130_fd_sc_hd__o21ai_1 _37859_ (.A1(_10225_),
    .A2(_10226_),
    .B1(_08918_),
    .Y(_10228_));
 sky130_fd_sc_hd__nand2_1 _37860_ (.A(_10227_),
    .B(_10228_),
    .Y(_10230_));
 sky130_fd_sc_hd__a21oi_2 _37861_ (.A1(_08925_),
    .A2(_08923_),
    .B1(_08920_),
    .Y(_10231_));
 sky130_fd_sc_hd__xnor2_2 _37862_ (.A(_10230_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__xor2_2 _37863_ (.A(_10193_),
    .B(_10232_),
    .X(_10233_));
 sky130_fd_sc_hd__a21bo_1 _37864_ (.A1(_06960_),
    .A2(_08873_),
    .B1_N(_08874_),
    .X(_10234_));
 sky130_fd_sc_hd__o21ai_1 _37865_ (.A1(_08857_),
    .A2(_08858_),
    .B1(_05409_),
    .Y(_10235_));
 sky130_fd_sc_hd__nor2_1 _37866_ (.A(_23213_),
    .B(_04353_),
    .Y(_10236_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _37867_ (.A(_00885_),
    .X(_10237_));
 sky130_fd_sc_hd__nor2_1 _37868_ (.A(_10237_),
    .B(_06957_),
    .Y(_10238_));
 sky130_fd_sc_hd__nor3_1 _37869_ (.A(_08865_),
    .B(_10236_),
    .C(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__a2bb2o_1 _37870_ (.A1_N(_10236_),
    .A2_N(_10238_),
    .B1(_05423_),
    .B2(_08864_),
    .X(_10241_));
 sky130_fd_sc_hd__or2b_1 _37871_ (.A(_10239_),
    .B_N(_10241_),
    .X(_10242_));
 sky130_fd_sc_hd__xor2_1 _37872_ (.A(_10235_),
    .B(_10242_),
    .X(_10243_));
 sky130_fd_sc_hd__buf_1 _37873_ (.A(_04351_),
    .X(_10244_));
 sky130_fd_sc_hd__buf_1 _37874_ (.A(_05409_),
    .X(_10245_));
 sky130_fd_sc_hd__nor2_1 _37875_ (.A(_08857_),
    .B(_08858_),
    .Y(_10246_));
 sky130_fd_sc_hd__a31o_1 _37876_ (.A1(_10244_),
    .A2(_10245_),
    .A3(_10246_),
    .B1(_08870_),
    .X(_10247_));
 sky130_fd_sc_hd__nor2_1 _37877_ (.A(_10243_),
    .B(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__and2_1 _37878_ (.A(_10247_),
    .B(_10243_),
    .X(_10249_));
 sky130_fd_sc_hd__nor2_1 _37879_ (.A(_10248_),
    .B(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__and4_1 _37880_ (.A(_08865_),
    .B(_10250_),
    .C(_08862_),
    .D(_08863_),
    .X(_10252_));
 sky130_fd_sc_hd__nor2_1 _37881_ (.A(_08867_),
    .B(_10250_),
    .Y(_10253_));
 sky130_fd_sc_hd__nor2_1 _37882_ (.A(_10252_),
    .B(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__nor2_1 _37883_ (.A(_10234_),
    .B(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__and2_1 _37884_ (.A(_10254_),
    .B(_10234_),
    .X(_10256_));
 sky130_fd_sc_hd__nor2_1 _37885_ (.A(_08883_),
    .B(_08884_),
    .Y(_10257_));
 sky130_fd_sc_hd__nor2_1 _37886_ (.A(_08881_),
    .B(_10257_),
    .Y(_10258_));
 sky130_fd_sc_hd__o21ai_1 _37887_ (.A1(_10255_),
    .A2(_10256_),
    .B1(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__or2_1 _37888_ (.A(_10255_),
    .B(_10256_),
    .X(_10260_));
 sky130_fd_sc_hd__o21bai_1 _37889_ (.A1(_08881_),
    .A2(_10257_),
    .B1_N(_10260_),
    .Y(_10261_));
 sky130_fd_sc_hd__and2_1 _37890_ (.A(_10259_),
    .B(_10261_),
    .X(_10263_));
 sky130_fd_sc_hd__xor2_2 _37891_ (.A(_08878_),
    .B(_10263_),
    .X(_10264_));
 sky130_fd_sc_hd__xnor2_2 _37892_ (.A(_10233_),
    .B(_10264_),
    .Y(_10265_));
 sky130_fd_sc_hd__and2_1 _37893_ (.A(_10182_),
    .B(_10265_),
    .X(_10266_));
 sky130_fd_sc_hd__or2_1 _37894_ (.A(_10182_),
    .B(_10265_),
    .X(_10267_));
 sky130_fd_sc_hd__inv_2 _37895_ (.A(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__o221a_1 _37896_ (.A1(_08397_),
    .A2(_08519_),
    .B1(_10266_),
    .B2(_10268_),
    .C1(_08521_),
    .X(_10269_));
 sky130_fd_sc_hd__o21a_1 _37897_ (.A1(_08397_),
    .A2(_08519_),
    .B1(_08521_),
    .X(_10270_));
 sky130_fd_sc_hd__or3_1 _37898_ (.A(_10270_),
    .B(_10266_),
    .C(_10268_),
    .X(_10271_));
 sky130_fd_sc_hd__and2b_1 _37899_ (.A_N(_10269_),
    .B(_10271_),
    .X(_10272_));
 sky130_fd_sc_hd__xor2_2 _37900_ (.A(_10127_),
    .B(_10272_),
    .X(_10274_));
 sky130_fd_sc_hd__xor2_1 _37901_ (.A(_10126_),
    .B(_10274_),
    .X(_10275_));
 sky130_fd_sc_hd__o21a_1 _37902_ (.A1(_08937_),
    .A2(_08774_),
    .B1(_08775_),
    .X(_10276_));
 sky130_fd_sc_hd__xor2_1 _37903_ (.A(_10275_),
    .B(_10276_),
    .X(_10277_));
 sky130_fd_sc_hd__o21ba_1 _37904_ (.A1(_09750_),
    .A2(_09751_),
    .B1_N(_10277_),
    .X(_10278_));
 sky130_fd_sc_hd__nor3b_1 _37905_ (.A(_09750_),
    .B(_09751_),
    .C_N(_10277_),
    .Y(_10279_));
 sky130_fd_sc_hd__or2_2 _37906_ (.A(_10278_),
    .B(_10279_),
    .X(_10280_));
 sky130_fd_sc_hd__xor2_1 _37907_ (.A(_09572_),
    .B(_10280_),
    .X(_10281_));
 sky130_fd_sc_hd__nand3_1 _37908_ (.A(_09562_),
    .B(_09566_),
    .C(_09567_),
    .Y(_10282_));
 sky130_fd_sc_hd__nand2_2 _37909_ (.A(_10281_),
    .B(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__a21oi_2 _37910_ (.A1(_09571_),
    .A2(_08941_),
    .B1(_10280_),
    .Y(_10285_));
 sky130_fd_sc_hd__and3_1 _37911_ (.A(_09571_),
    .B(_08941_),
    .C(_10280_),
    .X(_10286_));
 sky130_fd_sc_hd__inv_2 _37912_ (.A(_08176_),
    .Y(_10287_));
 sky130_fd_sc_hd__o211a_1 _37913_ (.A1(_08177_),
    .A2(_10287_),
    .B1(_09562_),
    .C1(_09566_),
    .X(_10288_));
 sky130_fd_sc_hd__o22ai_4 _37914_ (.A1(_10285_),
    .A2(_10286_),
    .B1(_09568_),
    .B2(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__o22ai_4 _37915_ (.A1(_08190_),
    .A2(_08942_),
    .B1(_08188_),
    .B2(_08945_),
    .Y(_10290_));
 sky130_fd_sc_hd__o211ai_4 _37916_ (.A1(_09570_),
    .A2(_10283_),
    .B1(_10289_),
    .C1(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__o21ai_1 _37917_ (.A1(_09570_),
    .A2(_10283_),
    .B1(_10289_),
    .Y(_10292_));
 sky130_fd_sc_hd__o22a_1 _37918_ (.A1(_08190_),
    .A2(_08942_),
    .B1(_08188_),
    .B2(_08945_),
    .X(_10293_));
 sky130_fd_sc_hd__nand2_1 _37919_ (.A(_10292_),
    .B(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__buf_1 _37920_ (.A(_08959_),
    .X(_10296_));
 sky130_fd_sc_hd__buf_1 _37921_ (.A(_10296_),
    .X(_10297_));
 sky130_fd_sc_hd__o2bb2a_1 _37922_ (.A1_N(_08957_),
    .A2_N(_10297_),
    .B1(_03011_),
    .B2(_23691_),
    .X(_10298_));
 sky130_fd_sc_hd__and3_1 _37923_ (.A(_08957_),
    .B(_10297_),
    .C(_08971_),
    .X(_10299_));
 sky130_fd_sc_hd__nor2_1 _37924_ (.A(_04558_),
    .B(_25224_),
    .Y(_10300_));
 sky130_fd_sc_hd__and2_1 _37925_ (.A(_25224_),
    .B(_04558_),
    .X(_10301_));
 sky130_fd_sc_hd__clkbuf_2 _37926_ (.A(_04559_),
    .X(_10302_));
 sky130_fd_sc_hd__and3_1 _37927_ (.A(_04533_),
    .B(_07537_),
    .C(_09002_),
    .X(_10303_));
 sky130_fd_sc_hd__buf_4 _37928_ (.A(_07537_),
    .X(_10304_));
 sky130_fd_sc_hd__a21oi_4 _37929_ (.A1(_10304_),
    .A2(_09002_),
    .B1(_04533_),
    .Y(_10305_));
 sky130_fd_sc_hd__or3_2 _37930_ (.A(_10302_),
    .B(_10303_),
    .C(_10305_),
    .X(_10307_));
 sky130_fd_sc_hd__o21ai_2 _37931_ (.A1(_10303_),
    .A2(_10305_),
    .B1(_10302_),
    .Y(_10308_));
 sky130_fd_sc_hd__nor3_1 _37932_ (.A(_08982_),
    .B(_08977_),
    .C(_08980_),
    .Y(_10309_));
 sky130_fd_sc_hd__a211o_1 _37933_ (.A1(_10307_),
    .A2(_10308_),
    .B1(_08977_),
    .C1(_10309_),
    .X(_10310_));
 sky130_fd_sc_hd__o211ai_4 _37934_ (.A1(_08977_),
    .A2(net196),
    .B1(_10307_),
    .C1(_10308_),
    .Y(_10311_));
 sky130_fd_sc_hd__or4bb_4 _37935_ (.A(_10300_),
    .B(_10301_),
    .C_N(_10310_),
    .D_N(_10311_),
    .X(_10312_));
 sky130_fd_sc_hd__a2bb2o_1 _37936_ (.A1_N(_10300_),
    .A2_N(_10301_),
    .B1(_10310_),
    .B2(_10311_),
    .X(_10313_));
 sky130_fd_sc_hd__a211oi_1 _37937_ (.A1(_10312_),
    .A2(_10313_),
    .B1(_08986_),
    .C1(net166),
    .Y(_10314_));
 sky130_fd_sc_hd__o211a_1 _37938_ (.A1(_08986_),
    .A2(net166),
    .B1(_10312_),
    .C1(_10313_),
    .X(_10315_));
 sky130_fd_sc_hd__o22a_1 _37939_ (.A1(_10298_),
    .A2(_10299_),
    .B1(_10314_),
    .B2(_10315_),
    .X(_10316_));
 sky130_fd_sc_hd__nor4_1 _37940_ (.A(_10298_),
    .B(_10299_),
    .C(_10314_),
    .D(_10315_),
    .Y(_10318_));
 sky130_fd_sc_hd__a211oi_1 _37941_ (.A1(_06643_),
    .A2(_08997_),
    .B1(_09013_),
    .C1(_09014_),
    .Y(_10319_));
 sky130_fd_sc_hd__nor4_2 _37942_ (.A(_06636_),
    .B(_09000_),
    .C(_04528_),
    .D(_08158_),
    .Y(_10320_));
 sky130_fd_sc_hd__buf_1 _37943_ (.A(_04528_),
    .X(_10321_));
 sky130_fd_sc_hd__o22a_1 _37944_ (.A1(_08158_),
    .A2(_06636_),
    .B1(_09000_),
    .B2(_10321_),
    .X(_10322_));
 sky130_fd_sc_hd__or4b_2 _37945_ (.A(_07541_),
    .B(_10320_),
    .C(_10322_),
    .D_N(_09007_),
    .X(_10323_));
 sky130_fd_sc_hd__clkbuf_4 _37946_ (.A(_07541_),
    .X(_10324_));
 sky130_fd_sc_hd__o32ai_4 _37947_ (.A1(_09004_),
    .A2(_10324_),
    .A3(_09001_),
    .B1(_10320_),
    .B2(_10322_),
    .Y(_10325_));
 sky130_fd_sc_hd__a221o_1 _37948_ (.A1(_08159_),
    .A2(_08166_),
    .B1(_10323_),
    .B2(_10325_),
    .C1(_08164_),
    .X(_10326_));
 sky130_fd_sc_hd__o211ai_1 _37949_ (.A1(_08164_),
    .A2(_08167_),
    .B1(_10323_),
    .C1(_10325_),
    .Y(_10327_));
 sky130_fd_sc_hd__nor4_1 _37950_ (.A(_06633_),
    .B(_09005_),
    .C(_06635_),
    .D(_09008_),
    .Y(_10329_));
 sky130_fd_sc_hd__or2_1 _37951_ (.A(_10329_),
    .B(_09014_),
    .X(_10330_));
 sky130_fd_sc_hd__and3_1 _37952_ (.A(_10326_),
    .B(_10327_),
    .C(_10330_),
    .X(_10331_));
 sky130_fd_sc_hd__a21oi_1 _37953_ (.A1(_10326_),
    .A2(_10327_),
    .B1(_10330_),
    .Y(_10332_));
 sky130_fd_sc_hd__nor2_1 _37954_ (.A(_10331_),
    .B(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__nor3_1 _37955_ (.A(_10319_),
    .B(_09017_),
    .C(_10333_),
    .Y(_10334_));
 sky130_fd_sc_hd__o21a_1 _37956_ (.A1(_10319_),
    .A2(_09017_),
    .B1(_10333_),
    .X(_10335_));
 sky130_fd_sc_hd__nor2_1 _37957_ (.A(_10334_),
    .B(_10335_),
    .Y(_10336_));
 sky130_fd_sc_hd__or3b_1 _37958_ (.A(_10316_),
    .B(net146),
    .C_N(_10336_),
    .X(_10337_));
 sky130_fd_sc_hd__nor2_1 _37959_ (.A(_10316_),
    .B(net146),
    .Y(_10338_));
 sky130_fd_sc_hd__or2_1 _37960_ (.A(_10336_),
    .B(_10338_),
    .X(_10340_));
 sky130_fd_sc_hd__nand2_1 _37961_ (.A(_10337_),
    .B(_10340_),
    .Y(_10341_));
 sky130_fd_sc_hd__nand2_1 _37962_ (.A(_08181_),
    .B(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__a21oi_2 _37963_ (.A1(_08186_),
    .A2(_08175_),
    .B1(_10342_),
    .Y(_10343_));
 sky130_fd_sc_hd__nand2_1 _37964_ (.A(_08186_),
    .B(_08175_),
    .Y(_10344_));
 sky130_fd_sc_hd__a21oi_1 _37965_ (.A1(_08181_),
    .A2(_10344_),
    .B1(_10341_),
    .Y(_10345_));
 sky130_fd_sc_hd__a21o_1 _37966_ (.A1(_08995_),
    .A2(_09019_),
    .B1(_09024_),
    .X(_10346_));
 sky130_fd_sc_hd__inv_2 _37967_ (.A(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__o21ai_1 _37968_ (.A1(_10343_),
    .A2(_10345_),
    .B1(_10347_),
    .Y(_10348_));
 sky130_fd_sc_hd__o21ai_2 _37969_ (.A1(_06651_),
    .A2(_06653_),
    .B1(_06655_),
    .Y(_10349_));
 sky130_fd_sc_hd__a32oi_4 _37970_ (.A1(_08170_),
    .A2(_08171_),
    .A3(_08172_),
    .B1(_10349_),
    .B2(_06654_),
    .Y(_10351_));
 sky130_fd_sc_hd__o211a_1 _37971_ (.A1(_08176_),
    .A2(_08177_),
    .B1(_08178_),
    .C1(_08179_),
    .X(_10352_));
 sky130_fd_sc_hd__o21bai_4 _37972_ (.A1(_10352_),
    .A2(_10351_),
    .B1_N(_10341_),
    .Y(_10353_));
 sky130_fd_sc_hd__o211ai_1 _37973_ (.A1(_10342_),
    .A2(_10351_),
    .B1(_10346_),
    .C1(_10353_),
    .Y(_10354_));
 sky130_fd_sc_hd__nand2_1 _37974_ (.A(_10348_),
    .B(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__a21o_1 _37975_ (.A1(_10291_),
    .A2(_10294_),
    .B1(_10355_),
    .X(_10356_));
 sky130_fd_sc_hd__nand3_2 _37976_ (.A(_10355_),
    .B(_10291_),
    .C(_10294_),
    .Y(_10357_));
 sky130_fd_sc_hd__a22o_1 _37977_ (.A1(_08950_),
    .A2(_09114_),
    .B1(_10356_),
    .B2(_10357_),
    .X(_10358_));
 sky130_fd_sc_hd__o2111ai_4 _37978_ (.A1(_09039_),
    .A2(_09040_),
    .B1(_10356_),
    .C1(_10357_),
    .D1(_08950_),
    .Y(_10359_));
 sky130_fd_sc_hd__inv_2 _37979_ (.A(_09077_),
    .Y(_10360_));
 sky130_fd_sc_hd__o21ai_2 _37980_ (.A1(_07563_),
    .A2(_07571_),
    .B1(_09027_),
    .Y(_10362_));
 sky130_fd_sc_hd__or2_1 _37981_ (.A(_09069_),
    .B(_09070_),
    .X(_10363_));
 sky130_fd_sc_hd__a211o_1 _37982_ (.A1(_08958_),
    .A2(_08962_),
    .B1(_07510_),
    .C1(_08960_),
    .X(_10364_));
 sky130_fd_sc_hd__and3_1 _37983_ (.A(_10364_),
    .B(_08957_),
    .C(_07502_),
    .X(_10365_));
 sky130_fd_sc_hd__a21o_1 _37984_ (.A1(_20957_),
    .A2(_20958_),
    .B1(_04573_),
    .X(_10366_));
 sky130_fd_sc_hd__nand2_1 _37985_ (.A(_04575_),
    .B(_20959_),
    .Y(_10367_));
 sky130_fd_sc_hd__a21o_1 _37986_ (.A1(_04572_),
    .A2(_09059_),
    .B1(_23604_),
    .X(_10368_));
 sky130_fd_sc_hd__and3_1 _37987_ (.A(_10366_),
    .B(_10367_),
    .C(_10368_),
    .X(_10369_));
 sky130_fd_sc_hd__a21oi_1 _37988_ (.A1(_10366_),
    .A2(_10367_),
    .B1(_10368_),
    .Y(_10370_));
 sky130_fd_sc_hd__nor2_1 _37989_ (.A(_10369_),
    .B(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__o21a_1 _37990_ (.A1(_08968_),
    .A2(_10365_),
    .B1(_10371_),
    .X(_10373_));
 sky130_fd_sc_hd__a221oi_4 _37991_ (.A1(_08958_),
    .A2(_08960_),
    .B1(_10364_),
    .B2(_08969_),
    .C1(_10371_),
    .Y(_10374_));
 sky130_fd_sc_hd__o21ai_1 _37992_ (.A1(_10373_),
    .A2(_10374_),
    .B1(_09061_),
    .Y(_10375_));
 sky130_fd_sc_hd__or3_1 _37993_ (.A(_10374_),
    .B(_09061_),
    .C(_10373_),
    .X(_10376_));
 sky130_fd_sc_hd__a211oi_2 _37994_ (.A1(_10375_),
    .A2(_10376_),
    .B1(_08993_),
    .C1(_08994_),
    .Y(_10377_));
 sky130_fd_sc_hd__o211a_2 _37995_ (.A1(_08993_),
    .A2(_08994_),
    .B1(_10375_),
    .C1(_10376_),
    .X(_10378_));
 sky130_fd_sc_hd__o211a_1 _37996_ (.A1(_10377_),
    .A2(_10378_),
    .B1(_09065_),
    .C1(_09067_),
    .X(_10379_));
 sky130_fd_sc_hd__a211oi_4 _37997_ (.A1(_09065_),
    .A2(_09067_),
    .B1(_10377_),
    .C1(_10378_),
    .Y(_10380_));
 sky130_fd_sc_hd__a211oi_2 _37998_ (.A1(_10363_),
    .A2(_09072_),
    .B1(_10379_),
    .C1(_10380_),
    .Y(_10381_));
 sky130_fd_sc_hd__o221a_2 _37999_ (.A1(_10379_),
    .A2(_10380_),
    .B1(_09055_),
    .B2(_09071_),
    .C1(_10363_),
    .X(_10382_));
 sky130_fd_sc_hd__or2_1 _38000_ (.A(_10381_),
    .B(_10382_),
    .X(_10384_));
 sky130_fd_sc_hd__a21o_1 _38001_ (.A1(_09045_),
    .A2(_10362_),
    .B1(_10384_),
    .X(_10385_));
 sky130_fd_sc_hd__buf_2 _38002_ (.A(_10381_),
    .X(_10386_));
 sky130_fd_sc_hd__o211ai_2 _38003_ (.A1(_10386_),
    .A2(_10382_),
    .B1(_09045_),
    .C1(_10362_),
    .Y(_10387_));
 sky130_fd_sc_hd__nand2_1 _38004_ (.A(_10385_),
    .B(_10387_),
    .Y(_10388_));
 sky130_fd_sc_hd__a31o_1 _38005_ (.A1(_09045_),
    .A2(_10362_),
    .A3(_10384_),
    .B1(_10360_),
    .X(_10389_));
 sky130_fd_sc_hd__a21oi_2 _38006_ (.A1(_09045_),
    .A2(_10362_),
    .B1(_10384_),
    .Y(_10390_));
 sky130_fd_sc_hd__o2bb2ai_2 _38007_ (.A1_N(_10360_),
    .A2_N(_10388_),
    .B1(_10389_),
    .B2(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__nand3_1 _38008_ (.A(_10358_),
    .B(_10359_),
    .C(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__a22oi_2 _38009_ (.A1(_08950_),
    .A2(_09114_),
    .B1(_10356_),
    .B2(_10357_),
    .Y(_10393_));
 sky130_fd_sc_hd__nand3b_1 _38010_ (.A_N(_09570_),
    .B(_10282_),
    .C(_10281_),
    .Y(_10395_));
 sky130_fd_sc_hd__a21oi_1 _38011_ (.A1(_10289_),
    .A2(_10395_),
    .B1(_10290_),
    .Y(_10396_));
 sky130_fd_sc_hd__nor2_1 _38012_ (.A(_10396_),
    .B(_10355_),
    .Y(_10397_));
 sky130_fd_sc_hd__o21ai_1 _38013_ (.A1(_10293_),
    .A2(_10292_),
    .B1(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__a22o_1 _38014_ (.A1(_10348_),
    .A2(_10354_),
    .B1(_10291_),
    .B2(_10294_),
    .X(_10399_));
 sky130_fd_sc_hd__nand2_1 _38015_ (.A(_08950_),
    .B(_09114_),
    .Y(_10400_));
 sky130_fd_sc_hd__a21oi_2 _38016_ (.A1(_10398_),
    .A2(_10399_),
    .B1(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__o21bai_1 _38017_ (.A1(_10393_),
    .A2(_10401_),
    .B1_N(_10391_),
    .Y(_10402_));
 sky130_fd_sc_hd__nand3_2 _38018_ (.A(_09113_),
    .B(_10392_),
    .C(_10402_),
    .Y(_10403_));
 sky130_fd_sc_hd__a31oi_1 _38019_ (.A1(_09044_),
    .A2(_09049_),
    .A3(_09050_),
    .B1(_09093_),
    .Y(_10404_));
 sky130_fd_sc_hd__a2bb2oi_1 _38020_ (.A1_N(_10389_),
    .A2_N(_10390_),
    .B1(_10360_),
    .B2(_10388_),
    .Y(_10406_));
 sky130_fd_sc_hd__nand3_1 _38021_ (.A(_10358_),
    .B(_10359_),
    .C(_10406_),
    .Y(_10407_));
 sky130_fd_sc_hd__o21ai_1 _38022_ (.A1(_10393_),
    .A2(_10401_),
    .B1(_10391_),
    .Y(_10408_));
 sky130_fd_sc_hd__o211ai_1 _38023_ (.A1(_09092_),
    .A2(_10404_),
    .B1(_10407_),
    .C1(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__clkbuf_2 _38024_ (.A(_10409_),
    .X(_10410_));
 sky130_fd_sc_hd__a2bb2oi_1 _38025_ (.A1_N(_09110_),
    .A2_N(_09112_),
    .B1(_10403_),
    .B2(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__and4_1 _38026_ (.A(_07611_),
    .B(_07612_),
    .C(_07615_),
    .D(_09081_),
    .X(_10412_));
 sky130_fd_sc_hd__o211a_1 _38027_ (.A1(_09111_),
    .A2(_10412_),
    .B1(_10410_),
    .C1(_10403_),
    .X(_10413_));
 sky130_fd_sc_hd__a21o_1 _38028_ (.A1(_09101_),
    .A2(_09096_),
    .B1(_09091_),
    .X(_10414_));
 sky130_fd_sc_hd__o21ai_1 _38029_ (.A1(_10411_),
    .A2(_10413_),
    .B1(_10414_),
    .Y(_10415_));
 sky130_fd_sc_hd__a2bb2o_1 _38030_ (.A1_N(_09110_),
    .A2_N(_09112_),
    .B1(_10403_),
    .B2(_10409_),
    .X(_10417_));
 sky130_fd_sc_hd__o211ai_1 _38031_ (.A1(_09111_),
    .A2(_10412_),
    .B1(_10410_),
    .C1(_10403_),
    .Y(_10418_));
 sky130_fd_sc_hd__a21oi_1 _38032_ (.A1(_09101_),
    .A2(_09096_),
    .B1(_09091_),
    .Y(_10419_));
 sky130_fd_sc_hd__nand3_1 _38033_ (.A(_10417_),
    .B(_10418_),
    .C(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__nand2_2 _38034_ (.A(_10415_),
    .B(_10420_),
    .Y(_10421_));
 sky130_fd_sc_hd__inv_2 _38035_ (.A(_07640_),
    .Y(_10422_));
 sky130_fd_sc_hd__a21boi_2 _38036_ (.A1(_10422_),
    .A2(_09106_),
    .B1_N(_09107_),
    .Y(_10423_));
 sky130_fd_sc_hd__xor2_4 _38037_ (.A(_10421_),
    .B(_10423_),
    .X(_00011_));
 sky130_fd_sc_hd__a21oi_1 _38038_ (.A1(_10359_),
    .A2(_10406_),
    .B1(_10393_),
    .Y(_10424_));
 sky130_fd_sc_hd__inv_2 _38039_ (.A(_10291_),
    .Y(_10425_));
 sky130_fd_sc_hd__o211a_1 _38040_ (.A1(_09551_),
    .A2(_09555_),
    .B1(_09557_),
    .C1(_09561_),
    .X(_10427_));
 sky130_fd_sc_hd__a32oi_4 _38041_ (.A1(_09564_),
    .A2(_09556_),
    .A3(_09565_),
    .B1(_08176_),
    .B2(_08149_),
    .Y(_10428_));
 sky130_fd_sc_hd__buf_1 _38042_ (.A(_09007_),
    .X(_10429_));
 sky130_fd_sc_hd__nor4b_1 _38043_ (.A(_10324_),
    .B(net248),
    .C(_10322_),
    .D_N(_10429_),
    .Y(_10430_));
 sky130_fd_sc_hd__and4b_1 _38044_ (.A_N(_24251_),
    .B(_07543_),
    .C(_22782_),
    .D(_24286_),
    .X(_10431_));
 sky130_fd_sc_hd__and2_1 _38045_ (.A(_07549_),
    .B(_09541_),
    .X(_10432_));
 sky130_fd_sc_hd__xnor2_1 _38046_ (.A(_08978_),
    .B(_07549_),
    .Y(_10433_));
 sky130_fd_sc_hd__or4bb_2 _38047_ (.A(_10431_),
    .B(_10432_),
    .C_N(_10433_),
    .D_N(_08999_),
    .X(_10434_));
 sky130_fd_sc_hd__buf_1 _38048_ (.A(_10433_),
    .X(_10435_));
 sky130_fd_sc_hd__buf_1 _38049_ (.A(_08999_),
    .X(_10436_));
 sky130_fd_sc_hd__a2bb2o_1 _38050_ (.A1_N(_10431_),
    .A2_N(_10432_),
    .B1(_10435_),
    .B2(_10436_),
    .X(_10438_));
 sky130_fd_sc_hd__o211ai_2 _38051_ (.A1(_09545_),
    .A2(_09546_),
    .B1(_10434_),
    .C1(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__a221o_1 _38052_ (.A1(_08161_),
    .A2(_09543_),
    .B1(_10434_),
    .B2(_10438_),
    .C1(_09546_),
    .X(_10440_));
 sky130_fd_sc_hd__and2_1 _38053_ (.A(_10439_),
    .B(_10440_),
    .X(_10441_));
 sky130_fd_sc_hd__or3_1 _38054_ (.A(net248),
    .B(net195),
    .C(_10441_),
    .X(_10442_));
 sky130_fd_sc_hd__o21ai_2 _38055_ (.A1(net248),
    .A2(net194),
    .B1(_10441_),
    .Y(_10443_));
 sky130_fd_sc_hd__o211a_1 _38056_ (.A1(_08164_),
    .A2(_08167_),
    .B1(_10323_),
    .C1(_10325_),
    .X(_10444_));
 sky130_fd_sc_hd__a221o_1 _38057_ (.A1(_10326_),
    .A2(_10330_),
    .B1(_10442_),
    .B2(_10443_),
    .C1(_10444_),
    .X(_10445_));
 sky130_fd_sc_hd__o211ai_1 _38058_ (.A1(_10444_),
    .A2(_10331_),
    .B1(_10442_),
    .C1(_10443_),
    .Y(_10446_));
 sky130_fd_sc_hd__and2_1 _38059_ (.A(_10445_),
    .B(_10446_),
    .X(_10447_));
 sky130_fd_sc_hd__nor2_1 _38060_ (.A(_07520_),
    .B(_01452_),
    .Y(_10449_));
 sky130_fd_sc_hd__and2_1 _38061_ (.A(_01452_),
    .B(_07520_),
    .X(_10450_));
 sky130_fd_sc_hd__a21boi_1 _38062_ (.A1(_07543_),
    .A2(_07539_),
    .B1_N(_07541_),
    .Y(_10451_));
 sky130_fd_sc_hd__or2_2 _38063_ (.A(_07545_),
    .B(_10451_),
    .X(_10452_));
 sky130_fd_sc_hd__nand2_1 _38064_ (.A(_07550_),
    .B(_10451_),
    .Y(_10453_));
 sky130_fd_sc_hd__nand3b_4 _38065_ (.A_N(_07516_),
    .B(_10452_),
    .C(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__a221o_1 _38066_ (.A1(_25216_),
    .A2(_01448_),
    .B1(_10452_),
    .B2(_10453_),
    .C1(_01447_),
    .X(_10455_));
 sky130_fd_sc_hd__nor3_1 _38067_ (.A(_10302_),
    .B(_10303_),
    .C(_10305_),
    .Y(_10456_));
 sky130_fd_sc_hd__a211o_1 _38068_ (.A1(_10454_),
    .A2(_10455_),
    .B1(_10305_),
    .C1(_10456_),
    .X(_10457_));
 sky130_fd_sc_hd__o211ai_4 _38069_ (.A1(_10305_),
    .A2(net193),
    .B1(_10454_),
    .C1(_10455_),
    .Y(_10458_));
 sky130_fd_sc_hd__and4bb_1 _38070_ (.A_N(_10449_),
    .B_N(_10450_),
    .C(_10457_),
    .D(_10458_),
    .X(_10460_));
 sky130_fd_sc_hd__buf_1 _38071_ (.A(_10449_),
    .X(_10461_));
 sky130_fd_sc_hd__nand2_1 _38072_ (.A(_10457_),
    .B(_10458_),
    .Y(_10462_));
 sky130_fd_sc_hd__o21a_1 _38073_ (.A1(_10461_),
    .A2(_10450_),
    .B1(_10462_),
    .X(_10463_));
 sky130_fd_sc_hd__o211a_1 _38074_ (.A1(_10460_),
    .A2(_10463_),
    .B1(_10311_),
    .C1(_10312_),
    .X(_10464_));
 sky130_fd_sc_hd__a211oi_4 _38075_ (.A1(_10311_),
    .A2(_10312_),
    .B1(_10460_),
    .C1(_10463_),
    .Y(_10465_));
 sky130_fd_sc_hd__nor2_1 _38076_ (.A(_10464_),
    .B(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38077_ (.A(_08959_),
    .X(_10467_));
 sky130_fd_sc_hd__or3b_2 _38078_ (.A(_04558_),
    .B(_25224_),
    .C_N(_10467_),
    .X(_10468_));
 sky130_fd_sc_hd__or2_1 _38079_ (.A(_10467_),
    .B(_10300_),
    .X(_10469_));
 sky130_fd_sc_hd__and3_1 _38080_ (.A(_10466_),
    .B(_10468_),
    .C(_10469_),
    .X(_10471_));
 sky130_fd_sc_hd__o2bb2a_1 _38081_ (.A1_N(_10469_),
    .A2_N(_10468_),
    .B1(_10464_),
    .B2(_10465_),
    .X(_10472_));
 sky130_fd_sc_hd__nor2_2 _38082_ (.A(_10471_),
    .B(_10472_),
    .Y(_10473_));
 sky130_fd_sc_hd__xnor2_1 _38083_ (.A(_10447_),
    .B(_10473_),
    .Y(_10474_));
 sky130_fd_sc_hd__o21bai_4 _38084_ (.A1(_10427_),
    .A2(_10428_),
    .B1_N(_10474_),
    .Y(_10475_));
 sky130_fd_sc_hd__o21ai_1 _38085_ (.A1(_08177_),
    .A2(_10287_),
    .B1(_09566_),
    .Y(_10476_));
 sky130_fd_sc_hd__nand3_1 _38086_ (.A(_09562_),
    .B(_10476_),
    .C(_10474_),
    .Y(_10477_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38087_ (.A(_10477_),
    .X(_10478_));
 sky130_fd_sc_hd__a21o_1 _38088_ (.A1(_10336_),
    .A2(_10338_),
    .B1(_10335_),
    .X(_10479_));
 sky130_fd_sc_hd__a21oi_1 _38089_ (.A1(_10475_),
    .A2(_10478_),
    .B1(_10479_),
    .Y(_10480_));
 sky130_fd_sc_hd__inv_2 _38090_ (.A(_10337_),
    .Y(_10482_));
 sky130_fd_sc_hd__o211a_1 _38091_ (.A1(_10335_),
    .A2(_10482_),
    .B1(_10475_),
    .C1(_10477_),
    .X(_10483_));
 sky130_fd_sc_hd__nor2_1 _38092_ (.A(_10480_),
    .B(_10483_),
    .Y(_10484_));
 sky130_fd_sc_hd__o21a_1 _38093_ (.A1(_09538_),
    .A2(_09530_),
    .B1(_09535_),
    .X(_10485_));
 sky130_fd_sc_hd__a31o_1 _38094_ (.A1(_09523_),
    .A2(_08130_),
    .A3(_09511_),
    .B1(_09519_),
    .X(_10486_));
 sky130_fd_sc_hd__a21o_1 _38095_ (.A1(_09728_),
    .A2(_09735_),
    .B1(_09718_),
    .X(_10487_));
 sky130_fd_sc_hd__o21ai_4 _38096_ (.A1(_09728_),
    .A2(_09735_),
    .B1(_10487_),
    .Y(_10488_));
 sky130_fd_sc_hd__o21a_1 _38097_ (.A1(_09498_),
    .A2(_09502_),
    .B1(_09504_),
    .X(_10489_));
 sky130_fd_sc_hd__a21oi_1 _38098_ (.A1(_09523_),
    .A2(_09508_),
    .B1(_10489_),
    .Y(_10490_));
 sky130_fd_sc_hd__nand4_1 _38099_ (.A(_08109_),
    .B(_09523_),
    .C(_09505_),
    .D(_09508_),
    .Y(_10491_));
 sky130_fd_sc_hd__a21oi_1 _38100_ (.A1(_07649_),
    .A2(_08120_),
    .B1(_10491_),
    .Y(_10493_));
 sky130_fd_sc_hd__a32o_1 _38101_ (.A1(_09119_),
    .A2(_09333_),
    .A3(_09336_),
    .B1(_09343_),
    .B2(_09438_),
    .X(_10494_));
 sky130_fd_sc_hd__nor2_1 _38102_ (.A(_09323_),
    .B(_09324_),
    .Y(_10495_));
 sky130_fd_sc_hd__a32o_1 _38103_ (.A1(_09221_),
    .A2(_09311_),
    .A3(_09314_),
    .B1(_09321_),
    .B2(_10495_),
    .X(_10496_));
 sky130_fd_sc_hd__and3_1 _38104_ (.A(_09213_),
    .B(_09200_),
    .C(_09199_),
    .X(_10497_));
 sky130_fd_sc_hd__a31o_1 _38105_ (.A1(_09224_),
    .A2(_09225_),
    .A3(_09227_),
    .B1(_09312_),
    .X(_10498_));
 sky130_fd_sc_hd__buf_1 _38106_ (.A(_07729_),
    .X(_10499_));
 sky130_fd_sc_hd__clkbuf_2 _38107_ (.A(_07728_),
    .X(_10500_));
 sky130_fd_sc_hd__and4_1 _38108_ (.A(_07884_),
    .B(_10499_),
    .C(_10500_),
    .D(_07730_),
    .X(_10501_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38109_ (.A(_09203_),
    .X(_10502_));
 sky130_fd_sc_hd__and4bb_1 _38110_ (.A_N(_07891_),
    .B_N(_09207_),
    .C(_10502_),
    .D(_25373_),
    .X(_10504_));
 sky130_fd_sc_hd__or2b_1 _38111_ (.A(_07730_),
    .B_N(_09203_),
    .X(_10505_));
 sky130_fd_sc_hd__or4_1 _38112_ (.A(_07891_),
    .B(_03131_),
    .C(_10499_),
    .D(_10505_),
    .X(_10506_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38113_ (.A(_03131_),
    .X(_10507_));
 sky130_fd_sc_hd__a2bb2o_1 _38114_ (.A1_N(_10507_),
    .A2_N(_10499_),
    .B1(_01529_),
    .B2(_09204_),
    .X(_10508_));
 sky130_fd_sc_hd__o211a_1 _38115_ (.A1(_10501_),
    .A2(_10504_),
    .B1(_10506_),
    .C1(_10508_),
    .X(_10509_));
 sky130_fd_sc_hd__a211oi_1 _38116_ (.A1(_10506_),
    .A2(_10508_),
    .B1(_10501_),
    .C1(_10504_),
    .Y(_10510_));
 sky130_fd_sc_hd__nor2_1 _38117_ (.A(_04844_),
    .B(_07869_),
    .Y(_10511_));
 sky130_fd_sc_hd__nor2_1 _38118_ (.A(_07695_),
    .B(_23762_),
    .Y(_10512_));
 sky130_fd_sc_hd__or3_2 _38119_ (.A(_09193_),
    .B(_10511_),
    .C(_10512_),
    .X(_10513_));
 sky130_fd_sc_hd__a2bb2o_1 _38120_ (.A1_N(_10511_),
    .A2_N(_10512_),
    .B1(_01702_),
    .B2(_07867_),
    .X(_10515_));
 sky130_fd_sc_hd__and4_1 _38121_ (.A(_06341_),
    .B(_10513_),
    .C(_10515_),
    .D(_09154_),
    .X(_10516_));
 sky130_fd_sc_hd__o2bb2a_1 _38122_ (.A1_N(_10513_),
    .A2_N(_10515_),
    .B1(_01694_),
    .B2(_07878_),
    .X(_10517_));
 sky130_fd_sc_hd__nor2_1 _38123_ (.A(_03283_),
    .B(_07861_),
    .Y(_10518_));
 sky130_fd_sc_hd__and2_1 _38124_ (.A(_03281_),
    .B(_07861_),
    .X(_10519_));
 sky130_fd_sc_hd__nor2_1 _38125_ (.A(_10518_),
    .B(_10519_),
    .Y(_10520_));
 sky130_fd_sc_hd__or2_1 _38126_ (.A(_09202_),
    .B(_10520_),
    .X(_10521_));
 sky130_fd_sc_hd__or3b_1 _38127_ (.A(_10518_),
    .B(_10519_),
    .C_N(_09202_),
    .X(_10522_));
 sky130_fd_sc_hd__nand2_1 _38128_ (.A(_10521_),
    .B(_10522_),
    .Y(_10523_));
 sky130_fd_sc_hd__nor2_1 _38129_ (.A(_09196_),
    .B(_10523_),
    .Y(_10524_));
 sky130_fd_sc_hd__buf_1 _38130_ (.A(_06364_),
    .X(_10526_));
 sky130_fd_sc_hd__clkbuf_2 _38131_ (.A(_10526_),
    .X(_10527_));
 sky130_fd_sc_hd__a32oi_1 _38132_ (.A1(_10527_),
    .A2(_09192_),
    .A3(_09193_),
    .B1(_10521_),
    .B2(_10522_),
    .Y(_10528_));
 sky130_fd_sc_hd__or4_1 _38133_ (.A(_10516_),
    .B(_10517_),
    .C(_10524_),
    .D(_10528_),
    .X(_10529_));
 sky130_fd_sc_hd__o22ai_1 _38134_ (.A1(_10516_),
    .A2(_10517_),
    .B1(_10524_),
    .B2(_10528_),
    .Y(_10530_));
 sky130_fd_sc_hd__or4bb_1 _38135_ (.A(_10509_),
    .B(_10510_),
    .C_N(_10529_),
    .D_N(_10530_),
    .X(_10531_));
 sky130_fd_sc_hd__a2bb2o_1 _38136_ (.A1_N(_10509_),
    .A2_N(_10510_),
    .B1(_10529_),
    .B2(_10530_),
    .X(_10532_));
 sky130_fd_sc_hd__nand2_1 _38137_ (.A(_10531_),
    .B(_10532_),
    .Y(_10533_));
 sky130_fd_sc_hd__xor2_1 _38138_ (.A(_10498_),
    .B(_10533_),
    .X(_10534_));
 sky130_fd_sc_hd__o21ba_2 _38139_ (.A1(_09211_),
    .A2(_10497_),
    .B1_N(_10534_),
    .X(_10535_));
 sky130_fd_sc_hd__nor3b_2 _38140_ (.A(_09211_),
    .B(_10497_),
    .C_N(_10534_),
    .Y(_10537_));
 sky130_fd_sc_hd__nand2_1 _38141_ (.A(_09288_),
    .B(_09303_),
    .Y(_10538_));
 sky130_fd_sc_hd__a21o_1 _38142_ (.A1(_09292_),
    .A2(_09289_),
    .B1(_09276_),
    .X(_10539_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38143_ (.A(_07807_),
    .X(_10540_));
 sky130_fd_sc_hd__buf_1 _38144_ (.A(_10540_),
    .X(_10541_));
 sky130_fd_sc_hd__and3_1 _38145_ (.A(_06272_),
    .B(_10541_),
    .C(_04734_),
    .X(_10542_));
 sky130_fd_sc_hd__nand2_1 _38146_ (.A(_06266_),
    .B(_10540_),
    .Y(_10543_));
 sky130_fd_sc_hd__nand2_1 _38147_ (.A(_06272_),
    .B(_09278_),
    .Y(_10544_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38148_ (.A(_09278_),
    .X(_10545_));
 sky130_fd_sc_hd__o2bb2a_1 _38149_ (.A1_N(_10543_),
    .A2_N(_10544_),
    .B1(_04745_),
    .B2(_10545_),
    .X(_10546_));
 sky130_fd_sc_hd__and2_1 _38150_ (.A(_09233_),
    .B(\delay_line[4][15] ),
    .X(_10548_));
 sky130_fd_sc_hd__buf_1 _38151_ (.A(\delay_line[4][15] ),
    .X(_10549_));
 sky130_fd_sc_hd__nor2_1 _38152_ (.A(_10549_),
    .B(_09233_),
    .Y(_10550_));
 sky130_fd_sc_hd__nor2_1 _38153_ (.A(_10548_),
    .B(_10550_),
    .Y(_10551_));
 sky130_fd_sc_hd__and3b_1 _38154_ (.A_N(_06225_),
    .B(\delay_line[4][13] ),
    .C(_09236_),
    .X(_10552_));
 sky130_fd_sc_hd__a21oi_1 _38155_ (.A1(_07767_),
    .A2(net432),
    .B1(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__xor2_1 _38156_ (.A(_10551_),
    .B(_10553_),
    .X(_10554_));
 sky130_fd_sc_hd__clkbuf_4 _38157_ (.A(_10554_),
    .X(_10555_));
 sky130_fd_sc_hd__inv_2 _38158_ (.A(net432),
    .Y(_10556_));
 sky130_fd_sc_hd__clkbuf_2 _38159_ (.A(_10556_),
    .X(_10557_));
 sky130_fd_sc_hd__or4b_4 _38160_ (.A(_04701_),
    .B(_07767_),
    .C(_10557_),
    .D_N(_07771_),
    .X(_10559_));
 sky130_fd_sc_hd__nand3_4 _38161_ (.A(_09264_),
    .B(_10555_),
    .C(_10559_),
    .Y(_10560_));
 sky130_fd_sc_hd__and4b_2 _38162_ (.A_N(_04701_),
    .B(\delay_line[4][12] ),
    .C(net432),
    .D(_07771_),
    .X(_10561_));
 sky130_fd_sc_hd__o21bai_4 _38163_ (.A1(_09245_),
    .A2(_10561_),
    .B1_N(_10555_),
    .Y(_10562_));
 sky130_fd_sc_hd__nor3_1 _38164_ (.A(_07752_),
    .B(_07753_),
    .C(_09251_),
    .Y(_10563_));
 sky130_fd_sc_hd__nand2_1 _38165_ (.A(_07763_),
    .B(net178),
    .Y(_10564_));
 sky130_fd_sc_hd__or3b_1 _38166_ (.A(_07746_),
    .B(_09246_),
    .C_N(_09247_),
    .X(_10565_));
 sky130_fd_sc_hd__o31a_2 _38167_ (.A1(_09246_),
    .A2(_07748_),
    .A3(_09249_),
    .B1(_10565_),
    .X(_10566_));
 sky130_fd_sc_hd__clkbuf_2 _38168_ (.A(\delay_line[11][11] ),
    .X(_10567_));
 sky130_fd_sc_hd__inv_2 _38169_ (.A(net408),
    .Y(_10568_));
 sky130_fd_sc_hd__or2_2 _38170_ (.A(_10567_),
    .B(_10568_),
    .X(_10570_));
 sky130_fd_sc_hd__nand3b_1 _38171_ (.A_N(_06233_),
    .B(net409),
    .C(_09247_),
    .Y(_10571_));
 sky130_fd_sc_hd__xor2_2 _38172_ (.A(\delay_line[11][12] ),
    .B(net408),
    .X(_10572_));
 sky130_fd_sc_hd__a21oi_1 _38173_ (.A1(_10570_),
    .A2(_10571_),
    .B1(_10572_),
    .Y(_10573_));
 sky130_fd_sc_hd__and3_1 _38174_ (.A(_10570_),
    .B(_10571_),
    .C(_10572_),
    .X(_10574_));
 sky130_fd_sc_hd__or2_2 _38175_ (.A(_10573_),
    .B(_10574_),
    .X(_10575_));
 sky130_fd_sc_hd__a21oi_4 _38176_ (.A1(_10564_),
    .A2(_10566_),
    .B1(_10575_),
    .Y(_10576_));
 sky130_fd_sc_hd__and3_1 _38177_ (.A(_10575_),
    .B(_10564_),
    .C(_10566_),
    .X(_10577_));
 sky130_fd_sc_hd__o2bb2ai_4 _38178_ (.A1_N(_10560_),
    .A2_N(_10562_),
    .B1(_10576_),
    .B2(_10577_),
    .Y(_10578_));
 sky130_fd_sc_hd__inv_2 _38179_ (.A(net178),
    .Y(_10579_));
 sky130_fd_sc_hd__nor2_1 _38180_ (.A(_10579_),
    .B(_07759_),
    .Y(_10581_));
 sky130_fd_sc_hd__nand2_1 _38181_ (.A(_10566_),
    .B(_10575_),
    .Y(_10582_));
 sky130_fd_sc_hd__inv_2 _38182_ (.A(_10566_),
    .Y(_10583_));
 sky130_fd_sc_hd__o21bai_1 _38183_ (.A1(_10579_),
    .A2(_07759_),
    .B1_N(_10583_),
    .Y(_10584_));
 sky130_fd_sc_hd__inv_2 _38184_ (.A(_10575_),
    .Y(_10585_));
 sky130_fd_sc_hd__nand2_1 _38185_ (.A(_10584_),
    .B(_10585_),
    .Y(_10586_));
 sky130_fd_sc_hd__o21ai_1 _38186_ (.A1(_10581_),
    .A2(_10582_),
    .B1(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__a31oi_4 _38187_ (.A1(_09264_),
    .A2(_10555_),
    .A3(_10559_),
    .B1(_10587_),
    .Y(_10588_));
 sky130_fd_sc_hd__nand2_1 _38188_ (.A(_10588_),
    .B(_10562_),
    .Y(_10589_));
 sky130_fd_sc_hd__o21ai_1 _38189_ (.A1(_07786_),
    .A2(_09269_),
    .B1(_09262_),
    .Y(_10590_));
 sky130_fd_sc_hd__a21o_2 _38190_ (.A1(_10578_),
    .A2(_10589_),
    .B1(_10590_),
    .X(_10592_));
 sky130_fd_sc_hd__a31oi_4 _38191_ (.A1(_09267_),
    .A2(_09264_),
    .A3(_09257_),
    .B1(_07786_),
    .Y(_10593_));
 sky130_fd_sc_hd__a21oi_2 _38192_ (.A1(_09264_),
    .A2(_10559_),
    .B1(_10555_),
    .Y(_10594_));
 sky130_fd_sc_hd__o21a_1 _38193_ (.A1(_10581_),
    .A2(_10582_),
    .B1(_10586_),
    .X(_10595_));
 sky130_fd_sc_hd__nand2_2 _38194_ (.A(_10560_),
    .B(_10595_),
    .Y(_10596_));
 sky130_fd_sc_hd__o221ai_4 _38195_ (.A1(_09268_),
    .A2(_10593_),
    .B1(_10594_),
    .B2(_10596_),
    .C1(_10578_),
    .Y(_10597_));
 sky130_fd_sc_hd__buf_2 _38196_ (.A(_07786_),
    .X(_10598_));
 sky130_fd_sc_hd__o21a_1 _38197_ (.A1(_09245_),
    .A2(_09258_),
    .B1(_09262_),
    .X(_10599_));
 sky130_fd_sc_hd__o21ai_4 _38198_ (.A1(_10598_),
    .A2(_10599_),
    .B1(_09263_),
    .Y(_10600_));
 sky130_fd_sc_hd__a21oi_4 _38199_ (.A1(_10592_),
    .A2(_10597_),
    .B1(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__o2bb2ai_4 _38200_ (.A1_N(_10562_),
    .A2_N(_10588_),
    .B1(_09268_),
    .B2(_10593_),
    .Y(_10603_));
 sky130_fd_sc_hd__a21oi_4 _38201_ (.A1(_10560_),
    .A2(_10562_),
    .B1(_10595_),
    .Y(_10604_));
 sky130_fd_sc_hd__o211a_1 _38202_ (.A1(_10603_),
    .A2(_10604_),
    .B1(_10600_),
    .C1(_10592_),
    .X(_10605_));
 sky130_fd_sc_hd__o22ai_2 _38203_ (.A1(_10542_),
    .A2(_10546_),
    .B1(_10601_),
    .B2(_10605_),
    .Y(_10606_));
 sky130_fd_sc_hd__clkbuf_2 _38204_ (.A(_06266_),
    .X(_10607_));
 sky130_fd_sc_hd__buf_1 _38205_ (.A(_10540_),
    .X(_10608_));
 sky130_fd_sc_hd__a22o_1 _38206_ (.A1(_04734_),
    .A2(_10608_),
    .B1(_10543_),
    .B2(_10544_),
    .X(_10609_));
 sky130_fd_sc_hd__a21oi_1 _38207_ (.A1(_10578_),
    .A2(_10589_),
    .B1(_10590_),
    .Y(_10610_));
 sky130_fd_sc_hd__nor2_1 _38208_ (.A(_10604_),
    .B(_10603_),
    .Y(_10611_));
 sky130_fd_sc_hd__o21bai_2 _38209_ (.A1(_10610_),
    .A2(_10611_),
    .B1_N(_10600_),
    .Y(_10612_));
 sky130_fd_sc_hd__o211ai_4 _38210_ (.A1(_10603_),
    .A2(_10604_),
    .B1(_10600_),
    .C1(_10592_),
    .Y(_10614_));
 sky130_fd_sc_hd__o2111ai_4 _38211_ (.A1(_10607_),
    .A2(_09277_),
    .B1(_10609_),
    .C1(_10612_),
    .D1(_10614_),
    .Y(_10615_));
 sky130_fd_sc_hd__nand3_2 _38212_ (.A(_10539_),
    .B(_10606_),
    .C(_10615_),
    .Y(_10616_));
 sky130_fd_sc_hd__o21a_1 _38213_ (.A1(_10607_),
    .A2(_09277_),
    .B1(_10609_),
    .X(_10617_));
 sky130_fd_sc_hd__o21ai_1 _38214_ (.A1(_10601_),
    .A2(_10605_),
    .B1(_10617_),
    .Y(_10618_));
 sky130_fd_sc_hd__a21oi_1 _38215_ (.A1(_09292_),
    .A2(_09289_),
    .B1(_09276_),
    .Y(_10619_));
 sky130_fd_sc_hd__o211ai_1 _38216_ (.A1(_10542_),
    .A2(_10546_),
    .B1(_10612_),
    .C1(_10614_),
    .Y(_10620_));
 sky130_fd_sc_hd__nand3_1 _38217_ (.A(_10618_),
    .B(_10619_),
    .C(_10620_),
    .Y(_10621_));
 sky130_fd_sc_hd__clkbuf_2 _38218_ (.A(_10621_),
    .X(_10622_));
 sky130_fd_sc_hd__xnor2_1 _38219_ (.A(_03148_),
    .B(_10540_),
    .Y(_10623_));
 sky130_fd_sc_hd__and4b_1 _38220_ (.A_N(_03148_),
    .B(_04745_),
    .C(_07807_),
    .D(_03206_),
    .X(_10625_));
 sky130_fd_sc_hd__a21oi_1 _38221_ (.A1(_09281_),
    .A2(_10623_),
    .B1(_10625_),
    .Y(_10626_));
 sky130_fd_sc_hd__and3_2 _38222_ (.A(_04762_),
    .B(_10608_),
    .C(_10626_),
    .X(_10627_));
 sky130_fd_sc_hd__clkbuf_2 _38223_ (.A(_10541_),
    .X(_10628_));
 sky130_fd_sc_hd__a21oi_2 _38224_ (.A1(_04789_),
    .A2(_10628_),
    .B1(_10626_),
    .Y(_10629_));
 sky130_fd_sc_hd__o2bb2ai_2 _38225_ (.A1_N(_10616_),
    .A2_N(_10622_),
    .B1(_10627_),
    .B2(_10629_),
    .Y(_10630_));
 sky130_fd_sc_hd__nor2_1 _38226_ (.A(_10627_),
    .B(_10629_),
    .Y(_10631_));
 sky130_fd_sc_hd__nand3_2 _38227_ (.A(_10616_),
    .B(_10622_),
    .C(_10631_),
    .Y(_10632_));
 sky130_fd_sc_hd__nand3_2 _38228_ (.A(_10538_),
    .B(_10630_),
    .C(_10632_),
    .Y(_10633_));
 sky130_fd_sc_hd__a21bo_1 _38229_ (.A1(_10616_),
    .A2(_10621_),
    .B1_N(_10631_),
    .X(_10634_));
 sky130_fd_sc_hd__o211ai_2 _38230_ (.A1(_10627_),
    .A2(_10629_),
    .B1(_10616_),
    .C1(_10622_),
    .Y(_10636_));
 sky130_fd_sc_hd__and2_1 _38231_ (.A(_09288_),
    .B(_09303_),
    .X(_10637_));
 sky130_fd_sc_hd__nand3_4 _38232_ (.A(_10634_),
    .B(_10636_),
    .C(_10637_),
    .Y(_10638_));
 sky130_fd_sc_hd__or3_1 _38233_ (.A(_04786_),
    .B(_03206_),
    .C(_06280_),
    .X(_10639_));
 sky130_fd_sc_hd__buf_2 _38234_ (.A(_06287_),
    .X(_10640_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38235_ (.A(_03221_),
    .X(_10641_));
 sky130_fd_sc_hd__nand4_1 _38236_ (.A(_09298_),
    .B(_10640_),
    .C(_10641_),
    .D(_10639_),
    .Y(_10642_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38237_ (.A(_06200_),
    .X(_10643_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38238_ (.A(_10499_),
    .X(_10644_));
 sky130_fd_sc_hd__and2_1 _38239_ (.A(_10643_),
    .B(_10644_),
    .X(_10645_));
 sky130_fd_sc_hd__o21a_2 _38240_ (.A1(_07888_),
    .A2(_10645_),
    .B1(_10641_),
    .X(_10647_));
 sky130_fd_sc_hd__clkbuf_2 _38241_ (.A(_07888_),
    .X(_10648_));
 sky130_fd_sc_hd__nor3_1 _38242_ (.A(_10641_),
    .B(_10648_),
    .C(_10645_),
    .Y(_10649_));
 sky130_fd_sc_hd__a211o_1 _38243_ (.A1(_10639_),
    .A2(_10642_),
    .B1(_10647_),
    .C1(_10649_),
    .X(_10650_));
 sky130_fd_sc_hd__o211ai_2 _38244_ (.A1(_10647_),
    .A2(_10649_),
    .B1(_10639_),
    .C1(_10642_),
    .Y(_10651_));
 sky130_fd_sc_hd__nand2_1 _38245_ (.A(_10650_),
    .B(_10651_),
    .Y(_10652_));
 sky130_fd_sc_hd__and2_1 _38246_ (.A(_09224_),
    .B(_10652_),
    .X(_10653_));
 sky130_fd_sc_hd__o2111a_1 _38247_ (.A1(_09222_),
    .A2(_09223_),
    .B1(_10651_),
    .C1(_01537_),
    .D1(_10650_),
    .X(_10654_));
 sky130_fd_sc_hd__o2bb2ai_2 _38248_ (.A1_N(_10633_),
    .A2_N(_10638_),
    .B1(_10653_),
    .B2(_10654_),
    .Y(_10655_));
 sky130_fd_sc_hd__a21oi_2 _38249_ (.A1(_09224_),
    .A2(_10652_),
    .B1(_10654_),
    .Y(_10656_));
 sky130_fd_sc_hd__nand3_2 _38250_ (.A(_10633_),
    .B(_10638_),
    .C(_10656_),
    .Y(_10658_));
 sky130_fd_sc_hd__nand2_2 _38251_ (.A(_09306_),
    .B(_09311_),
    .Y(_10659_));
 sky130_fd_sc_hd__a21oi_2 _38252_ (.A1(_10655_),
    .A2(_10658_),
    .B1(_10659_),
    .Y(_10660_));
 sky130_fd_sc_hd__a21oi_2 _38253_ (.A1(_10633_),
    .A2(_10638_),
    .B1(_10656_),
    .Y(_10661_));
 sky130_fd_sc_hd__nand2_1 _38254_ (.A(_10658_),
    .B(_10659_),
    .Y(_10662_));
 sky130_fd_sc_hd__nor2_2 _38255_ (.A(_10661_),
    .B(_10662_),
    .Y(_10663_));
 sky130_fd_sc_hd__o22ai_2 _38256_ (.A1(_10535_),
    .A2(_10537_),
    .B1(_10660_),
    .B2(_10663_),
    .Y(_10664_));
 sky130_fd_sc_hd__or2_2 _38257_ (.A(_10535_),
    .B(_10537_),
    .X(_10665_));
 sky130_fd_sc_hd__a21o_1 _38258_ (.A1(_10655_),
    .A2(_10658_),
    .B1(_10659_),
    .X(_10666_));
 sky130_fd_sc_hd__nand3_1 _38259_ (.A(_10655_),
    .B(_10658_),
    .C(_10659_),
    .Y(_10667_));
 sky130_fd_sc_hd__nand3b_1 _38260_ (.A_N(_10665_),
    .B(_10666_),
    .C(_10667_),
    .Y(_10669_));
 sky130_fd_sc_hd__nand3_2 _38261_ (.A(_10496_),
    .B(_10664_),
    .C(_10669_),
    .Y(_10670_));
 sky130_fd_sc_hd__o21bai_4 _38262_ (.A1(_10660_),
    .A2(_10663_),
    .B1_N(_10665_),
    .Y(_10671_));
 sky130_fd_sc_hd__o221ai_4 _38263_ (.A1(_10535_),
    .A2(_10537_),
    .B1(_10661_),
    .B2(_10662_),
    .C1(_10666_),
    .Y(_10672_));
 sky130_fd_sc_hd__a32oi_4 _38264_ (.A1(_09221_),
    .A2(_09311_),
    .A3(_09314_),
    .B1(_09321_),
    .B2(_10495_),
    .Y(_10673_));
 sky130_fd_sc_hd__nand3_4 _38265_ (.A(_10671_),
    .B(_10672_),
    .C(_10673_),
    .Y(_10674_));
 sky130_fd_sc_hd__o21a_1 _38266_ (.A1(_09152_),
    .A2(_09169_),
    .B1(_09167_),
    .X(_10675_));
 sky130_fd_sc_hd__o21a_2 _38267_ (.A1(_09183_),
    .A2(_09218_),
    .B1(_09216_),
    .X(_10676_));
 sky130_fd_sc_hd__buf_1 _38268_ (.A(_09121_),
    .X(_10677_));
 sky130_fd_sc_hd__nor2_1 _38269_ (.A(_01788_),
    .B(_23970_),
    .Y(_10678_));
 sky130_fd_sc_hd__and3_1 _38270_ (.A(_23974_),
    .B(_10677_),
    .C(_10678_),
    .X(_10680_));
 sky130_fd_sc_hd__a21oi_1 _38271_ (.A1(_25337_),
    .A2(_09128_),
    .B1(_07703_),
    .Y(_10681_));
 sky130_fd_sc_hd__a31o_1 _38272_ (.A1(_23976_),
    .A2(_09128_),
    .A3(_01789_),
    .B1(_10681_),
    .X(_10682_));
 sky130_fd_sc_hd__nand2_1 _38273_ (.A(_10682_),
    .B(_03349_),
    .Y(_10683_));
 sky130_fd_sc_hd__a311o_1 _38274_ (.A1(_23976_),
    .A2(_10677_),
    .A3(_01789_),
    .B1(_03349_),
    .C1(_10681_),
    .X(_10684_));
 sky130_fd_sc_hd__o211a_1 _38275_ (.A1(_09132_),
    .A2(_10680_),
    .B1(_10683_),
    .C1(_10684_),
    .X(_10685_));
 sky130_fd_sc_hd__a211oi_2 _38276_ (.A1(_10684_),
    .A2(_10683_),
    .B1(_10680_),
    .C1(_09132_),
    .Y(_10686_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38277_ (.A(_06430_),
    .X(_10687_));
 sky130_fd_sc_hd__nand2_1 _38278_ (.A(_09141_),
    .B(_10687_),
    .Y(_10688_));
 sky130_fd_sc_hd__a21oi_1 _38279_ (.A1(_01740_),
    .A2(_06430_),
    .B1(_01741_),
    .Y(_10689_));
 sky130_fd_sc_hd__and3_1 _38280_ (.A(_01740_),
    .B(_01741_),
    .C(_06428_),
    .X(_10691_));
 sky130_fd_sc_hd__a21bo_1 _38281_ (.A1(_01757_),
    .A2(_09122_),
    .B1_N(_09123_),
    .X(_10692_));
 sky130_fd_sc_hd__or3_1 _38282_ (.A(_10689_),
    .B(_10691_),
    .C(_10692_),
    .X(_10693_));
 sky130_fd_sc_hd__o21ai_2 _38283_ (.A1(_10689_),
    .A2(_10691_),
    .B1(_10692_),
    .Y(_10694_));
 sky130_fd_sc_hd__or4bb_2 _38284_ (.A(_04642_),
    .B(_10688_),
    .C_N(_10693_),
    .D_N(_10694_),
    .X(_10695_));
 sky130_fd_sc_hd__a2bb2o_1 _38285_ (.A1_N(_10688_),
    .A2_N(_04642_),
    .B1(_10694_),
    .B2(_10693_),
    .X(_10696_));
 sky130_fd_sc_hd__nand2_1 _38286_ (.A(_10695_),
    .B(_10696_),
    .Y(_10697_));
 sky130_fd_sc_hd__o21ai_1 _38287_ (.A1(_10685_),
    .A2(_10686_),
    .B1(_10697_),
    .Y(_10698_));
 sky130_fd_sc_hd__inv_2 _38288_ (.A(_10698_),
    .Y(_10699_));
 sky130_fd_sc_hd__nor3_1 _38289_ (.A(_10685_),
    .B(_10686_),
    .C(_10697_),
    .Y(_10700_));
 sky130_fd_sc_hd__o21ai_4 _38290_ (.A1(_09165_),
    .A2(_09164_),
    .B1(_09163_),
    .Y(_10702_));
 sky130_fd_sc_hd__nand3b_1 _38291_ (.A_N(_07862_),
    .B(_09194_),
    .C(_09196_),
    .Y(_10703_));
 sky130_fd_sc_hd__nor2_1 _38292_ (.A(net417),
    .B(_07695_),
    .Y(_10704_));
 sky130_fd_sc_hd__clkbuf_2 _38293_ (.A(\delay_line[9][12] ),
    .X(_10705_));
 sky130_fd_sc_hd__a21boi_1 _38294_ (.A1(_09188_),
    .A2(_07871_),
    .B1_N(_09189_),
    .Y(_10706_));
 sky130_fd_sc_hd__a21o_1 _38295_ (.A1(_10705_),
    .A2(_07695_),
    .B1(_10706_),
    .X(_10707_));
 sky130_fd_sc_hd__nor2_1 _38296_ (.A(_03265_),
    .B(_07869_),
    .Y(_10708_));
 sky130_fd_sc_hd__o21ai_1 _38297_ (.A1(_10708_),
    .A2(_10704_),
    .B1(_10706_),
    .Y(_10709_));
 sky130_fd_sc_hd__o21a_1 _38298_ (.A1(_10704_),
    .A2(_10707_),
    .B1(_10709_),
    .X(_10710_));
 sky130_fd_sc_hd__xnor2_1 _38299_ (.A(_09155_),
    .B(_10710_),
    .Y(_10711_));
 sky130_fd_sc_hd__and3_1 _38300_ (.A(_10703_),
    .B(_09199_),
    .C(_10711_),
    .X(_10713_));
 sky130_fd_sc_hd__a21o_1 _38301_ (.A1(_10703_),
    .A2(_09199_),
    .B1(_10711_),
    .X(_10714_));
 sky130_fd_sc_hd__and2b_1 _38302_ (.A_N(_10713_),
    .B(_10714_),
    .X(_10715_));
 sky130_fd_sc_hd__or3_2 _38303_ (.A(_09158_),
    .B(_09160_),
    .C(_10715_),
    .X(_10716_));
 sky130_fd_sc_hd__o21ai_4 _38304_ (.A1(_09158_),
    .A2(_09160_),
    .B1(_10715_),
    .Y(_10717_));
 sky130_fd_sc_hd__and2_1 _38305_ (.A(_10716_),
    .B(_10717_),
    .X(_10718_));
 sky130_fd_sc_hd__xnor2_1 _38306_ (.A(_10702_),
    .B(_10718_),
    .Y(_10719_));
 sky130_fd_sc_hd__o21a_1 _38307_ (.A1(_10699_),
    .A2(_10700_),
    .B1(_10719_),
    .X(_10720_));
 sky130_fd_sc_hd__nor3_1 _38308_ (.A(_10699_),
    .B(_10700_),
    .C(_10719_),
    .Y(_10721_));
 sky130_fd_sc_hd__buf_2 _38309_ (.A(_10721_),
    .X(_10722_));
 sky130_fd_sc_hd__nor3_4 _38310_ (.A(_10676_),
    .B(_10720_),
    .C(_10722_),
    .Y(_10724_));
 sky130_fd_sc_hd__o21ai_1 _38311_ (.A1(_10720_),
    .A2(_10721_),
    .B1(_10676_),
    .Y(_10725_));
 sky130_fd_sc_hd__inv_2 _38312_ (.A(_10725_),
    .Y(_10726_));
 sky130_fd_sc_hd__nor3_4 _38313_ (.A(_10675_),
    .B(_10724_),
    .C(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__o21a_1 _38314_ (.A1(_10724_),
    .A2(_10726_),
    .B1(_10675_),
    .X(_10728_));
 sky130_fd_sc_hd__o2bb2ai_4 _38315_ (.A1_N(_10670_),
    .A2_N(_10674_),
    .B1(_10727_),
    .B2(_10728_),
    .Y(_10729_));
 sky130_fd_sc_hd__nor2_2 _38316_ (.A(_10727_),
    .B(_10728_),
    .Y(_10730_));
 sky130_fd_sc_hd__nand3_4 _38317_ (.A(_10670_),
    .B(_10674_),
    .C(_10730_),
    .Y(_10731_));
 sky130_fd_sc_hd__nand2_2 _38318_ (.A(_09328_),
    .B(_09333_),
    .Y(_10732_));
 sky130_fd_sc_hd__a21oi_2 _38319_ (.A1(_10729_),
    .A2(_10731_),
    .B1(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__inv_2 _38320_ (.A(_10730_),
    .Y(_10735_));
 sky130_fd_sc_hd__a31o_2 _38321_ (.A1(_10671_),
    .A2(_10672_),
    .A3(_10673_),
    .B1(_10735_),
    .X(_10736_));
 sky130_fd_sc_hd__a21oi_4 _38322_ (.A1(_10671_),
    .A2(_10672_),
    .B1(_10673_),
    .Y(_10737_));
 sky130_fd_sc_hd__o211a_1 _38323_ (.A1(_10736_),
    .A2(_10737_),
    .B1(_10732_),
    .C1(_10729_),
    .X(_10738_));
 sky130_fd_sc_hd__nor2_1 _38324_ (.A(_09172_),
    .B(_09170_),
    .Y(_10739_));
 sky130_fd_sc_hd__a21oi_1 _38325_ (.A1(_09170_),
    .A2(_09171_),
    .B1(_09174_),
    .Y(_10740_));
 sky130_fd_sc_hd__nor2_1 _38326_ (.A(_10739_),
    .B(_10740_),
    .Y(_10741_));
 sky130_fd_sc_hd__and2b_1 _38327_ (.A_N(_09413_),
    .B(_09422_),
    .X(_10742_));
 sky130_fd_sc_hd__and3b_1 _38328_ (.A_N(_09423_),
    .B(_09411_),
    .C(_09410_),
    .X(_10743_));
 sky130_fd_sc_hd__buf_1 _38329_ (.A(_09399_),
    .X(_10744_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38330_ (.A(_10744_),
    .X(_10746_));
 sky130_fd_sc_hd__nor2_2 _38331_ (.A(_04945_),
    .B(_06148_),
    .Y(_10747_));
 sky130_fd_sc_hd__and2_1 _38332_ (.A(_06148_),
    .B(_04945_),
    .X(_10748_));
 sky130_fd_sc_hd__nor2_1 _38333_ (.A(_10747_),
    .B(_10748_),
    .Y(_10749_));
 sky130_fd_sc_hd__xnor2_1 _38334_ (.A(_10746_),
    .B(_10749_),
    .Y(_10750_));
 sky130_fd_sc_hd__and2b_1 _38335_ (.A_N(_03464_),
    .B(_10744_),
    .X(_10751_));
 sky130_fd_sc_hd__o21ai_1 _38336_ (.A1(_04927_),
    .A2(_10744_),
    .B1(_09406_),
    .Y(_10752_));
 sky130_fd_sc_hd__a21oi_1 _38337_ (.A1(_04933_),
    .A2(_10744_),
    .B1(_10752_),
    .Y(_10753_));
 sky130_fd_sc_hd__a21o_1 _38338_ (.A1(_04933_),
    .A2(_10751_),
    .B1(_10753_),
    .X(_10754_));
 sky130_fd_sc_hd__xnor2_1 _38339_ (.A(_10750_),
    .B(_10754_),
    .Y(_10755_));
 sky130_fd_sc_hd__or2_1 _38340_ (.A(_09414_),
    .B(_09421_),
    .X(_10757_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38341_ (.A(_07947_),
    .X(_10758_));
 sky130_fd_sc_hd__nand3_2 _38342_ (.A(_09358_),
    .B(_09356_),
    .C(_09357_),
    .Y(_10759_));
 sky130_fd_sc_hd__o21a_1 _38343_ (.A1(_06097_),
    .A2(_07947_),
    .B1(_08010_),
    .X(_10760_));
 sky130_fd_sc_hd__o221ai_4 _38344_ (.A1(_04980_),
    .A2(_07947_),
    .B1(_07940_),
    .B2(_09359_),
    .C1(_10759_),
    .Y(_10761_));
 sky130_fd_sc_hd__o311a_1 _38345_ (.A1(_04980_),
    .A2(_10758_),
    .A3(_10759_),
    .B1(_10760_),
    .C1(_10761_),
    .X(_10762_));
 sky130_fd_sc_hd__or3_1 _38346_ (.A(_04980_),
    .B(_07947_),
    .C(_10759_),
    .X(_10763_));
 sky130_fd_sc_hd__a21oi_2 _38347_ (.A1(_10761_),
    .A2(_10763_),
    .B1(_10760_),
    .Y(_10764_));
 sky130_fd_sc_hd__a211oi_2 _38348_ (.A1(_09420_),
    .A2(_10757_),
    .B1(_10762_),
    .C1(_10764_),
    .Y(_10765_));
 sky130_fd_sc_hd__o221a_1 _38349_ (.A1(_09414_),
    .A2(_09421_),
    .B1(_10762_),
    .B2(_10764_),
    .C1(_09420_),
    .X(_10766_));
 sky130_fd_sc_hd__nor2_1 _38350_ (.A(_10765_),
    .B(_10766_),
    .Y(_10768_));
 sky130_fd_sc_hd__xnor2_1 _38351_ (.A(_10755_),
    .B(_10768_),
    .Y(_10769_));
 sky130_fd_sc_hd__o21a_1 _38352_ (.A1(_10742_),
    .A2(_10743_),
    .B1(_10769_),
    .X(_10770_));
 sky130_fd_sc_hd__o221a_1 _38353_ (.A1(_07998_),
    .A2(_07999_),
    .B1(_09381_),
    .B2(_09383_),
    .C1(_06157_),
    .X(_10771_));
 sky130_fd_sc_hd__and3_1 _38354_ (.A(_01865_),
    .B(_04941_),
    .C(_06125_),
    .X(_10772_));
 sky130_fd_sc_hd__buf_1 _38355_ (.A(_06148_),
    .X(_10773_));
 sky130_fd_sc_hd__a2111oi_1 _38356_ (.A1(_10744_),
    .A2(_09402_),
    .B1(_10772_),
    .C1(_10773_),
    .D1(_09400_),
    .Y(_10774_));
 sky130_fd_sc_hd__o22a_1 _38357_ (.A1(_10772_),
    .A2(_06148_),
    .B1(_09400_),
    .B2(_09405_),
    .X(_10775_));
 sky130_fd_sc_hd__o211a_1 _38358_ (.A1(net265),
    .A2(_10775_),
    .B1(_09408_),
    .C1(_09410_),
    .X(_10776_));
 sky130_fd_sc_hd__a211oi_1 _38359_ (.A1(_09408_),
    .A2(_09410_),
    .B1(net264),
    .C1(_10775_),
    .Y(_10777_));
 sky130_fd_sc_hd__a2111o_1 _38360_ (.A1(_09386_),
    .A2(_09385_),
    .B1(_10771_),
    .C1(_10776_),
    .D1(_10777_),
    .X(_10779_));
 sky130_fd_sc_hd__a21oi_1 _38361_ (.A1(_09385_),
    .A2(_09386_),
    .B1(_10771_),
    .Y(_10780_));
 sky130_fd_sc_hd__o21bai_1 _38362_ (.A1(_10777_),
    .A2(_10776_),
    .B1_N(_10780_),
    .Y(_10781_));
 sky130_fd_sc_hd__nand2_1 _38363_ (.A(_10779_),
    .B(_10781_),
    .Y(_10782_));
 sky130_fd_sc_hd__or3_1 _38364_ (.A(_10742_),
    .B(_10743_),
    .C(_10769_),
    .X(_10783_));
 sky130_fd_sc_hd__inv_2 _38365_ (.A(_10783_),
    .Y(_10784_));
 sky130_fd_sc_hd__or3_1 _38366_ (.A(_10770_),
    .B(_10782_),
    .C(_10784_),
    .X(_10785_));
 sky130_fd_sc_hd__o21ai_1 _38367_ (.A1(_10784_),
    .A2(_10770_),
    .B1(_10782_),
    .Y(_10786_));
 sky130_fd_sc_hd__and2_1 _38368_ (.A(_10785_),
    .B(_10786_),
    .X(_10787_));
 sky130_fd_sc_hd__a21o_1 _38369_ (.A1(_09376_),
    .A2(_09347_),
    .B1(_09374_),
    .X(_10788_));
 sky130_fd_sc_hd__a21bo_1 _38370_ (.A1(_09346_),
    .A2(_09367_),
    .B1_N(_09366_),
    .X(_10790_));
 sky130_fd_sc_hd__o211ai_2 _38371_ (.A1(_09120_),
    .A2(_07676_),
    .B1(_09134_),
    .C1(_07682_),
    .Y(_10791_));
 sky130_fd_sc_hd__a21o_1 _38372_ (.A1(_09150_),
    .A2(_10791_),
    .B1(_09137_),
    .X(_10792_));
 sky130_fd_sc_hd__o21a_1 _38373_ (.A1(_01744_),
    .A2(_03334_),
    .B1(_25296_),
    .X(_10793_));
 sky130_fd_sc_hd__or2_1 _38374_ (.A(_04973_),
    .B(_06091_),
    .X(_10794_));
 sky130_fd_sc_hd__nand2_1 _38375_ (.A(_09355_),
    .B(_24091_),
    .Y(_10795_));
 sky130_fd_sc_hd__o211a_2 _38376_ (.A1(_09352_),
    .A2(_10793_),
    .B1(_10794_),
    .C1(_10795_),
    .X(_10796_));
 sky130_fd_sc_hd__buf_1 _38377_ (.A(_09355_),
    .X(_10797_));
 sky130_fd_sc_hd__a221oi_2 _38378_ (.A1(_03341_),
    .A2(_03338_),
    .B1(_10794_),
    .B2(_10795_),
    .C1(_10793_),
    .Y(_10798_));
 sky130_fd_sc_hd__nor4_1 _38379_ (.A(_04971_),
    .B(_10796_),
    .C(_10797_),
    .D(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__o22a_1 _38380_ (.A1(_10797_),
    .A2(_04971_),
    .B1(_10796_),
    .B2(_10798_),
    .X(_10801_));
 sky130_fd_sc_hd__buf_1 _38381_ (.A(_03334_),
    .X(_10802_));
 sky130_fd_sc_hd__and2_1 _38382_ (.A(_10802_),
    .B(_06432_),
    .X(_10803_));
 sky130_fd_sc_hd__nor2_1 _38383_ (.A(\delay_line[7][13] ),
    .B(\delay_line[7][14] ),
    .Y(_10804_));
 sky130_fd_sc_hd__o21ba_1 _38384_ (.A1(_10803_),
    .A2(_10804_),
    .B1_N(_03341_),
    .X(_10805_));
 sky130_fd_sc_hd__nand2_2 _38385_ (.A(\delay_line[7][13] ),
    .B(_04659_),
    .Y(_10806_));
 sky130_fd_sc_hd__nand3b_2 _38386_ (.A_N(_10804_),
    .B(_01744_),
    .C(_10806_),
    .Y(_10807_));
 sky130_fd_sc_hd__inv_2 _38387_ (.A(_10807_),
    .Y(_10808_));
 sky130_fd_sc_hd__o22ai_1 _38388_ (.A1(_10799_),
    .A2(_10801_),
    .B1(_10805_),
    .B2(_10808_),
    .Y(_10809_));
 sky130_fd_sc_hd__or4_2 _38389_ (.A(_10799_),
    .B(_10801_),
    .C(_10805_),
    .D(_10808_),
    .X(_10810_));
 sky130_fd_sc_hd__a21boi_1 _38390_ (.A1(_09145_),
    .A2(_09149_),
    .B1_N(_09146_),
    .Y(_10812_));
 sky130_fd_sc_hd__a21boi_1 _38391_ (.A1(_10809_),
    .A2(_10810_),
    .B1_N(_10812_),
    .Y(_10813_));
 sky130_fd_sc_hd__and3b_1 _38392_ (.A_N(_10812_),
    .B(_10809_),
    .C(_10810_),
    .X(_10814_));
 sky130_fd_sc_hd__o21bai_1 _38393_ (.A1(_10813_),
    .A2(_10814_),
    .B1_N(_09364_),
    .Y(_10815_));
 sky130_fd_sc_hd__or3b_1 _38394_ (.A(_10813_),
    .B(_10814_),
    .C_N(_09364_),
    .X(_10816_));
 sky130_fd_sc_hd__nand3_2 _38395_ (.A(_10792_),
    .B(_10815_),
    .C(_10816_),
    .Y(_10817_));
 sky130_fd_sc_hd__a221o_1 _38396_ (.A1(_09150_),
    .A2(_10791_),
    .B1(_10816_),
    .B2(_10815_),
    .C1(_09137_),
    .X(_10818_));
 sky130_fd_sc_hd__and3_1 _38397_ (.A(_10790_),
    .B(_10817_),
    .C(_10818_),
    .X(_10819_));
 sky130_fd_sc_hd__a21oi_1 _38398_ (.A1(_10817_),
    .A2(_10818_),
    .B1(_10790_),
    .Y(_10820_));
 sky130_fd_sc_hd__a211o_1 _38399_ (.A1(_09373_),
    .A2(_10788_),
    .B1(_10819_),
    .C1(_10820_),
    .X(_10821_));
 sky130_fd_sc_hd__o221ai_2 _38400_ (.A1(_09348_),
    .A2(_09370_),
    .B1(_10820_),
    .B2(_10819_),
    .C1(_10788_),
    .Y(_10823_));
 sky130_fd_sc_hd__nand2_2 _38401_ (.A(_10821_),
    .B(_10823_),
    .Y(_10824_));
 sky130_fd_sc_hd__xnor2_2 _38402_ (.A(_10787_),
    .B(_10824_),
    .Y(_10825_));
 sky130_fd_sc_hd__or2_1 _38403_ (.A(_10741_),
    .B(_10825_),
    .X(_10826_));
 sky130_fd_sc_hd__nand2_1 _38404_ (.A(_10825_),
    .B(_10741_),
    .Y(_10827_));
 sky130_fd_sc_hd__a221o_1 _38405_ (.A1(_09427_),
    .A2(_09379_),
    .B1(_10826_),
    .B2(_10827_),
    .C1(_09378_),
    .X(_10828_));
 sky130_fd_sc_hd__a21oi_1 _38406_ (.A1(_09427_),
    .A2(_09379_),
    .B1(_09378_),
    .Y(_10829_));
 sky130_fd_sc_hd__nand3b_2 _38407_ (.A_N(_10829_),
    .B(_10826_),
    .C(_10827_),
    .Y(_10830_));
 sky130_fd_sc_hd__nand2_1 _38408_ (.A(_10828_),
    .B(_10830_),
    .Y(_10831_));
 sky130_fd_sc_hd__clkbuf_2 _38409_ (.A(_10831_),
    .X(_10832_));
 sky130_fd_sc_hd__o21ai_2 _38410_ (.A1(_10733_),
    .A2(_10738_),
    .B1(_10832_),
    .Y(_10834_));
 sky130_fd_sc_hd__a21o_1 _38411_ (.A1(_10729_),
    .A2(_10731_),
    .B1(_10732_),
    .X(_10835_));
 sky130_fd_sc_hd__o211ai_2 _38412_ (.A1(_10737_),
    .A2(_10736_),
    .B1(_10729_),
    .C1(_10732_),
    .Y(_10836_));
 sky130_fd_sc_hd__nand3b_2 _38413_ (.A_N(_10832_),
    .B(_10835_),
    .C(_10836_),
    .Y(_10837_));
 sky130_fd_sc_hd__nand3_1 _38414_ (.A(_10494_),
    .B(_10834_),
    .C(_10837_),
    .Y(_10838_));
 sky130_fd_sc_hd__o21bai_1 _38415_ (.A1(_10733_),
    .A2(_10738_),
    .B1_N(_10831_),
    .Y(_10839_));
 sky130_fd_sc_hd__nand3_1 _38416_ (.A(_10832_),
    .B(_10835_),
    .C(_10836_),
    .Y(_10840_));
 sky130_fd_sc_hd__inv_2 _38417_ (.A(_09337_),
    .Y(_10841_));
 sky130_fd_sc_hd__a21oi_1 _38418_ (.A1(_09439_),
    .A2(_09343_),
    .B1(_10841_),
    .Y(_10842_));
 sky130_fd_sc_hd__nand3_1 _38419_ (.A(_10839_),
    .B(_10840_),
    .C(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__o22ai_2 _38420_ (.A1(_08067_),
    .A2(_08071_),
    .B1(_09469_),
    .B2(_09467_),
    .Y(_10845_));
 sky130_fd_sc_hd__or2_1 _38421_ (.A(_09454_),
    .B(_09466_),
    .X(_10846_));
 sky130_fd_sc_hd__o21a_1 _38422_ (.A1(_09464_),
    .A2(_09465_),
    .B1(_10846_),
    .X(_10847_));
 sky130_fd_sc_hd__a211oi_1 _38423_ (.A1(_08055_),
    .A2(_09461_),
    .B1(_09458_),
    .C1(_09460_),
    .Y(_10848_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38424_ (.A(_06125_),
    .X(_10849_));
 sky130_fd_sc_hd__o31a_1 _38425_ (.A1(_08047_),
    .A2(_04908_),
    .A3(_08046_),
    .B1(_06511_),
    .X(_10850_));
 sky130_fd_sc_hd__o21ai_1 _38426_ (.A1(net446),
    .A2(_06510_),
    .B1(_06125_),
    .Y(_10851_));
 sky130_fd_sc_hd__or3_1 _38427_ (.A(\delay_line[1][14] ),
    .B(_06125_),
    .C(_06510_),
    .X(_10852_));
 sky130_fd_sc_hd__a21bo_1 _38428_ (.A1(_10851_),
    .A2(_10852_),
    .B1_N(_10850_),
    .X(_10853_));
 sky130_fd_sc_hd__o21a_1 _38429_ (.A1(_10849_),
    .A2(_10850_),
    .B1(_10853_),
    .X(_10854_));
 sky130_fd_sc_hd__or3_1 _38430_ (.A(_09389_),
    .B(_09396_),
    .C(_10854_),
    .X(_10856_));
 sky130_fd_sc_hd__o21ai_1 _38431_ (.A1(_09389_),
    .A2(_09396_),
    .B1(_10854_),
    .Y(_10857_));
 sky130_fd_sc_hd__o211a_1 _38432_ (.A1(_09460_),
    .A2(_10848_),
    .B1(_10856_),
    .C1(_10857_),
    .X(_10858_));
 sky130_fd_sc_hd__a211oi_1 _38433_ (.A1(_10856_),
    .A2(_10857_),
    .B1(_09460_),
    .C1(_10848_),
    .Y(_10859_));
 sky130_fd_sc_hd__nor2_1 _38434_ (.A(_10858_),
    .B(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__or2_1 _38435_ (.A(_09424_),
    .B(_09398_),
    .X(_10861_));
 sky130_fd_sc_hd__o21ai_1 _38436_ (.A1(_09397_),
    .A2(_09425_),
    .B1(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__xor2_1 _38437_ (.A(_10860_),
    .B(_10862_),
    .X(_10863_));
 sky130_fd_sc_hd__xor2_2 _38438_ (.A(_10847_),
    .B(_10863_),
    .X(_10864_));
 sky130_fd_sc_hd__a21oi_2 _38439_ (.A1(_09471_),
    .A2(_10845_),
    .B1(_10864_),
    .Y(_10865_));
 sky130_fd_sc_hd__and3_1 _38440_ (.A(_10864_),
    .B(_10845_),
    .C(_09471_),
    .X(_10867_));
 sky130_fd_sc_hd__or2_1 _38441_ (.A(_10865_),
    .B(_10867_),
    .X(_10868_));
 sky130_fd_sc_hd__a21o_1 _38442_ (.A1(_09431_),
    .A2(_09436_),
    .B1(_10868_),
    .X(_10869_));
 sky130_fd_sc_hd__or2_1 _38443_ (.A(_09453_),
    .B(_09475_),
    .X(_10870_));
 sky130_fd_sc_hd__o211ai_2 _38444_ (.A1(_09434_),
    .A2(_09432_),
    .B1(_09431_),
    .C1(_10868_),
    .Y(_10871_));
 sky130_fd_sc_hd__inv_2 _38445_ (.A(_10871_),
    .Y(_10872_));
 sky130_fd_sc_hd__nor2_1 _38446_ (.A(_10870_),
    .B(_10872_),
    .Y(_10873_));
 sky130_fd_sc_hd__nand2_1 _38447_ (.A(_10869_),
    .B(_10871_),
    .Y(_10874_));
 sky130_fd_sc_hd__a22oi_1 _38448_ (.A1(_10869_),
    .A2(_10873_),
    .B1(_10874_),
    .B2(_10870_),
    .Y(_10875_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38449_ (.A(_10875_),
    .X(_10876_));
 sky130_fd_sc_hd__a21bo_1 _38450_ (.A1(_10838_),
    .A2(_10843_),
    .B1_N(_10876_),
    .X(_10878_));
 sky130_fd_sc_hd__nand2_1 _38451_ (.A(_09344_),
    .B(_09439_),
    .Y(_10879_));
 sky130_fd_sc_hd__o21ai_1 _38452_ (.A1(_10879_),
    .A2(_10841_),
    .B1(_09449_),
    .Y(_10880_));
 sky130_fd_sc_hd__a21oi_1 _38453_ (.A1(_07928_),
    .A2(_08031_),
    .B1(_09445_),
    .Y(_10881_));
 sky130_fd_sc_hd__nand2_1 _38454_ (.A(_10880_),
    .B(_10881_),
    .Y(_10882_));
 sky130_fd_sc_hd__o221a_1 _38455_ (.A1(_10879_),
    .A2(_10841_),
    .B1(_09446_),
    .B2(_09445_),
    .C1(_09449_),
    .X(_10883_));
 sky130_fd_sc_hd__a21oi_1 _38456_ (.A1(_10882_),
    .A2(_09483_),
    .B1(_10883_),
    .Y(_10884_));
 sky130_fd_sc_hd__clkbuf_2 _38457_ (.A(_10843_),
    .X(_10885_));
 sky130_fd_sc_hd__nand3b_1 _38458_ (.A_N(_10875_),
    .B(_10838_),
    .C(_10885_),
    .Y(_10886_));
 sky130_fd_sc_hd__nand3_1 _38459_ (.A(_10878_),
    .B(_10884_),
    .C(_10886_),
    .Y(_10887_));
 sky130_fd_sc_hd__clkbuf_2 _38460_ (.A(_10887_),
    .X(_10889_));
 sky130_fd_sc_hd__a21oi_1 _38461_ (.A1(_10881_),
    .A2(_10880_),
    .B1(_09487_),
    .Y(_10890_));
 sky130_fd_sc_hd__nand3_1 _38462_ (.A(_10838_),
    .B(_10885_),
    .C(_10876_),
    .Y(_10891_));
 sky130_fd_sc_hd__a21o_1 _38463_ (.A1(_10838_),
    .A2(_10885_),
    .B1(_10876_),
    .X(_10892_));
 sky130_fd_sc_hd__o211ai_4 _38464_ (.A1(_10883_),
    .A2(_10890_),
    .B1(_10891_),
    .C1(_10892_),
    .Y(_10893_));
 sky130_fd_sc_hd__or2_1 _38465_ (.A(_09477_),
    .B(net89),
    .X(_10894_));
 sky130_fd_sc_hd__a21oi_1 _38466_ (.A1(_10889_),
    .A2(_10893_),
    .B1(_10894_),
    .Y(_10895_));
 sky130_fd_sc_hd__clkbuf_2 _38467_ (.A(_10893_),
    .X(_10896_));
 sky130_fd_sc_hd__a21oi_2 _38468_ (.A1(_09494_),
    .A2(_09497_),
    .B1(_09500_),
    .Y(_10897_));
 sky130_fd_sc_hd__a31o_2 _38469_ (.A1(_10894_),
    .A2(_10889_),
    .A3(_10896_),
    .B1(_10897_),
    .X(_10898_));
 sky130_fd_sc_hd__o211a_1 _38470_ (.A1(_09477_),
    .A2(net89),
    .B1(_10887_),
    .C1(_10893_),
    .X(_10900_));
 sky130_fd_sc_hd__o21ai_1 _38471_ (.A1(_10895_),
    .A2(_10900_),
    .B1(_10897_),
    .Y(_10901_));
 sky130_fd_sc_hd__clkbuf_2 _38472_ (.A(_10901_),
    .X(_10902_));
 sky130_fd_sc_hd__o21a_1 _38473_ (.A1(_10895_),
    .A2(_10898_),
    .B1(_10902_),
    .X(_10903_));
 sky130_fd_sc_hd__o21ai_1 _38474_ (.A1(_10490_),
    .A2(_10493_),
    .B1(_10903_),
    .Y(_10904_));
 sky130_fd_sc_hd__buf_2 _38475_ (.A(_10895_),
    .X(_10905_));
 sky130_fd_sc_hd__o21ai_2 _38476_ (.A1(_10905_),
    .A2(_10898_),
    .B1(_10902_),
    .Y(_10906_));
 sky130_fd_sc_hd__a21o_1 _38477_ (.A1(_09523_),
    .A2(_09508_),
    .B1(_10489_),
    .X(_10907_));
 sky130_fd_sc_hd__and4_2 _38478_ (.A(_08109_),
    .B(_08114_),
    .C(_09505_),
    .D(_09508_),
    .X(_10908_));
 sky130_fd_sc_hd__nand2_1 _38479_ (.A(_08127_),
    .B(_10908_),
    .Y(_10909_));
 sky130_fd_sc_hd__nand3_1 _38480_ (.A(_10906_),
    .B(_10907_),
    .C(_10909_),
    .Y(_10911_));
 sky130_fd_sc_hd__nand3_1 _38481_ (.A(_10488_),
    .B(_10904_),
    .C(_10911_),
    .Y(_10912_));
 sky130_fd_sc_hd__o21ai_1 _38482_ (.A1(_10490_),
    .A2(_10493_),
    .B1(_10906_),
    .Y(_10913_));
 sky130_fd_sc_hd__o2111ai_2 _38483_ (.A1(_10898_),
    .A2(_10905_),
    .B1(_10902_),
    .C1(_10907_),
    .D1(_10909_),
    .Y(_10914_));
 sky130_fd_sc_hd__inv_2 _38484_ (.A(_10488_),
    .Y(_10915_));
 sky130_fd_sc_hd__nand3_2 _38485_ (.A(_10913_),
    .B(_10914_),
    .C(_10915_),
    .Y(_10916_));
 sky130_fd_sc_hd__a21o_1 _38486_ (.A1(_10912_),
    .A2(_10916_),
    .B1(_09526_),
    .X(_10917_));
 sky130_fd_sc_hd__a21oi_1 _38487_ (.A1(_10907_),
    .A2(_10909_),
    .B1(_10906_),
    .Y(_10918_));
 sky130_fd_sc_hd__nand2_1 _38488_ (.A(_10488_),
    .B(_10911_),
    .Y(_10919_));
 sky130_fd_sc_hd__o211ai_2 _38489_ (.A1(_10918_),
    .A2(_10919_),
    .B1(_10916_),
    .C1(_09526_),
    .Y(_10920_));
 sky130_fd_sc_hd__o21bai_1 _38490_ (.A1(_09710_),
    .A2(_09709_),
    .B1_N(_09737_),
    .Y(_10922_));
 sky130_fd_sc_hd__inv_2 _38491_ (.A(_10922_),
    .Y(_10923_));
 sky130_fd_sc_hd__a31o_1 _38492_ (.A1(_08267_),
    .A2(_08270_),
    .A3(_09709_),
    .B1(_10923_),
    .X(_10924_));
 sky130_fd_sc_hd__inv_2 _38493_ (.A(_10924_),
    .Y(_10925_));
 sky130_fd_sc_hd__nand3_2 _38494_ (.A(_10917_),
    .B(_10920_),
    .C(_10925_),
    .Y(_10926_));
 sky130_fd_sc_hd__inv_2 _38495_ (.A(_09711_),
    .Y(_10927_));
 sky130_fd_sc_hd__a21oi_2 _38496_ (.A1(_10912_),
    .A2(_10916_),
    .B1(_09526_),
    .Y(_10928_));
 sky130_fd_sc_hd__o211a_1 _38497_ (.A1(_10918_),
    .A2(_10919_),
    .B1(_10916_),
    .C1(_09521_),
    .X(_10929_));
 sky130_fd_sc_hd__o22ai_4 _38498_ (.A1(_10927_),
    .A2(_10923_),
    .B1(_10928_),
    .B2(_10929_),
    .Y(_10930_));
 sky130_fd_sc_hd__a22o_2 _38499_ (.A1(_10486_),
    .A2(_09528_),
    .B1(_10926_),
    .B2(_10930_),
    .X(_10931_));
 sky130_fd_sc_hd__inv_2 _38500_ (.A(\delay_line[23][15] ),
    .Y(_10933_));
 sky130_fd_sc_hd__clkbuf_2 _38501_ (.A(_10933_),
    .X(_10934_));
 sky130_fd_sc_hd__buf_2 _38502_ (.A(_10934_),
    .X(_10935_));
 sky130_fd_sc_hd__o2111ai_4 _38503_ (.A1(_10935_),
    .A2(_09515_),
    .B1(_10486_),
    .C1(_10926_),
    .D1(_10930_),
    .Y(_10936_));
 sky130_fd_sc_hd__nand3_1 _38504_ (.A(_10485_),
    .B(_10931_),
    .C(_10936_),
    .Y(_10937_));
 sky130_fd_sc_hd__and3_2 _38505_ (.A(_10917_),
    .B(_10920_),
    .C(_10925_),
    .X(_10938_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38506_ (.A(_09521_),
    .X(_10939_));
 sky130_fd_sc_hd__a2bb2o_1 _38507_ (.A1_N(_09524_),
    .A2_N(_09519_),
    .B1(_10939_),
    .B2(_09527_),
    .X(_10940_));
 sky130_fd_sc_hd__nand2_2 _38508_ (.A(_10940_),
    .B(_10930_),
    .Y(_10941_));
 sky130_fd_sc_hd__a21oi_2 _38509_ (.A1(_09533_),
    .A2(_09529_),
    .B1(_09538_),
    .Y(_10942_));
 sky130_fd_sc_hd__a21o_1 _38510_ (.A1(_10926_),
    .A2(_10930_),
    .B1(_10940_),
    .X(_10944_));
 sky130_fd_sc_hd__o221ai_4 _38511_ (.A1(_10938_),
    .A2(_10941_),
    .B1(_09531_),
    .B2(_10942_),
    .C1(_10944_),
    .Y(_10945_));
 sky130_fd_sc_hd__o2bb2a_1 _38512_ (.A1_N(_08158_),
    .A2_N(_00437_),
    .B1(_24256_),
    .B2(_22750_),
    .X(_10946_));
 sky130_fd_sc_hd__nand2_1 _38513_ (.A(_08158_),
    .B(_00437_),
    .Y(_10947_));
 sky130_fd_sc_hd__nor2_1 _38514_ (.A(_06644_),
    .B(_10947_),
    .Y(_10948_));
 sky130_fd_sc_hd__o21ai_1 _38515_ (.A1(_03565_),
    .A2(_10933_),
    .B1(_08163_),
    .Y(_10949_));
 sky130_fd_sc_hd__or3_1 _38516_ (.A(_03564_),
    .B(_03066_),
    .C(_10933_),
    .X(_10950_));
 sky130_fd_sc_hd__and2_1 _38517_ (.A(_10949_),
    .B(_10950_),
    .X(_10951_));
 sky130_fd_sc_hd__or3_2 _38518_ (.A(_10946_),
    .B(_10948_),
    .C(_10951_),
    .X(_10952_));
 sky130_fd_sc_hd__inv_2 _38519_ (.A(_10952_),
    .Y(_10953_));
 sky130_fd_sc_hd__o21a_2 _38520_ (.A1(_10946_),
    .A2(_10948_),
    .B1(_10951_),
    .X(_10955_));
 sky130_fd_sc_hd__nor2_1 _38521_ (.A(_10953_),
    .B(_10955_),
    .Y(_10956_));
 sky130_fd_sc_hd__a21bo_1 _38522_ (.A1(_10937_),
    .A2(_10945_),
    .B1_N(_10956_),
    .X(_10957_));
 sky130_fd_sc_hd__o21a_1 _38523_ (.A1(_09749_),
    .A2(_09746_),
    .B1(_09748_),
    .X(_10958_));
 sky130_fd_sc_hd__clkbuf_2 _38524_ (.A(_10937_),
    .X(_10959_));
 sky130_fd_sc_hd__clkbuf_2 _38525_ (.A(_10945_),
    .X(_10960_));
 sky130_fd_sc_hd__o211ai_1 _38526_ (.A1(_10953_),
    .A2(_10955_),
    .B1(_10959_),
    .C1(_10960_),
    .Y(_10961_));
 sky130_fd_sc_hd__nand3_1 _38527_ (.A(_10957_),
    .B(_10958_),
    .C(_10961_),
    .Y(_10962_));
 sky130_fd_sc_hd__inv_2 _38528_ (.A(_09748_),
    .Y(_10963_));
 sky130_fd_sc_hd__nand3_1 _38529_ (.A(_10959_),
    .B(_10960_),
    .C(_10956_),
    .Y(_10964_));
 sky130_fd_sc_hd__o2bb2ai_1 _38530_ (.A1_N(_10959_),
    .A2_N(_10960_),
    .B1(_10953_),
    .B2(_10955_),
    .Y(_10966_));
 sky130_fd_sc_hd__o211ai_2 _38531_ (.A1(_10963_),
    .A2(_09751_),
    .B1(_10964_),
    .C1(_10966_),
    .Y(_10967_));
 sky130_fd_sc_hd__a32o_1 _38532_ (.A1(_09552_),
    .A2(_09553_),
    .A3(_09554_),
    .B1(_09560_),
    .B2(_09549_),
    .X(_10968_));
 sky130_fd_sc_hd__a21oi_1 _38533_ (.A1(_10962_),
    .A2(_10967_),
    .B1(_10968_),
    .Y(_10969_));
 sky130_fd_sc_hd__o21bai_2 _38534_ (.A1(_10275_),
    .A2(_10276_),
    .B1_N(_10279_),
    .Y(_10970_));
 sky130_fd_sc_hd__a21oi_1 _38535_ (.A1(_10125_),
    .A2(_10274_),
    .B1(_10124_),
    .Y(_10971_));
 sky130_fd_sc_hd__o32ai_2 _38536_ (.A1(_09991_),
    .A2(_09993_),
    .A3(_09990_),
    .B1(_09995_),
    .B2(_09895_),
    .Y(_10972_));
 sky130_fd_sc_hd__clkbuf_2 _38537_ (.A(_22954_),
    .X(_10973_));
 sky130_fd_sc_hd__a211o_1 _38538_ (.A1(_07409_),
    .A2(_10973_),
    .B1(_22944_),
    .C1(_09819_),
    .X(_10974_));
 sky130_fd_sc_hd__nand2_1 _38539_ (.A(_09817_),
    .B(_09823_),
    .Y(_10975_));
 sky130_fd_sc_hd__o21ai_1 _38540_ (.A1(_10973_),
    .A2(_00653_),
    .B1(_04043_),
    .Y(_10977_));
 sky130_fd_sc_hd__or3_1 _38541_ (.A(_24661_),
    .B(_02588_),
    .C(_02589_),
    .X(_10978_));
 sky130_fd_sc_hd__buf_1 _38542_ (.A(_02588_),
    .X(_10979_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38543_ (.A(_24661_),
    .X(_10980_));
 sky130_fd_sc_hd__o21ai_1 _38544_ (.A1(_10979_),
    .A2(_02589_),
    .B1(_10980_),
    .Y(_10981_));
 sky130_fd_sc_hd__and3_1 _38545_ (.A(_10977_),
    .B(_10978_),
    .C(_10981_),
    .X(_10982_));
 sky130_fd_sc_hd__a21oi_1 _38546_ (.A1(_10978_),
    .A2(_10981_),
    .B1(_10977_),
    .Y(_10983_));
 sky130_fd_sc_hd__xor2_1 _38547_ (.A(_05698_),
    .B(_08735_),
    .X(_10984_));
 sky130_fd_sc_hd__nand3b_1 _38548_ (.A_N(_05698_),
    .B(_08733_),
    .C(_09799_),
    .Y(_10985_));
 sky130_fd_sc_hd__o21a_1 _38549_ (.A1(_09802_),
    .A2(_10984_),
    .B1(_10985_),
    .X(_10986_));
 sky130_fd_sc_hd__or3b_1 _38550_ (.A(_10982_),
    .B(_10983_),
    .C_N(_10986_),
    .X(_10988_));
 sky130_fd_sc_hd__o21bai_1 _38551_ (.A1(_10982_),
    .A2(_10983_),
    .B1_N(_10986_),
    .Y(_10989_));
 sky130_fd_sc_hd__a21bo_1 _38552_ (.A1(_09805_),
    .A2(_09810_),
    .B1_N(_09806_),
    .X(_10990_));
 sky130_fd_sc_hd__a21oi_1 _38553_ (.A1(_10988_),
    .A2(_10989_),
    .B1(_10990_),
    .Y(_10991_));
 sky130_fd_sc_hd__and3_1 _38554_ (.A(_10990_),
    .B(_10988_),
    .C(_10989_),
    .X(_10992_));
 sky130_fd_sc_hd__nor2_1 _38555_ (.A(_10991_),
    .B(_10992_),
    .Y(_10993_));
 sky130_fd_sc_hd__a21o_1 _38556_ (.A1(_22944_),
    .A2(_10980_),
    .B1(_09807_),
    .X(_10994_));
 sky130_fd_sc_hd__a21o_1 _38557_ (.A1(_04055_),
    .A2(_07423_),
    .B1(_07427_),
    .X(_10995_));
 sky130_fd_sc_hd__and3_1 _38558_ (.A(_10993_),
    .B(_10994_),
    .C(_10995_),
    .X(_10996_));
 sky130_fd_sc_hd__a21oi_1 _38559_ (.A1(_10994_),
    .A2(_10995_),
    .B1(_10993_),
    .Y(_10997_));
 sky130_fd_sc_hd__nor2_1 _38560_ (.A(_10996_),
    .B(_10997_),
    .Y(_10999_));
 sky130_fd_sc_hd__xnor2_1 _38561_ (.A(_10975_),
    .B(_10999_),
    .Y(_11000_));
 sky130_fd_sc_hd__xor2_1 _38562_ (.A(_10974_),
    .B(_11000_),
    .X(_11001_));
 sky130_fd_sc_hd__a311o_2 _38563_ (.A1(_08719_),
    .A2(_09827_),
    .A3(_09828_),
    .B1(_09826_),
    .C1(_11001_),
    .X(_11002_));
 sky130_fd_sc_hd__o21a_1 _38564_ (.A1(_09826_),
    .A2(_09829_),
    .B1(_11001_),
    .X(_11003_));
 sky130_fd_sc_hd__inv_2 _38565_ (.A(_11003_),
    .Y(_11004_));
 sky130_fd_sc_hd__a2bb2o_1 _38566_ (.A1_N(_09834_),
    .A2_N(_09840_),
    .B1(_11002_),
    .B2(_11004_),
    .X(_11005_));
 sky130_fd_sc_hd__or4bb_1 _38567_ (.A(_09834_),
    .B(_09840_),
    .C_N(_11002_),
    .D_N(_11004_),
    .X(_11006_));
 sky130_fd_sc_hd__or4b_1 _38568_ (.A(_07375_),
    .B(_07376_),
    .C(_09753_),
    .D_N(_09784_),
    .X(_11007_));
 sky130_fd_sc_hd__or3b_1 _38569_ (.A(_07376_),
    .B(_09755_),
    .C_N(_09753_),
    .X(_11008_));
 sky130_fd_sc_hd__o21ai_1 _38570_ (.A1(_09757_),
    .A2(_09777_),
    .B1(_09776_),
    .Y(_11010_));
 sky130_fd_sc_hd__clkbuf_2 _38571_ (.A(_09768_),
    .X(_11011_));
 sky130_fd_sc_hd__inv_2 _38572_ (.A(_11011_),
    .Y(_11012_));
 sky130_fd_sc_hd__clkbuf_2 _38573_ (.A(_09766_),
    .X(_11013_));
 sky130_fd_sc_hd__a21oi_1 _38574_ (.A1(_11012_),
    .A2(_08687_),
    .B1(_11013_),
    .Y(_11014_));
 sky130_fd_sc_hd__o21ai_1 _38575_ (.A1(_09764_),
    .A2(_08694_),
    .B1(_09771_),
    .Y(_11015_));
 sky130_fd_sc_hd__clkbuf_2 _38576_ (.A(_05646_),
    .X(_11016_));
 sky130_fd_sc_hd__a21oi_2 _38577_ (.A1(_09766_),
    .A2(_09768_),
    .B1(_02638_),
    .Y(_11017_));
 sky130_fd_sc_hd__and3_1 _38578_ (.A(_09766_),
    .B(_02638_),
    .C(_09768_),
    .X(_11018_));
 sky130_fd_sc_hd__nor2_1 _38579_ (.A(_05646_),
    .B(_09758_),
    .Y(_11019_));
 sky130_fd_sc_hd__and2_1 _38580_ (.A(_05646_),
    .B(net372),
    .X(_11021_));
 sky130_fd_sc_hd__a2bb2o_1 _38581_ (.A1_N(_11019_),
    .A2_N(_11021_),
    .B1(_09764_),
    .B2(_09758_),
    .X(_11022_));
 sky130_fd_sc_hd__o221ai_4 _38582_ (.A1(_11016_),
    .A2(_09759_),
    .B1(_11017_),
    .B2(_11018_),
    .C1(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__buf_1 _38583_ (.A(_09760_),
    .X(_11024_));
 sky130_fd_sc_hd__or3_1 _38584_ (.A(_11016_),
    .B(_09761_),
    .C(_11024_),
    .X(_11025_));
 sky130_fd_sc_hd__a211o_1 _38585_ (.A1(_11022_),
    .A2(_11025_),
    .B1(_11017_),
    .C1(_11018_),
    .X(_11026_));
 sky130_fd_sc_hd__and4_2 _38586_ (.A(_09763_),
    .B(_11015_),
    .C(_11023_),
    .D(_11026_),
    .X(_11027_));
 sky130_fd_sc_hd__a22o_1 _38587_ (.A1(_09763_),
    .A2(_11015_),
    .B1(_11023_),
    .B2(_11026_),
    .X(_11028_));
 sky130_fd_sc_hd__and2b_1 _38588_ (.A_N(_11027_),
    .B(_11028_),
    .X(_11029_));
 sky130_fd_sc_hd__xor2_1 _38589_ (.A(_11014_),
    .B(_11029_),
    .X(_11030_));
 sky130_fd_sc_hd__nor2_1 _38590_ (.A(_11010_),
    .B(_11030_),
    .Y(_11032_));
 sky130_fd_sc_hd__nand2_1 _38591_ (.A(_11030_),
    .B(_11010_),
    .Y(_11033_));
 sky130_fd_sc_hd__and2b_1 _38592_ (.A_N(_11032_),
    .B(_11033_),
    .X(_11034_));
 sky130_fd_sc_hd__xnor2_1 _38593_ (.A(_11008_),
    .B(_11034_),
    .Y(_11035_));
 sky130_fd_sc_hd__a21bo_1 _38594_ (.A1(_09783_),
    .A2(_11007_),
    .B1_N(_11035_),
    .X(_11036_));
 sky130_fd_sc_hd__a211o_1 _38595_ (.A1(_09779_),
    .A2(_09781_),
    .B1(_09788_),
    .C1(_11035_),
    .X(_11037_));
 sky130_fd_sc_hd__nand2_1 _38596_ (.A(_11036_),
    .B(_11037_),
    .Y(_11038_));
 sky130_fd_sc_hd__o221a_1 _38597_ (.A1(_09785_),
    .A2(_09787_),
    .B1(_09791_),
    .B2(_09793_),
    .C1(_11038_),
    .X(_11039_));
 sky130_fd_sc_hd__o22ai_1 _38598_ (.A1(_09785_),
    .A2(_09787_),
    .B1(_09791_),
    .B2(_09793_),
    .Y(_11040_));
 sky130_fd_sc_hd__inv_2 _38599_ (.A(_11038_),
    .Y(_11041_));
 sky130_fd_sc_hd__nand2_1 _38600_ (.A(_11040_),
    .B(_11041_),
    .Y(_11043_));
 sky130_fd_sc_hd__or2b_1 _38601_ (.A(_11039_),
    .B_N(_11043_),
    .X(_11044_));
 sky130_fd_sc_hd__a21o_1 _38602_ (.A1(_11005_),
    .A2(_11006_),
    .B1(_11044_),
    .X(_11045_));
 sky130_fd_sc_hd__nand3_1 _38603_ (.A(_11044_),
    .B(_11005_),
    .C(_11006_),
    .Y(_11046_));
 sky130_fd_sc_hd__and2_1 _38604_ (.A(_11045_),
    .B(_11046_),
    .X(_11047_));
 sky130_fd_sc_hd__buf_1 _38605_ (.A(_04094_),
    .X(_11048_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38606_ (.A(_08652_),
    .X(_11049_));
 sky130_fd_sc_hd__buf_1 _38607_ (.A(_09845_),
    .X(_11050_));
 sky130_fd_sc_hd__and4b_2 _38608_ (.A_N(_11048_),
    .B(_11049_),
    .C(_11050_),
    .D(_09846_),
    .X(_11051_));
 sky130_fd_sc_hd__nand2_1 _38609_ (.A(_11048_),
    .B(_11050_),
    .Y(_11052_));
 sky130_fd_sc_hd__or2_1 _38610_ (.A(_11048_),
    .B(_09845_),
    .X(_11054_));
 sky130_fd_sc_hd__a21oi_1 _38611_ (.A1(_11052_),
    .A2(_11054_),
    .B1(_09848_),
    .Y(_11055_));
 sky130_fd_sc_hd__a21o_1 _38612_ (.A1(_05609_),
    .A2(_09854_),
    .B1(_09853_),
    .X(_11056_));
 sky130_fd_sc_hd__buf_1 _38613_ (.A(_02540_),
    .X(_11057_));
 sky130_fd_sc_hd__buf_1 _38614_ (.A(_02541_),
    .X(_11058_));
 sky130_fd_sc_hd__buf_1 _38615_ (.A(_24635_),
    .X(_11059_));
 sky130_fd_sc_hd__or3b_1 _38616_ (.A(_11057_),
    .B(_11058_),
    .C_N(_11059_),
    .X(_11060_));
 sky130_fd_sc_hd__nor2_1 _38617_ (.A(_11057_),
    .B(_02541_),
    .Y(_11061_));
 sky130_fd_sc_hd__or2_1 _38618_ (.A(_11059_),
    .B(_11061_),
    .X(_11062_));
 sky130_fd_sc_hd__and3_1 _38619_ (.A(_11056_),
    .B(_11060_),
    .C(_11062_),
    .X(_11063_));
 sky130_fd_sc_hd__a21oi_1 _38620_ (.A1(_11060_),
    .A2(_11062_),
    .B1(_11056_),
    .Y(_11065_));
 sky130_fd_sc_hd__nor4_1 _38621_ (.A(_11051_),
    .B(_11055_),
    .C(_11063_),
    .D(_11065_),
    .Y(_11066_));
 sky130_fd_sc_hd__o22a_1 _38622_ (.A1(_11051_),
    .A2(_11055_),
    .B1(_11063_),
    .B2(_11065_),
    .X(_11067_));
 sky130_fd_sc_hd__a211oi_4 _38623_ (.A1(_09852_),
    .A2(_09859_),
    .B1(net222),
    .C1(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38624_ (.A(_11059_),
    .X(_11069_));
 sky130_fd_sc_hd__o22a_1 _38625_ (.A1(_09867_),
    .A2(_11069_),
    .B1(_00614_),
    .B2(_09853_),
    .X(_11070_));
 sky130_fd_sc_hd__or3_1 _38626_ (.A(_07340_),
    .B(_08645_),
    .C(_11070_),
    .X(_11071_));
 sky130_fd_sc_hd__o211ai_1 _38627_ (.A1(net222),
    .A2(_11067_),
    .B1(_09852_),
    .C1(_09859_),
    .Y(_11072_));
 sky130_fd_sc_hd__inv_2 _38628_ (.A(_11072_),
    .Y(_11073_));
 sky130_fd_sc_hd__nor3_2 _38629_ (.A(_11068_),
    .B(_11071_),
    .C(_11073_),
    .Y(_11074_));
 sky130_fd_sc_hd__o32a_1 _38630_ (.A1(_07340_),
    .A2(_08645_),
    .A3(_11070_),
    .B1(_11073_),
    .B2(_11068_),
    .X(_11076_));
 sky130_fd_sc_hd__o211ai_2 _38631_ (.A1(_11074_),
    .A2(_11076_),
    .B1(_09863_),
    .C1(_09873_),
    .Y(_11077_));
 sky130_fd_sc_hd__a211o_1 _38632_ (.A1(_09863_),
    .A2(_09873_),
    .B1(_11074_),
    .C1(_11076_),
    .X(_11078_));
 sky130_fd_sc_hd__o221a_1 _38633_ (.A1(_07324_),
    .A2(_09865_),
    .B1(_08644_),
    .B2(_08645_),
    .C1(_09867_),
    .X(_11079_));
 sky130_fd_sc_hd__a21oi_1 _38634_ (.A1(_11077_),
    .A2(_11078_),
    .B1(_11079_),
    .Y(_11080_));
 sky130_fd_sc_hd__and3_1 _38635_ (.A(_11078_),
    .B(_11079_),
    .C(_11077_),
    .X(_11081_));
 sky130_fd_sc_hd__nor2_1 _38636_ (.A(_11080_),
    .B(_11081_),
    .Y(_11082_));
 sky130_fd_sc_hd__a311o_2 _38637_ (.A1(_09871_),
    .A2(_09873_),
    .A3(_09876_),
    .B1(_09881_),
    .C1(_11082_),
    .X(_11083_));
 sky130_fd_sc_hd__o21ai_1 _38638_ (.A1(_09879_),
    .A2(_09881_),
    .B1(_11082_),
    .Y(_11084_));
 sky130_fd_sc_hd__nand2_1 _38639_ (.A(_11083_),
    .B(_11084_),
    .Y(_11085_));
 sky130_fd_sc_hd__a21oi_1 _38640_ (.A1(_09892_),
    .A2(_09891_),
    .B1(_09885_),
    .Y(_11087_));
 sky130_fd_sc_hd__xor2_2 _38641_ (.A(_11085_),
    .B(_11087_),
    .X(_11088_));
 sky130_fd_sc_hd__nand3_2 _38642_ (.A(_11088_),
    .B(_11045_),
    .C(_11046_),
    .Y(_11089_));
 sky130_fd_sc_hd__a21oi_2 _38643_ (.A1(_09918_),
    .A2(_09950_),
    .B1(_09993_),
    .Y(_11090_));
 sky130_fd_sc_hd__o21bai_1 _38644_ (.A1(_09983_),
    .A2(_09988_),
    .B1_N(_09984_),
    .Y(_11091_));
 sky130_fd_sc_hd__a21o_1 _38645_ (.A1(_09956_),
    .A2(_09978_),
    .B1(_09975_),
    .X(_11092_));
 sky130_fd_sc_hd__buf_1 _38646_ (.A(_09970_),
    .X(_11093_));
 sky130_fd_sc_hd__o211a_1 _38647_ (.A1(_09969_),
    .A2(_11093_),
    .B1(_08529_),
    .C1(_09971_),
    .X(_11094_));
 sky130_fd_sc_hd__o21ba_1 _38648_ (.A1(_02498_),
    .A2(_08540_),
    .B1_N(_08529_),
    .X(_11095_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38649_ (.A(_05747_),
    .X(_11096_));
 sky130_fd_sc_hd__a21oi_1 _38650_ (.A1(_03885_),
    .A2(_11096_),
    .B1(_02494_),
    .Y(_11098_));
 sky130_fd_sc_hd__nor2_1 _38651_ (.A(\delay_line[16][13] ),
    .B(net380),
    .Y(_11099_));
 sky130_fd_sc_hd__and2_1 _38652_ (.A(\delay_line[16][13] ),
    .B(net380),
    .X(_11100_));
 sky130_fd_sc_hd__o21ai_1 _38653_ (.A1(_11099_),
    .A2(_11100_),
    .B1(_03885_),
    .Y(_11101_));
 sky130_fd_sc_hd__or3_2 _38654_ (.A(_08535_),
    .B(_11099_),
    .C(_11100_),
    .X(_11102_));
 sky130_fd_sc_hd__nand2_1 _38655_ (.A(_11101_),
    .B(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__a21oi_1 _38656_ (.A1(_09966_),
    .A2(_09958_),
    .B1(_11103_),
    .Y(_11104_));
 sky130_fd_sc_hd__and3_1 _38657_ (.A(_09964_),
    .B(_11103_),
    .C(\delay_line[16][15] ),
    .X(_11105_));
 sky130_fd_sc_hd__o22a_1 _38658_ (.A1(_09960_),
    .A2(_11098_),
    .B1(_11104_),
    .B2(_11105_),
    .X(_11106_));
 sky130_fd_sc_hd__inv_2 _38659_ (.A(_11106_),
    .Y(_11107_));
 sky130_fd_sc_hd__or4_1 _38660_ (.A(_09960_),
    .B(_11098_),
    .C(_11104_),
    .D(_11105_),
    .X(_11109_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38661_ (.A(_09958_),
    .X(_11110_));
 sky130_fd_sc_hd__nand2_1 _38662_ (.A(_09966_),
    .B(_11110_),
    .Y(_11111_));
 sky130_fd_sc_hd__o21ai_1 _38663_ (.A1(_08543_),
    .A2(_11111_),
    .B1(_09973_),
    .Y(_11112_));
 sky130_fd_sc_hd__nand3_1 _38664_ (.A(_11107_),
    .B(_11109_),
    .C(_11112_),
    .Y(_11113_));
 sky130_fd_sc_hd__a21oi_1 _38665_ (.A1(_11107_),
    .A2(_11109_),
    .B1(_11112_),
    .Y(_11114_));
 sky130_fd_sc_hd__inv_2 _38666_ (.A(_11114_),
    .Y(_11115_));
 sky130_fd_sc_hd__or4bb_1 _38667_ (.A(_11094_),
    .B(_11095_),
    .C_N(_11113_),
    .D_N(_11115_),
    .X(_11116_));
 sky130_fd_sc_hd__a2bb2o_1 _38668_ (.A1_N(_11094_),
    .A2_N(_11095_),
    .B1(_11113_),
    .B2(_11115_),
    .X(_11117_));
 sky130_fd_sc_hd__nand2_1 _38669_ (.A(_11116_),
    .B(_11117_),
    .Y(_11118_));
 sky130_fd_sc_hd__xnor2_1 _38670_ (.A(_11092_),
    .B(_11118_),
    .Y(_11120_));
 sky130_fd_sc_hd__xnor2_1 _38671_ (.A(_09955_),
    .B(_11120_),
    .Y(_11121_));
 sky130_fd_sc_hd__nor2_1 _38672_ (.A(_09980_),
    .B(_09979_),
    .Y(_11122_));
 sky130_fd_sc_hd__a41o_1 _38673_ (.A1(_05740_),
    .A2(_09981_),
    .A3(_03874_),
    .A4(_08529_),
    .B1(_11122_),
    .X(_11123_));
 sky130_fd_sc_hd__and2b_1 _38674_ (.A_N(_11121_),
    .B(_11123_),
    .X(_11124_));
 sky130_fd_sc_hd__and2b_1 _38675_ (.A_N(_11123_),
    .B(_11121_),
    .X(_11125_));
 sky130_fd_sc_hd__nor2_1 _38676_ (.A(_11124_),
    .B(_11125_),
    .Y(_11126_));
 sky130_fd_sc_hd__xnor2_1 _38677_ (.A(_11091_),
    .B(_11126_),
    .Y(_11127_));
 sky130_fd_sc_hd__a21o_1 _38678_ (.A1(_08619_),
    .A2(_08625_),
    .B1(_09946_),
    .X(_11128_));
 sky130_fd_sc_hd__o211ai_2 _38679_ (.A1(_05823_),
    .A2(_08611_),
    .B1(_09922_),
    .C1(_09938_),
    .Y(_11129_));
 sky130_fd_sc_hd__buf_1 _38680_ (.A(_09930_),
    .X(_11131_));
 sky130_fd_sc_hd__and3b_1 _38681_ (.A_N(_11131_),
    .B(_08611_),
    .C(_09922_),
    .X(_11132_));
 sky130_fd_sc_hd__o2bb2a_1 _38682_ (.A1_N(_09925_),
    .A2_N(_05809_),
    .B1(_07251_),
    .B2(_07252_),
    .X(_11133_));
 sky130_fd_sc_hd__and3_1 _38683_ (.A(_09925_),
    .B(_05809_),
    .C(_08606_),
    .X(_11134_));
 sky130_fd_sc_hd__nor2_1 _38684_ (.A(_00775_),
    .B(_00778_),
    .Y(_11135_));
 sky130_fd_sc_hd__nor2_1 _38685_ (.A(_09930_),
    .B(_08597_),
    .Y(_11136_));
 sky130_fd_sc_hd__a21o_1 _38686_ (.A1(_09930_),
    .A2(_11135_),
    .B1(_11136_),
    .X(_11137_));
 sky130_fd_sc_hd__or3_1 _38687_ (.A(_11133_),
    .B(_11134_),
    .C(_11137_),
    .X(_11138_));
 sky130_fd_sc_hd__o21ai_1 _38688_ (.A1(_11133_),
    .A2(_11134_),
    .B1(_11137_),
    .Y(_11139_));
 sky130_fd_sc_hd__o211a_1 _38689_ (.A1(_09934_),
    .A2(_09935_),
    .B1(_11138_),
    .C1(_11139_),
    .X(_11140_));
 sky130_fd_sc_hd__a211oi_1 _38690_ (.A1(_11138_),
    .A2(_11139_),
    .B1(_09934_),
    .C1(_09935_),
    .Y(_11142_));
 sky130_fd_sc_hd__nor4_1 _38691_ (.A(_24740_),
    .B(_11132_),
    .C(_11140_),
    .D(_11142_),
    .Y(_11143_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38692_ (.A(_11140_),
    .X(_11144_));
 sky130_fd_sc_hd__o22a_1 _38693_ (.A1(_11132_),
    .A2(_24740_),
    .B1(_11142_),
    .B2(_11144_),
    .X(_11145_));
 sky130_fd_sc_hd__a211oi_2 _38694_ (.A1(_09937_),
    .A2(_11129_),
    .B1(net165),
    .C1(_11145_),
    .Y(_11146_));
 sky130_fd_sc_hd__o211a_1 _38695_ (.A1(net165),
    .A2(_11145_),
    .B1(_09937_),
    .C1(_11129_),
    .X(_11147_));
 sky130_fd_sc_hd__nor3_1 _38696_ (.A(_09923_),
    .B(_11146_),
    .C(_11147_),
    .Y(_11148_));
 sky130_fd_sc_hd__o21a_1 _38697_ (.A1(_11146_),
    .A2(_11147_),
    .B1(_09923_),
    .X(_11149_));
 sky130_fd_sc_hd__a21boi_1 _38698_ (.A1(_08595_),
    .A2(_09941_),
    .B1_N(_09942_),
    .Y(_11150_));
 sky130_fd_sc_hd__or3b_1 _38699_ (.A(_11148_),
    .B(_11149_),
    .C_N(_11150_),
    .X(_11151_));
 sky130_fd_sc_hd__o21bai_1 _38700_ (.A1(_11148_),
    .A2(_11149_),
    .B1_N(_11150_),
    .Y(_11153_));
 sky130_fd_sc_hd__nand2_1 _38701_ (.A(_11151_),
    .B(_11153_),
    .Y(_11154_));
 sky130_fd_sc_hd__nand3_1 _38702_ (.A(_11128_),
    .B(_09948_),
    .C(_11154_),
    .Y(_11155_));
 sky130_fd_sc_hd__a21o_1 _38703_ (.A1(_11128_),
    .A2(_09948_),
    .B1(_11154_),
    .X(_11156_));
 sky130_fd_sc_hd__buf_1 _38704_ (.A(_09897_),
    .X(_11157_));
 sky130_fd_sc_hd__clkbuf_2 _38705_ (.A(_11157_),
    .X(_11158_));
 sky130_fd_sc_hd__buf_1 _38706_ (.A(_09902_),
    .X(_11159_));
 sky130_fd_sc_hd__buf_1 _38707_ (.A(net388),
    .X(_11160_));
 sky130_fd_sc_hd__and3b_1 _38708_ (.A_N(_11159_),
    .B(_08573_),
    .C(_11160_),
    .X(_11161_));
 sky130_fd_sc_hd__clkbuf_2 _38709_ (.A(\delay_line[14][12] ),
    .X(_11162_));
 sky130_fd_sc_hd__clkbuf_2 _38710_ (.A(_07293_),
    .X(_11164_));
 sky130_fd_sc_hd__xor2_2 _38711_ (.A(_11162_),
    .B(_11164_),
    .X(_11165_));
 sky130_fd_sc_hd__o21a_1 _38712_ (.A1(_09901_),
    .A2(_11159_),
    .B1(_11165_),
    .X(_11166_));
 sky130_fd_sc_hd__nor3_1 _38713_ (.A(_09901_),
    .B(_11159_),
    .C(_11165_),
    .Y(_11167_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38714_ (.A(_11162_),
    .X(_11168_));
 sky130_fd_sc_hd__nand3_1 _38715_ (.A(_08568_),
    .B(_11157_),
    .C(_11168_),
    .Y(_11169_));
 sky130_fd_sc_hd__a21o_1 _38716_ (.A1(_09897_),
    .A2(_11168_),
    .B1(_08568_),
    .X(_11170_));
 sky130_fd_sc_hd__o211ai_2 _38717_ (.A1(_11166_),
    .A2(_11167_),
    .B1(_11169_),
    .C1(_11170_),
    .Y(_11171_));
 sky130_fd_sc_hd__a211o_1 _38718_ (.A1(_11169_),
    .A2(_11170_),
    .B1(_11166_),
    .C1(_11167_),
    .X(_11172_));
 sky130_fd_sc_hd__o211ai_2 _38719_ (.A1(_09906_),
    .A2(_11161_),
    .B1(_11171_),
    .C1(_11172_),
    .Y(_11173_));
 sky130_fd_sc_hd__a211o_1 _38720_ (.A1(_11172_),
    .A2(_11171_),
    .B1(_11161_),
    .C1(_09906_),
    .X(_11175_));
 sky130_fd_sc_hd__a32o_1 _38721_ (.A1(_07285_),
    .A2(_08570_),
    .A3(_11158_),
    .B1(_11173_),
    .B2(_11175_),
    .X(_11176_));
 sky130_fd_sc_hd__nand2_1 _38722_ (.A(_11175_),
    .B(_09900_),
    .Y(_11177_));
 sky130_fd_sc_hd__nand2_1 _38723_ (.A(_11176_),
    .B(_11177_),
    .Y(_11178_));
 sky130_fd_sc_hd__a31o_1 _38724_ (.A1(_03923_),
    .A2(_07290_),
    .A3(_09909_),
    .B1(_09908_),
    .X(_11179_));
 sky130_fd_sc_hd__xnor2_1 _38725_ (.A(_11178_),
    .B(_11179_),
    .Y(_11180_));
 sky130_fd_sc_hd__o21ba_1 _38726_ (.A1(_09917_),
    .A2(_09896_),
    .B1_N(_11180_),
    .X(_11181_));
 sky130_fd_sc_hd__nand3_1 _38727_ (.A(_08566_),
    .B(_08587_),
    .C(_08588_),
    .Y(_11182_));
 sky130_fd_sc_hd__a21o_1 _38728_ (.A1(_08587_),
    .A2(_11182_),
    .B1(_09917_),
    .X(_11183_));
 sky130_fd_sc_hd__a21boi_1 _38729_ (.A1(_09915_),
    .A2(_11183_),
    .B1_N(_11180_),
    .Y(_11184_));
 sky130_fd_sc_hd__a21oi_2 _38730_ (.A1(_11181_),
    .A2(_09915_),
    .B1(_11184_),
    .Y(_11186_));
 sky130_fd_sc_hd__a21oi_1 _38731_ (.A1(_11155_),
    .A2(_11156_),
    .B1(_11186_),
    .Y(_11187_));
 sky130_fd_sc_hd__and3_1 _38732_ (.A(_11186_),
    .B(_11156_),
    .C(_11155_),
    .X(_11188_));
 sky130_fd_sc_hd__nor3_2 _38733_ (.A(_11127_),
    .B(_11187_),
    .C(_11188_),
    .Y(_11189_));
 sky130_fd_sc_hd__o21a_1 _38734_ (.A1(_11188_),
    .A2(_11187_),
    .B1(_11127_),
    .X(_11190_));
 sky130_fd_sc_hd__or3_4 _38735_ (.A(_11090_),
    .B(_11189_),
    .C(_11190_),
    .X(_11191_));
 sky130_fd_sc_hd__o21ai_4 _38736_ (.A1(_11189_),
    .A2(_11190_),
    .B1(_11090_),
    .Y(_11192_));
 sky130_fd_sc_hd__o2111ai_4 _38737_ (.A1(_11047_),
    .A2(_11088_),
    .B1(_11089_),
    .C1(_11191_),
    .D1(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__o21a_1 _38738_ (.A1(_11088_),
    .A2(_11047_),
    .B1(_11089_),
    .X(_11194_));
 sky130_fd_sc_hd__a21o_4 _38739_ (.A1(_11191_),
    .A2(_11192_),
    .B1(_11194_),
    .X(_11195_));
 sky130_fd_sc_hd__a21oi_1 _38740_ (.A1(_11193_),
    .A2(_11195_),
    .B1(net81),
    .Y(_11197_));
 sky130_fd_sc_hd__a211o_1 _38741_ (.A1(_09794_),
    .A2(_09841_),
    .B1(_09890_),
    .C1(_09893_),
    .X(_11198_));
 sky130_fd_sc_hd__o21a_4 _38742_ (.A1(_09794_),
    .A2(_09841_),
    .B1(_11198_),
    .X(_11199_));
 sky130_fd_sc_hd__and2_1 _38743_ (.A(_10001_),
    .B(_10027_),
    .X(_11200_));
 sky130_fd_sc_hd__o21bai_1 _38744_ (.A1(_08407_),
    .A2(_10024_),
    .B1_N(_10023_),
    .Y(_11201_));
 sky130_fd_sc_hd__buf_1 _38745_ (.A(_08410_),
    .X(_11202_));
 sky130_fd_sc_hd__a2111oi_1 _38746_ (.A1(_08402_),
    .A2(_11202_),
    .B1(_10002_),
    .C1(_10018_),
    .D1(_10019_),
    .Y(_11203_));
 sky130_fd_sc_hd__clkbuf_2 _38747_ (.A(_05867_),
    .X(_11204_));
 sky130_fd_sc_hd__buf_1 _38748_ (.A(_10010_),
    .X(_11205_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38749_ (.A(_08411_),
    .X(_11206_));
 sky130_fd_sc_hd__a32o_1 _38750_ (.A1(_11205_),
    .A2(_11206_),
    .A3(_10008_),
    .B1(_07080_),
    .B2(_07082_),
    .X(_11208_));
 sky130_fd_sc_hd__buf_1 _38751_ (.A(_05868_),
    .X(_11209_));
 sky130_fd_sc_hd__or3b_2 _38752_ (.A(_11209_),
    .B(_08413_),
    .C_N(_11205_),
    .X(_11210_));
 sky130_fd_sc_hd__or3b_2 _38753_ (.A(_00473_),
    .B(_00476_),
    .C_N(_10004_),
    .X(_11211_));
 sky130_fd_sc_hd__o2111ai_4 _38754_ (.A1(_10004_),
    .A2(_11204_),
    .B1(_11208_),
    .C1(_11210_),
    .D1(_11211_),
    .Y(_11212_));
 sky130_fd_sc_hd__or2_1 _38755_ (.A(_10004_),
    .B(_11204_),
    .X(_11213_));
 sky130_fd_sc_hd__a22o_1 _38756_ (.A1(_11208_),
    .A2(_11210_),
    .B1(_11211_),
    .B2(_11213_),
    .X(_11214_));
 sky130_fd_sc_hd__o211a_1 _38757_ (.A1(_10013_),
    .A2(_10015_),
    .B1(_11212_),
    .C1(_11214_),
    .X(_11215_));
 sky130_fd_sc_hd__a211o_1 _38758_ (.A1(_11212_),
    .A2(_11214_),
    .B1(_10013_),
    .C1(_10015_),
    .X(_11216_));
 sky130_fd_sc_hd__and2b_1 _38759_ (.A_N(_11215_),
    .B(_11216_),
    .X(_11217_));
 sky130_fd_sc_hd__buf_1 _38760_ (.A(_10004_),
    .X(_11219_));
 sky130_fd_sc_hd__o21ai_1 _38761_ (.A1(_11219_),
    .A2(_10002_),
    .B1(_10005_),
    .Y(_11220_));
 sky130_fd_sc_hd__xnor2_1 _38762_ (.A(_11217_),
    .B(_11220_),
    .Y(_11221_));
 sky130_fd_sc_hd__nor3_1 _38763_ (.A(_10018_),
    .B(net153),
    .C(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__o21a_1 _38764_ (.A1(_10018_),
    .A2(net152),
    .B1(_11221_),
    .X(_11223_));
 sky130_fd_sc_hd__nor2_1 _38765_ (.A(_11222_),
    .B(_11223_),
    .Y(_11224_));
 sky130_fd_sc_hd__xor2_1 _38766_ (.A(_10003_),
    .B(_11224_),
    .X(_11225_));
 sky130_fd_sc_hd__nor2_1 _38767_ (.A(_11201_),
    .B(_11225_),
    .Y(_11226_));
 sky130_fd_sc_hd__nand2_1 _38768_ (.A(_11225_),
    .B(_11201_),
    .Y(_11227_));
 sky130_fd_sc_hd__and2b_1 _38769_ (.A_N(_11226_),
    .B(_11227_),
    .X(_11228_));
 sky130_fd_sc_hd__or3_1 _38770_ (.A(_11200_),
    .B(_10029_),
    .C(_11228_),
    .X(_11230_));
 sky130_fd_sc_hd__o21ai_1 _38771_ (.A1(_11200_),
    .A2(_10029_),
    .B1(_11228_),
    .Y(_11231_));
 sky130_fd_sc_hd__a21boi_2 _38772_ (.A1(_10066_),
    .A2(_10069_),
    .B1_N(_10067_),
    .Y(_11232_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38773_ (.A(_10047_),
    .X(_11233_));
 sky130_fd_sc_hd__nand3_1 _38774_ (.A(_11233_),
    .B(_10034_),
    .C(_10033_),
    .Y(_11234_));
 sky130_fd_sc_hd__o21ai_1 _38775_ (.A1(_10039_),
    .A2(_08455_),
    .B1(_10049_),
    .Y(_11235_));
 sky130_fd_sc_hd__clkbuf_2 _38776_ (.A(_07121_),
    .X(_11236_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38777_ (.A(_00518_),
    .X(_11237_));
 sky130_fd_sc_hd__o21a_1 _38778_ (.A1(_08450_),
    .A2(_10047_),
    .B1(_11237_),
    .X(_11238_));
 sky130_fd_sc_hd__nor3_1 _38779_ (.A(_08450_),
    .B(_11237_),
    .C(_10047_),
    .Y(_11239_));
 sky130_fd_sc_hd__nor2_1 _38780_ (.A(_11236_),
    .B(_10037_),
    .Y(_11241_));
 sky130_fd_sc_hd__and2_1 _38781_ (.A(_07121_),
    .B(net350),
    .X(_11242_));
 sky130_fd_sc_hd__a2bb2o_1 _38782_ (.A1_N(_11241_),
    .A2_N(_11242_),
    .B1(_04179_),
    .B2(_10038_),
    .X(_11243_));
 sky130_fd_sc_hd__o221ai_4 _38783_ (.A1(_11236_),
    .A2(_10040_),
    .B1(_11238_),
    .B2(net263),
    .C1(_11243_),
    .Y(_11244_));
 sky130_fd_sc_hd__or3b_1 _38784_ (.A(_11236_),
    .B(_10044_),
    .C_N(_04179_),
    .X(_11245_));
 sky130_fd_sc_hd__a211o_1 _38785_ (.A1(_11243_),
    .A2(_11245_),
    .B1(_11238_),
    .C1(_11239_),
    .X(_11246_));
 sky130_fd_sc_hd__and4_1 _38786_ (.A(_10043_),
    .B(_11235_),
    .C(_11244_),
    .D(_11246_),
    .X(_11247_));
 sky130_fd_sc_hd__a22o_1 _38787_ (.A1(_10043_),
    .A2(_11235_),
    .B1(_11244_),
    .B2(_11246_),
    .X(_11248_));
 sky130_fd_sc_hd__inv_2 _38788_ (.A(_11248_),
    .Y(_11249_));
 sky130_fd_sc_hd__o2bb2a_1 _38789_ (.A1_N(_10057_),
    .A2_N(_11234_),
    .B1(_11247_),
    .B2(_11249_),
    .X(_11250_));
 sky130_fd_sc_hd__and4b_1 _38790_ (.A_N(_11247_),
    .B(_10057_),
    .C(_11234_),
    .D(_11248_),
    .X(_11252_));
 sky130_fd_sc_hd__a211o_1 _38791_ (.A1(_10055_),
    .A2(_10058_),
    .B1(_11250_),
    .C1(_11252_),
    .X(_11253_));
 sky130_fd_sc_hd__and3b_1 _38792_ (.A_N(_10057_),
    .B(_10033_),
    .C(_20450_),
    .X(_11254_));
 sky130_fd_sc_hd__nand2_1 _38793_ (.A(_10055_),
    .B(_10058_),
    .Y(_11255_));
 sky130_fd_sc_hd__nor2_1 _38794_ (.A(_11250_),
    .B(_11252_),
    .Y(_11256_));
 sky130_fd_sc_hd__or2_1 _38795_ (.A(_11255_),
    .B(_11256_),
    .X(_11257_));
 sky130_fd_sc_hd__nand3_1 _38796_ (.A(_11253_),
    .B(_11254_),
    .C(_11257_),
    .Y(_11258_));
 sky130_fd_sc_hd__inv_2 _38797_ (.A(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__a21oi_1 _38798_ (.A1(_11257_),
    .A2(_11253_),
    .B1(_11254_),
    .Y(_11260_));
 sky130_fd_sc_hd__a21boi_1 _38799_ (.A1(_10060_),
    .A2(_08449_),
    .B1_N(_10061_),
    .Y(_11261_));
 sky130_fd_sc_hd__nor3_1 _38800_ (.A(_11259_),
    .B(_11260_),
    .C(_11261_),
    .Y(_11263_));
 sky130_fd_sc_hd__o21a_1 _38801_ (.A1(_11259_),
    .A2(_11260_),
    .B1(_11261_),
    .X(_11264_));
 sky130_fd_sc_hd__or2_1 _38802_ (.A(_11263_),
    .B(_11264_),
    .X(_11265_));
 sky130_fd_sc_hd__xnor2_2 _38803_ (.A(_11232_),
    .B(_11265_),
    .Y(_11266_));
 sky130_fd_sc_hd__nand2_1 _38804_ (.A(_10098_),
    .B(_10100_),
    .Y(_11267_));
 sky130_fd_sc_hd__buf_1 _38805_ (.A(_10087_),
    .X(_11268_));
 sky130_fd_sc_hd__buf_1 _38806_ (.A(_07167_),
    .X(_11269_));
 sky130_fd_sc_hd__o211a_1 _38807_ (.A1(_10074_),
    .A2(_11268_),
    .B1(_07171_),
    .C1(_11269_),
    .X(_11270_));
 sky130_fd_sc_hd__o21ba_1 _38808_ (.A1(_08484_),
    .A2(_08483_),
    .B1_N(_07171_),
    .X(_11271_));
 sky130_fd_sc_hd__a21oi_1 _38809_ (.A1(_10087_),
    .A2(_07164_),
    .B1(_02322_),
    .Y(_11272_));
 sky130_fd_sc_hd__nor2_1 _38810_ (.A(\delay_line[24][13] ),
    .B(\delay_line[24][14] ),
    .Y(_11274_));
 sky130_fd_sc_hd__and2_1 _38811_ (.A(\delay_line[24][13] ),
    .B(\delay_line[24][14] ),
    .X(_11275_));
 sky130_fd_sc_hd__o21ai_1 _38812_ (.A1(_11274_),
    .A2(_11275_),
    .B1(_04214_),
    .Y(_11276_));
 sky130_fd_sc_hd__or3_1 _38813_ (.A(_04213_),
    .B(_11274_),
    .C(_11275_),
    .X(_11277_));
 sky130_fd_sc_hd__nand2_1 _38814_ (.A(_11276_),
    .B(_11277_),
    .Y(_11278_));
 sky130_fd_sc_hd__a21oi_1 _38815_ (.A1(_10083_),
    .A2(_08488_),
    .B1(_11278_),
    .Y(_11279_));
 sky130_fd_sc_hd__and3_1 _38816_ (.A(_10082_),
    .B(_11278_),
    .C(\delay_line[24][15] ),
    .X(_11280_));
 sky130_fd_sc_hd__o22a_1 _38817_ (.A1(_10080_),
    .A2(_11272_),
    .B1(_11279_),
    .B2(_11280_),
    .X(_11281_));
 sky130_fd_sc_hd__inv_2 _38818_ (.A(_11281_),
    .Y(_11282_));
 sky130_fd_sc_hd__or4_1 _38819_ (.A(_10080_),
    .B(_11272_),
    .C(_11279_),
    .D(_11280_),
    .X(_11283_));
 sky130_fd_sc_hd__or3b_1 _38820_ (.A(_08482_),
    .B(_08487_),
    .C_N(_10083_),
    .X(_11285_));
 sky130_fd_sc_hd__nand2_1 _38821_ (.A(_10089_),
    .B(_11285_),
    .Y(_11286_));
 sky130_fd_sc_hd__nand3_1 _38822_ (.A(_11282_),
    .B(_11283_),
    .C(_11286_),
    .Y(_11287_));
 sky130_fd_sc_hd__inv_2 _38823_ (.A(_11287_),
    .Y(_11288_));
 sky130_fd_sc_hd__a21oi_1 _38824_ (.A1(_11282_),
    .A2(_11283_),
    .B1(_11286_),
    .Y(_11289_));
 sky130_fd_sc_hd__or4_2 _38825_ (.A(_11270_),
    .B(_11271_),
    .C(_11288_),
    .D(_11289_),
    .X(_11290_));
 sky130_fd_sc_hd__o22ai_2 _38826_ (.A1(_11270_),
    .A2(_11271_),
    .B1(_11288_),
    .B2(_11289_),
    .Y(_11291_));
 sky130_fd_sc_hd__a211oi_1 _38827_ (.A1(_11290_),
    .A2(_11291_),
    .B1(_10092_),
    .C1(net154),
    .Y(_11292_));
 sky130_fd_sc_hd__inv_2 _38828_ (.A(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__o211ai_2 _38829_ (.A1(_10092_),
    .A2(net154),
    .B1(_11290_),
    .C1(_11291_),
    .Y(_11294_));
 sky130_fd_sc_hd__nand4_1 _38830_ (.A(_11293_),
    .B(_11294_),
    .C(_05961_),
    .D(_08491_),
    .Y(_11296_));
 sky130_fd_sc_hd__a22o_1 _38831_ (.A1(_05961_),
    .A2(_08491_),
    .B1(_11293_),
    .B2(_11294_),
    .X(_11297_));
 sky130_fd_sc_hd__nand2_1 _38832_ (.A(_11296_),
    .B(_11297_),
    .Y(_11298_));
 sky130_fd_sc_hd__xnor2_2 _38833_ (.A(_11267_),
    .B(_11298_),
    .Y(_11299_));
 sky130_fd_sc_hd__o22ai_4 _38834_ (.A1(_10103_),
    .A2(_10101_),
    .B1(_10105_),
    .B2(_10106_),
    .Y(_11300_));
 sky130_fd_sc_hd__xor2_2 _38835_ (.A(_11299_),
    .B(_11300_),
    .X(_11301_));
 sky130_fd_sc_hd__xnor2_1 _38836_ (.A(_11266_),
    .B(_11301_),
    .Y(_11302_));
 sky130_fd_sc_hd__a21oi_1 _38837_ (.A1(_11230_),
    .A2(_11231_),
    .B1(_11302_),
    .Y(_11303_));
 sky130_fd_sc_hd__nand3_1 _38838_ (.A(_11302_),
    .B(_11231_),
    .C(_11230_),
    .Y(_11304_));
 sky130_fd_sc_hd__inv_2 _38839_ (.A(_11304_),
    .Y(_11305_));
 sky130_fd_sc_hd__nor3_1 _38840_ (.A(_11199_),
    .B(_11303_),
    .C(_11305_),
    .Y(_11307_));
 sky130_fd_sc_hd__o21ai_1 _38841_ (.A1(_11303_),
    .A2(_11305_),
    .B1(_11199_),
    .Y(_11308_));
 sky130_fd_sc_hd__and2b_1 _38842_ (.A_N(_11307_),
    .B(_11308_),
    .X(_11309_));
 sky130_fd_sc_hd__o21ai_2 _38843_ (.A1(_10032_),
    .A2(_10112_),
    .B1(_10110_),
    .Y(_11310_));
 sky130_fd_sc_hd__xnor2_1 _38844_ (.A(_11309_),
    .B(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__or2_1 _38845_ (.A(_11197_),
    .B(_11311_),
    .X(_11312_));
 sky130_fd_sc_hd__a31o_1 _38846_ (.A1(net81),
    .A2(_11193_),
    .A3(_11195_),
    .B1(_11312_),
    .X(_11313_));
 sky130_fd_sc_hd__nand3_1 _38847_ (.A(net81),
    .B(_11193_),
    .C(_11195_),
    .Y(_11314_));
 sky130_fd_sc_hd__inv_2 _38848_ (.A(_11314_),
    .Y(_11315_));
 sky130_fd_sc_hd__o21ai_1 _38849_ (.A1(_11315_),
    .A2(_11197_),
    .B1(_11311_),
    .Y(_11316_));
 sky130_fd_sc_hd__nor2_1 _38850_ (.A(_09996_),
    .B(_09752_),
    .Y(_11318_));
 sky130_fd_sc_hd__o21ai_2 _38851_ (.A1(_08639_),
    .A2(_08766_),
    .B1(_09996_),
    .Y(_11319_));
 sky130_fd_sc_hd__o21ai_4 _38852_ (.A1(_11318_),
    .A2(_10120_),
    .B1(_11319_),
    .Y(_11320_));
 sky130_fd_sc_hd__a21o_1 _38853_ (.A1(_11313_),
    .A2(_11316_),
    .B1(_11320_),
    .X(_11321_));
 sky130_fd_sc_hd__a21oi_2 _38854_ (.A1(_10116_),
    .A2(_10118_),
    .B1(_10114_),
    .Y(_11322_));
 sky130_fd_sc_hd__inv_2 _38855_ (.A(_10166_),
    .Y(_11323_));
 sky130_fd_sc_hd__o21a_1 _38856_ (.A1(_10178_),
    .A2(_11323_),
    .B1(_10165_),
    .X(_11324_));
 sky130_fd_sc_hd__nor2_1 _38857_ (.A(_06999_),
    .B(_10170_),
    .Y(_11325_));
 sky130_fd_sc_hd__o21a_1 _38858_ (.A1(_04266_),
    .A2(_10168_),
    .B1(_06999_),
    .X(_11326_));
 sky130_fd_sc_hd__o211ai_1 _38859_ (.A1(_11325_),
    .A2(_11326_),
    .B1(_08785_),
    .C1(_10172_),
    .Y(_11327_));
 sky130_fd_sc_hd__a211o_1 _38860_ (.A1(_08785_),
    .A2(_10172_),
    .B1(_11325_),
    .C1(_11326_),
    .X(_11329_));
 sky130_fd_sc_hd__and4bb_1 _38861_ (.A_N(_10173_),
    .B_N(_10175_),
    .C(_11327_),
    .D(_11329_),
    .X(_11330_));
 sky130_fd_sc_hd__o2bb2a_1 _38862_ (.A1_N(_11327_),
    .A2_N(_11329_),
    .B1(_10173_),
    .B2(_10175_),
    .X(_11331_));
 sky130_fd_sc_hd__or2_1 _38863_ (.A(_11330_),
    .B(_11331_),
    .X(_11332_));
 sky130_fd_sc_hd__or2b_1 _38864_ (.A(_08793_),
    .B_N(_10176_),
    .X(_11333_));
 sky130_fd_sc_hd__o21a_1 _38865_ (.A1(_10177_),
    .A2(_10167_),
    .B1(_11333_),
    .X(_11334_));
 sky130_fd_sc_hd__xnor2_2 _38866_ (.A(_11332_),
    .B(_11334_),
    .Y(_11335_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38867_ (.A(_08803_),
    .X(_11336_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38868_ (.A(net336),
    .X(_11337_));
 sky130_fd_sc_hd__nor2_1 _38869_ (.A(_11337_),
    .B(net335),
    .Y(_11338_));
 sky130_fd_sc_hd__and2_1 _38870_ (.A(net336),
    .B(net335),
    .X(_11340_));
 sky130_fd_sc_hd__or3b_2 _38871_ (.A(_11338_),
    .B(_11340_),
    .C_N(_24337_),
    .X(_11341_));
 sky130_fd_sc_hd__o21bai_1 _38872_ (.A1(_11338_),
    .A2(_11340_),
    .B1_N(_24337_),
    .Y(_11342_));
 sky130_fd_sc_hd__o211a_1 _38873_ (.A1(_10149_),
    .A2(_10150_),
    .B1(_11341_),
    .C1(_11342_),
    .X(_11343_));
 sky130_fd_sc_hd__a221oi_2 _38874_ (.A1(_10146_),
    .A2(_11337_),
    .B1(_11341_),
    .B2(_11342_),
    .C1(_10150_),
    .Y(_11344_));
 sky130_fd_sc_hd__nor2_1 _38875_ (.A(_11343_),
    .B(_11344_),
    .Y(_11345_));
 sky130_fd_sc_hd__a21oi_1 _38876_ (.A1(_08810_),
    .A2(_10156_),
    .B1(_10154_),
    .Y(_11346_));
 sky130_fd_sc_hd__xor2_1 _38877_ (.A(_11345_),
    .B(_11346_),
    .X(_11347_));
 sky130_fd_sc_hd__xor2_1 _38878_ (.A(_11336_),
    .B(_11347_),
    .X(_11348_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38879_ (.A(_08802_),
    .X(_11349_));
 sky130_fd_sc_hd__a32o_1 _38880_ (.A1(_08814_),
    .A2(_08813_),
    .A3(_10156_),
    .B1(_10158_),
    .B2(_11349_),
    .X(_11351_));
 sky130_fd_sc_hd__nand2_1 _38881_ (.A(_11348_),
    .B(_11351_),
    .Y(_11352_));
 sky130_fd_sc_hd__or2_1 _38882_ (.A(_11351_),
    .B(_11348_),
    .X(_11353_));
 sky130_fd_sc_hd__and2_1 _38883_ (.A(_11352_),
    .B(_11353_),
    .X(_11354_));
 sky130_fd_sc_hd__a21oi_1 _38884_ (.A1(_10160_),
    .A2(_10162_),
    .B1(_11354_),
    .Y(_11355_));
 sky130_fd_sc_hd__and3_1 _38885_ (.A(_10160_),
    .B(_10162_),
    .C(_11354_),
    .X(_11356_));
 sky130_fd_sc_hd__nor2_1 _38886_ (.A(_11355_),
    .B(_11356_),
    .Y(_11357_));
 sky130_fd_sc_hd__a21oi_2 _38887_ (.A1(_05509_),
    .A2(_02221_),
    .B1(_07040_),
    .Y(_11358_));
 sky130_fd_sc_hd__and3_1 _38888_ (.A(_07040_),
    .B(_05509_),
    .C(_02221_),
    .X(_11359_));
 sky130_fd_sc_hd__a2111oi_1 _38889_ (.A1(_10131_),
    .A2(_00969_),
    .B1(_02228_),
    .C1(_11358_),
    .D1(_11359_),
    .Y(_11360_));
 sky130_fd_sc_hd__a31oi_2 _38890_ (.A1(_23155_),
    .A2(_00972_),
    .A3(_10136_),
    .B1(_10134_),
    .Y(_11362_));
 sky130_fd_sc_hd__o22a_1 _38891_ (.A1(_02228_),
    .A2(_10132_),
    .B1(_11359_),
    .B2(_11358_),
    .X(_11363_));
 sky130_fd_sc_hd__or2_1 _38892_ (.A(_11362_),
    .B(_11363_),
    .X(_11364_));
 sky130_fd_sc_hd__o21ai_1 _38893_ (.A1(_11363_),
    .A2(net192),
    .B1(_11362_),
    .Y(_11365_));
 sky130_fd_sc_hd__o21a_1 _38894_ (.A1(net191),
    .A2(_11364_),
    .B1(_11365_),
    .X(_11366_));
 sky130_fd_sc_hd__and2_1 _38895_ (.A(_10138_),
    .B(_11366_),
    .X(_11367_));
 sky130_fd_sc_hd__nor2_1 _38896_ (.A(_10138_),
    .B(_11366_),
    .Y(_11368_));
 sky130_fd_sc_hd__nor2_1 _38897_ (.A(_11367_),
    .B(_11368_),
    .Y(_11369_));
 sky130_fd_sc_hd__inv_2 _38898_ (.A(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__o21ba_1 _38899_ (.A1(_08839_),
    .A2(_08842_),
    .B1_N(_10140_),
    .X(_11371_));
 sky130_fd_sc_hd__a31oi_2 _38900_ (.A1(_08846_),
    .A2(_10142_),
    .A3(_08845_),
    .B1(_11371_),
    .Y(_11373_));
 sky130_fd_sc_hd__xor2_1 _38901_ (.A(_11370_),
    .B(_11373_),
    .X(_11374_));
 sky130_fd_sc_hd__and2b_1 _38902_ (.A_N(_11357_),
    .B(_11374_),
    .X(_11375_));
 sky130_fd_sc_hd__and2b_1 _38903_ (.A_N(_11374_),
    .B(_11357_),
    .X(_11376_));
 sky130_fd_sc_hd__or2_1 _38904_ (.A(_11375_),
    .B(_11376_),
    .X(_11377_));
 sky130_fd_sc_hd__xor2_1 _38905_ (.A(_11335_),
    .B(_11377_),
    .X(_11378_));
 sky130_fd_sc_hd__xnor2_1 _38906_ (.A(_11324_),
    .B(_11378_),
    .Y(_11379_));
 sky130_fd_sc_hd__o21ai_1 _38907_ (.A1(_08883_),
    .A2(_08884_),
    .B1(_10260_),
    .Y(_11380_));
 sky130_fd_sc_hd__nand2_1 _38908_ (.A(_11380_),
    .B(_08878_),
    .Y(_11381_));
 sky130_fd_sc_hd__buf_1 _38909_ (.A(_08858_),
    .X(_11382_));
 sky130_fd_sc_hd__or2b_1 _38910_ (.A(_08864_),
    .B_N(_10244_),
    .X(_11384_));
 sky130_fd_sc_hd__or2b_1 _38911_ (.A(_10244_),
    .B_N(_08864_),
    .X(_11385_));
 sky130_fd_sc_hd__nand4_1 _38912_ (.A(_06957_),
    .B(_11384_),
    .C(_11385_),
    .D(_10237_),
    .Y(_11386_));
 sky130_fd_sc_hd__inv_2 _38913_ (.A(_11386_),
    .Y(_11387_));
 sky130_fd_sc_hd__a22o_1 _38914_ (.A1(_06957_),
    .A2(_10237_),
    .B1(_11384_),
    .B2(_11385_),
    .X(_11388_));
 sky130_fd_sc_hd__or3b_1 _38915_ (.A(_11382_),
    .B(_11387_),
    .C_N(_11388_),
    .X(_11389_));
 sky130_fd_sc_hd__nand2_1 _38916_ (.A(_11386_),
    .B(_11388_),
    .Y(_11390_));
 sky130_fd_sc_hd__nand2_1 _38917_ (.A(_11390_),
    .B(_11382_),
    .Y(_11391_));
 sky130_fd_sc_hd__o32a_1 _38918_ (.A1(_08865_),
    .A2(_10236_),
    .A3(_10238_),
    .B1(_10242_),
    .B2(_10235_),
    .X(_11392_));
 sky130_fd_sc_hd__a21oi_2 _38919_ (.A1(_11389_),
    .A2(_11391_),
    .B1(_11392_),
    .Y(_11393_));
 sky130_fd_sc_hd__nand3_1 _38920_ (.A(_11392_),
    .B(_11389_),
    .C(_11391_),
    .Y(_11395_));
 sky130_fd_sc_hd__and2b_1 _38921_ (.A_N(_11393_),
    .B(_11395_),
    .X(_11396_));
 sky130_fd_sc_hd__a211oi_1 _38922_ (.A1(_08867_),
    .A2(_10250_),
    .B1(_11396_),
    .C1(_10249_),
    .Y(_11397_));
 sky130_fd_sc_hd__o21a_1 _38923_ (.A1(_10249_),
    .A2(_10252_),
    .B1(_11396_),
    .X(_11398_));
 sky130_fd_sc_hd__nor2_1 _38924_ (.A(_11397_),
    .B(_11398_),
    .Y(_11399_));
 sky130_fd_sc_hd__and3_1 _38925_ (.A(_11399_),
    .B(_10234_),
    .C(_10254_),
    .X(_11400_));
 sky130_fd_sc_hd__a21oi_1 _38926_ (.A1(_10234_),
    .A2(_10254_),
    .B1(_11399_),
    .Y(_11401_));
 sky130_fd_sc_hd__or2_1 _38927_ (.A(_11400_),
    .B(_11401_),
    .X(_11402_));
 sky130_fd_sc_hd__a21oi_1 _38928_ (.A1(_10261_),
    .A2(_11381_),
    .B1(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__o211ai_1 _38929_ (.A1(_10260_),
    .A2(_10258_),
    .B1(_11381_),
    .C1(_11402_),
    .Y(_11404_));
 sky130_fd_sc_hd__and2b_1 _38930_ (.A_N(_11403_),
    .B(_11404_),
    .X(_11406_));
 sky130_fd_sc_hd__or2_1 _38931_ (.A(_10230_),
    .B(_10231_),
    .X(_11407_));
 sky130_fd_sc_hd__a21bo_1 _38932_ (.A1(_05477_),
    .A2(_10203_),
    .B1_N(_10201_),
    .X(_11408_));
 sky130_fd_sc_hd__and3_1 _38933_ (.A(_10199_),
    .B(net319),
    .C(_10209_),
    .X(_11409_));
 sky130_fd_sc_hd__buf_1 _38934_ (.A(_10199_),
    .X(_11410_));
 sky130_fd_sc_hd__a21oi_1 _38935_ (.A1(_10211_),
    .A2(_10210_),
    .B1(_11410_),
    .Y(_11411_));
 sky130_fd_sc_hd__and3_1 _38936_ (.A(_06924_),
    .B(_08902_),
    .C(_10204_),
    .X(_11412_));
 sky130_fd_sc_hd__clkbuf_2 _38937_ (.A(_02101_),
    .X(_11413_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38938_ (.A(_10206_),
    .X(_11414_));
 sky130_fd_sc_hd__o21a_1 _38939_ (.A1(_11413_),
    .A2(_11414_),
    .B1(_06908_),
    .X(_11415_));
 sky130_fd_sc_hd__nor4_1 _38940_ (.A(_05477_),
    .B(_08895_),
    .C(_11412_),
    .D(_11415_),
    .Y(_11417_));
 sky130_fd_sc_hd__o22a_1 _38941_ (.A1(_05477_),
    .A2(_08895_),
    .B1(_11412_),
    .B2(_11415_),
    .X(_11418_));
 sky130_fd_sc_hd__or4_1 _38942_ (.A(_11409_),
    .B(_11411_),
    .C(net247),
    .D(_11418_),
    .X(_11419_));
 sky130_fd_sc_hd__nor2_1 _38943_ (.A(_11409_),
    .B(_11411_),
    .Y(_11420_));
 sky130_fd_sc_hd__nor2_1 _38944_ (.A(net247),
    .B(_11418_),
    .Y(_11421_));
 sky130_fd_sc_hd__or2_1 _38945_ (.A(_11420_),
    .B(_11421_),
    .X(_11422_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _38946_ (.A(_10217_),
    .X(_11423_));
 sky130_fd_sc_hd__nor4b_1 _38947_ (.A(_10203_),
    .B(_08898_),
    .C(_10210_),
    .D_N(_11423_),
    .Y(_11424_));
 sky130_fd_sc_hd__a211o_1 _38948_ (.A1(_11419_),
    .A2(_11422_),
    .B1(_10215_),
    .C1(net221),
    .X(_11425_));
 sky130_fd_sc_hd__o211ai_1 _38949_ (.A1(_10215_),
    .A2(net221),
    .B1(_11419_),
    .C1(_11422_),
    .Y(_11426_));
 sky130_fd_sc_hd__and3_1 _38950_ (.A(_11408_),
    .B(_11425_),
    .C(_11426_),
    .X(_11428_));
 sky130_fd_sc_hd__a21oi_1 _38951_ (.A1(_11425_),
    .A2(_11426_),
    .B1(_11408_),
    .Y(_11429_));
 sky130_fd_sc_hd__nor2_1 _38952_ (.A(_10220_),
    .B(_10223_),
    .Y(_11430_));
 sky130_fd_sc_hd__or3_1 _38953_ (.A(_11428_),
    .B(_11429_),
    .C(_11430_),
    .X(_11431_));
 sky130_fd_sc_hd__nor2_1 _38954_ (.A(_11428_),
    .B(_11429_),
    .Y(_11432_));
 sky130_fd_sc_hd__or3_1 _38955_ (.A(_10220_),
    .B(_10223_),
    .C(_11432_),
    .X(_11433_));
 sky130_fd_sc_hd__and2_1 _38956_ (.A(_11431_),
    .B(_11433_),
    .X(_11434_));
 sky130_fd_sc_hd__o2bb2a_1 _38957_ (.A1_N(_10227_),
    .A2_N(_11407_),
    .B1(_11434_),
    .B2(_10225_),
    .X(_11435_));
 sky130_fd_sc_hd__a21o_1 _38958_ (.A1(_11431_),
    .A2(_11433_),
    .B1(_10225_),
    .X(_11436_));
 sky130_fd_sc_hd__or4b_2 _38959_ (.A(_10195_),
    .B(_10223_),
    .C(_10224_),
    .D_N(_11434_),
    .X(_11437_));
 sky130_fd_sc_hd__and2_1 _38960_ (.A(_11436_),
    .B(_11437_),
    .X(_11439_));
 sky130_fd_sc_hd__o21ai_1 _38961_ (.A1(_10230_),
    .A2(_10231_),
    .B1(_10227_),
    .Y(_11440_));
 sky130_fd_sc_hd__nor2_1 _38962_ (.A(_11439_),
    .B(_11440_),
    .Y(_11441_));
 sky130_fd_sc_hd__buf_1 _38963_ (.A(\delay_line[29][12] ),
    .X(_11442_));
 sky130_fd_sc_hd__buf_1 _38964_ (.A(\delay_line[29][15] ),
    .X(_11443_));
 sky130_fd_sc_hd__nor2_1 _38965_ (.A(_11442_),
    .B(_11443_),
    .Y(_11444_));
 sky130_fd_sc_hd__and2_1 _38966_ (.A(\delay_line[29][12] ),
    .B(_11443_),
    .X(_11445_));
 sky130_fd_sc_hd__a21o_1 _38967_ (.A1(_08886_),
    .A2(_10186_),
    .B1(_10183_),
    .X(_11446_));
 sky130_fd_sc_hd__o21a_1 _38968_ (.A1(_11444_),
    .A2(_11445_),
    .B1(_11446_),
    .X(_11447_));
 sky130_fd_sc_hd__a2111oi_1 _38969_ (.A1(_08886_),
    .A2(_10186_),
    .B1(_11444_),
    .C1(_11445_),
    .D1(_10183_),
    .Y(_11448_));
 sky130_fd_sc_hd__or4_2 _38970_ (.A(_06943_),
    .B(_10183_),
    .C(_10184_),
    .D(_08889_),
    .X(_11450_));
 sky130_fd_sc_hd__o221a_1 _38971_ (.A1(_10188_),
    .A2(_10190_),
    .B1(_11447_),
    .B2(net262),
    .C1(_11450_),
    .X(_11451_));
 sky130_fd_sc_hd__a211oi_2 _38972_ (.A1(_10192_),
    .A2(_11450_),
    .B1(net262),
    .C1(_11447_),
    .Y(_11452_));
 sky130_fd_sc_hd__or2_1 _38973_ (.A(_11451_),
    .B(_11452_),
    .X(_11453_));
 sky130_fd_sc_hd__o21a_1 _38974_ (.A1(_11435_),
    .A2(_11441_),
    .B1(_11453_),
    .X(_11454_));
 sky130_fd_sc_hd__nor3_2 _38975_ (.A(_11441_),
    .B(_11453_),
    .C(_11435_),
    .Y(_11455_));
 sky130_fd_sc_hd__or3_1 _38976_ (.A(_11406_),
    .B(_11454_),
    .C(_11455_),
    .X(_11456_));
 sky130_fd_sc_hd__o21ai_1 _38977_ (.A1(_11454_),
    .A2(_11455_),
    .B1(_11406_),
    .Y(_11457_));
 sky130_fd_sc_hd__nand2_2 _38978_ (.A(_11456_),
    .B(_11457_),
    .Y(_11458_));
 sky130_fd_sc_hd__xnor2_1 _38979_ (.A(_11379_),
    .B(_11458_),
    .Y(_11459_));
 sky130_fd_sc_hd__or2_1 _38980_ (.A(_11322_),
    .B(_11459_),
    .X(_11461_));
 sky130_fd_sc_hd__nand2_1 _38981_ (.A(_11459_),
    .B(_11322_),
    .Y(_11462_));
 sky130_fd_sc_hd__a221oi_1 _38982_ (.A1(_10128_),
    .A2(_10181_),
    .B1(_11461_),
    .B2(_11462_),
    .C1(_10268_),
    .Y(_11463_));
 sky130_fd_sc_hd__a21oi_1 _38983_ (.A1(_10128_),
    .A2(_10181_),
    .B1(_10268_),
    .Y(_11464_));
 sky130_fd_sc_hd__and3b_1 _38984_ (.A_N(_11464_),
    .B(_11461_),
    .C(_11462_),
    .X(_11465_));
 sky130_fd_sc_hd__nor2_2 _38985_ (.A(_11463_),
    .B(_11465_),
    .Y(_11466_));
 sky130_fd_sc_hd__o211ai_1 _38986_ (.A1(_11315_),
    .A2(_11312_),
    .B1(_11316_),
    .C1(_11320_),
    .Y(_11467_));
 sky130_fd_sc_hd__nand3_1 _38987_ (.A(_11321_),
    .B(_11466_),
    .C(_11467_),
    .Y(_11468_));
 sky130_fd_sc_hd__a21o_1 _38988_ (.A1(_11467_),
    .A2(_11321_),
    .B1(_11466_),
    .X(_11469_));
 sky130_fd_sc_hd__nand2_1 _38989_ (.A(_11468_),
    .B(_11469_),
    .Y(_11470_));
 sky130_fd_sc_hd__xnor2_1 _38990_ (.A(_10971_),
    .B(_11470_),
    .Y(_11472_));
 sky130_fd_sc_hd__o21ba_1 _38991_ (.A1(_09683_),
    .A2(_09681_),
    .B1_N(_09740_),
    .X(_11473_));
 sky130_fd_sc_hd__a21oi_2 _38992_ (.A1(_09683_),
    .A2(_09681_),
    .B1(_11473_),
    .Y(_11474_));
 sky130_fd_sc_hd__a21oi_1 _38993_ (.A1(_08299_),
    .A2(_09652_),
    .B1(_09658_),
    .Y(_11475_));
 sky130_fd_sc_hd__buf_1 _38994_ (.A(_08291_),
    .X(_11476_));
 sky130_fd_sc_hd__buf_1 _38995_ (.A(_06779_),
    .X(_11477_));
 sky130_fd_sc_hd__a21oi_1 _38996_ (.A1(_11476_),
    .A2(_11477_),
    .B1(_08286_),
    .Y(_11478_));
 sky130_fd_sc_hd__and3_1 _38997_ (.A(_08286_),
    .B(_11476_),
    .C(_11477_),
    .X(_11479_));
 sky130_fd_sc_hd__o22a_1 _38998_ (.A1(_09653_),
    .A2(_11475_),
    .B1(_11478_),
    .B2(_11479_),
    .X(_11480_));
 sky130_fd_sc_hd__nor4_1 _38999_ (.A(_09653_),
    .B(_11475_),
    .C(_11478_),
    .D(_11479_),
    .Y(_11481_));
 sky130_fd_sc_hd__nor3_1 _39000_ (.A(_11480_),
    .B(_09651_),
    .C(_11481_),
    .Y(_11483_));
 sky130_fd_sc_hd__o21a_1 _39001_ (.A1(_11481_),
    .A2(_11480_),
    .B1(_09651_),
    .X(_11484_));
 sky130_fd_sc_hd__nor2_1 _39002_ (.A(_11483_),
    .B(_11484_),
    .Y(_11485_));
 sky130_fd_sc_hd__a31o_1 _39003_ (.A1(_08282_),
    .A2(_09662_),
    .A3(_06776_),
    .B1(_09661_),
    .X(_11486_));
 sky130_fd_sc_hd__xor2_1 _39004_ (.A(_11485_),
    .B(_11486_),
    .X(_11487_));
 sky130_fd_sc_hd__o21a_1 _39005_ (.A1(_09666_),
    .A2(_09671_),
    .B1(_11487_),
    .X(_11488_));
 sky130_fd_sc_hd__nor3_1 _39006_ (.A(_09666_),
    .B(_09671_),
    .C(_11487_),
    .Y(_11489_));
 sky130_fd_sc_hd__or2_1 _39007_ (.A(_11488_),
    .B(_11489_),
    .X(_11490_));
 sky130_fd_sc_hd__buf_1 _39008_ (.A(_09636_),
    .X(_11491_));
 sky130_fd_sc_hd__o21a_1 _39009_ (.A1(_08331_),
    .A2(_09620_),
    .B1(_09625_),
    .X(_11492_));
 sky130_fd_sc_hd__buf_1 _39010_ (.A(\delay_line[33][13] ),
    .X(_11494_));
 sky130_fd_sc_hd__nor3_1 _39011_ (.A(_08322_),
    .B(_11494_),
    .C(_08331_),
    .Y(_11495_));
 sky130_fd_sc_hd__buf_1 _39012_ (.A(_02845_),
    .X(_11496_));
 sky130_fd_sc_hd__o21a_1 _39013_ (.A1(_11494_),
    .A2(_08331_),
    .B1(_08321_),
    .X(_11497_));
 sky130_fd_sc_hd__or4_1 _39014_ (.A(_08320_),
    .B(_11495_),
    .C(_11496_),
    .D(_11497_),
    .X(_11498_));
 sky130_fd_sc_hd__o22ai_1 _39015_ (.A1(_11496_),
    .A2(_08320_),
    .B1(_11495_),
    .B2(_11497_),
    .Y(_11499_));
 sky130_fd_sc_hd__and2b_1 _39016_ (.A_N(_11494_),
    .B(net310),
    .X(_11500_));
 sky130_fd_sc_hd__and2b_1 _39017_ (.A_N(net310),
    .B(_11494_),
    .X(_11501_));
 sky130_fd_sc_hd__a211o_1 _39018_ (.A1(_09615_),
    .A2(_09617_),
    .B1(_11500_),
    .C1(_11501_),
    .X(_11502_));
 sky130_fd_sc_hd__o221ai_2 _39019_ (.A1(_09612_),
    .A2(_09614_),
    .B1(_11501_),
    .B2(_11500_),
    .C1(_09617_),
    .Y(_11503_));
 sky130_fd_sc_hd__nand4_1 _39020_ (.A(_11498_),
    .B(_11499_),
    .C(_11502_),
    .D(_11503_),
    .Y(_11505_));
 sky130_fd_sc_hd__a22o_1 _39021_ (.A1(_11498_),
    .A2(_11499_),
    .B1(_11502_),
    .B2(_11503_),
    .X(_11506_));
 sky130_fd_sc_hd__a31o_1 _39022_ (.A1(_09617_),
    .A2(_09611_),
    .A3(_09615_),
    .B1(_09626_),
    .X(_11507_));
 sky130_fd_sc_hd__a21oi_1 _39023_ (.A1(_11505_),
    .A2(_11506_),
    .B1(_11507_),
    .Y(_11508_));
 sky130_fd_sc_hd__nand3_1 _39024_ (.A(_11505_),
    .B(_11506_),
    .C(_11507_),
    .Y(_11509_));
 sky130_fd_sc_hd__or3b_1 _39025_ (.A(_11492_),
    .B(_11508_),
    .C_N(_11509_),
    .X(_11510_));
 sky130_fd_sc_hd__or2b_1 _39026_ (.A(_11508_),
    .B_N(_11509_),
    .X(_11511_));
 sky130_fd_sc_hd__nand2_1 _39027_ (.A(_11511_),
    .B(_11492_),
    .Y(_11512_));
 sky130_fd_sc_hd__nand2_1 _39028_ (.A(_11510_),
    .B(_11512_),
    .Y(_11513_));
 sky130_fd_sc_hd__o311a_1 _39029_ (.A1(_09629_),
    .A2(_09626_),
    .A3(_09627_),
    .B1(_11491_),
    .C1(_11513_),
    .X(_11514_));
 sky130_fd_sc_hd__a21oi_1 _39030_ (.A1(_09631_),
    .A2(_11491_),
    .B1(_11513_),
    .Y(_11516_));
 sky130_fd_sc_hd__nor2_1 _39031_ (.A(_11514_),
    .B(_11516_),
    .Y(_11517_));
 sky130_fd_sc_hd__and4_1 _39032_ (.A(_11517_),
    .B(_09638_),
    .C(_09637_),
    .D(_11491_),
    .X(_11518_));
 sky130_fd_sc_hd__a31o_1 _39033_ (.A1(_11491_),
    .A2(_09637_),
    .A3(_09638_),
    .B1(_11517_),
    .X(_11519_));
 sky130_fd_sc_hd__and2b_1 _39034_ (.A_N(_11518_),
    .B(_11519_),
    .X(_11520_));
 sky130_fd_sc_hd__o21a_1 _39035_ (.A1(_09642_),
    .A2(_09645_),
    .B1(_11520_),
    .X(_11521_));
 sky130_fd_sc_hd__nor3_1 _39036_ (.A(_09642_),
    .B(_09645_),
    .C(_11520_),
    .Y(_11522_));
 sky130_fd_sc_hd__nor2_1 _39037_ (.A(_11521_),
    .B(_11522_),
    .Y(_11523_));
 sky130_fd_sc_hd__buf_1 _39038_ (.A(_06856_),
    .X(_11524_));
 sky130_fd_sc_hd__or2b_1 _39039_ (.A(_09588_),
    .B_N(_11524_),
    .X(_11525_));
 sky130_fd_sc_hd__or2b_1 _39040_ (.A(_06856_),
    .B_N(_09588_),
    .X(_11527_));
 sky130_fd_sc_hd__o2bb2a_1 _39041_ (.A1_N(_11525_),
    .A2_N(_11527_),
    .B1(_01115_),
    .B2(_09586_),
    .X(_11528_));
 sky130_fd_sc_hd__nor2_1 _39042_ (.A(_01115_),
    .B(_09586_),
    .Y(_11529_));
 sky130_fd_sc_hd__and3_1 _39043_ (.A(_11529_),
    .B(_11525_),
    .C(_11527_),
    .X(_11530_));
 sky130_fd_sc_hd__o221a_1 _39044_ (.A1(_11528_),
    .A2(_11530_),
    .B1(_09584_),
    .B2(_09592_),
    .C1(_09583_),
    .X(_11531_));
 sky130_fd_sc_hd__a211oi_1 _39045_ (.A1(_09583_),
    .A2(_09593_),
    .B1(_11528_),
    .C1(_11530_),
    .Y(_11532_));
 sky130_fd_sc_hd__or3_1 _39046_ (.A(_09589_),
    .B(_11531_),
    .C(_11532_),
    .X(_11533_));
 sky130_fd_sc_hd__o21ai_1 _39047_ (.A1(_11531_),
    .A2(_11532_),
    .B1(_09589_),
    .Y(_11534_));
 sky130_fd_sc_hd__a211oi_1 _39048_ (.A1(_11533_),
    .A2(_11534_),
    .B1(_09597_),
    .C1(net155),
    .Y(_11535_));
 sky130_fd_sc_hd__o211a_1 _39049_ (.A1(_09597_),
    .A2(net155),
    .B1(_11533_),
    .C1(_11534_),
    .X(_11536_));
 sky130_fd_sc_hd__or4b_1 _39050_ (.A(_09601_),
    .B(_11535_),
    .C(_11536_),
    .D_N(_09600_),
    .X(_11538_));
 sky130_fd_sc_hd__o32ai_1 _39051_ (.A1(net155),
    .A2(_09599_),
    .A3(_09601_),
    .B1(_11535_),
    .B2(_11536_),
    .Y(_11539_));
 sky130_fd_sc_hd__and2_1 _39052_ (.A(_11538_),
    .B(_11539_),
    .X(_11540_));
 sky130_fd_sc_hd__nor2_1 _39053_ (.A(_08373_),
    .B(_08372_),
    .Y(_11541_));
 sky130_fd_sc_hd__o2bb2ai_1 _39054_ (.A1_N(_11541_),
    .A2_N(_09604_),
    .B1(_09603_),
    .B2(_09606_),
    .Y(_11542_));
 sky130_fd_sc_hd__xor2_1 _39055_ (.A(_11540_),
    .B(_11542_),
    .X(_11543_));
 sky130_fd_sc_hd__nand2_1 _39056_ (.A(_11523_),
    .B(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__or2_1 _39057_ (.A(_11523_),
    .B(_11543_),
    .X(_11545_));
 sky130_fd_sc_hd__and3_1 _39058_ (.A(_11490_),
    .B(_11544_),
    .C(_11545_),
    .X(_11546_));
 sky130_fd_sc_hd__a21oi_1 _39059_ (.A1(_11544_),
    .A2(_11545_),
    .B1(_11490_),
    .Y(_11547_));
 sky130_fd_sc_hd__inv_2 _39060_ (.A(_10232_),
    .Y(_11549_));
 sky130_fd_sc_hd__a32o_2 _39061_ (.A1(_10191_),
    .A2(_10192_),
    .A3(_11549_),
    .B1(_10264_),
    .B2(_10233_),
    .X(_11550_));
 sky130_fd_sc_hd__o21a_1 _39062_ (.A1(_11546_),
    .A2(_11547_),
    .B1(_11550_),
    .X(_11551_));
 sky130_fd_sc_hd__nor3_2 _39063_ (.A(_11547_),
    .B(_11550_),
    .C(_11546_),
    .Y(_11552_));
 sky130_fd_sc_hd__nor2_1 _39064_ (.A(_09649_),
    .B(_09674_),
    .Y(_11553_));
 sky130_fd_sc_hd__o21ai_1 _39065_ (.A1(_11551_),
    .A2(_11552_),
    .B1(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__or3_1 _39066_ (.A(_11553_),
    .B(_11551_),
    .C(_11552_),
    .X(_11555_));
 sky130_fd_sc_hd__a221o_2 _39067_ (.A1(_09574_),
    .A2(_09678_),
    .B1(_11554_),
    .B2(_11555_),
    .C1(_09677_),
    .X(_11556_));
 sky130_fd_sc_hd__a21o_1 _39068_ (.A1(_09574_),
    .A2(_09678_),
    .B1(_09677_),
    .X(_11557_));
 sky130_fd_sc_hd__nand3_2 _39069_ (.A(_11554_),
    .B(_11555_),
    .C(_11557_),
    .Y(_11558_));
 sky130_fd_sc_hd__nand2_1 _39070_ (.A(_09691_),
    .B(net294),
    .Y(_11560_));
 sky130_fd_sc_hd__or2_1 _39071_ (.A(net294),
    .B(_09691_),
    .X(_11561_));
 sky130_fd_sc_hd__nor4_1 _39072_ (.A(_06669_),
    .B(_09691_),
    .C(_09687_),
    .D(_09688_),
    .Y(_11562_));
 sky130_fd_sc_hd__a211o_1 _39073_ (.A1(_11560_),
    .A2(_11561_),
    .B1(net276),
    .C1(_09687_),
    .X(_11563_));
 sky130_fd_sc_hd__o211ai_1 _39074_ (.A1(_09687_),
    .A2(net276),
    .B1(_11561_),
    .C1(_11560_),
    .Y(_11564_));
 sky130_fd_sc_hd__nand2_1 _39075_ (.A(_11563_),
    .B(_11564_),
    .Y(_11565_));
 sky130_fd_sc_hd__a32o_2 _39076_ (.A1(net295),
    .A2(_08240_),
    .A3(_08242_),
    .B1(_09694_),
    .B2(_09695_),
    .X(_11566_));
 sky130_fd_sc_hd__xor2_2 _39077_ (.A(_11565_),
    .B(_11566_),
    .X(_11567_));
 sky130_fd_sc_hd__buf_1 _39078_ (.A(_08249_),
    .X(_11568_));
 sky130_fd_sc_hd__and2b_1 _39079_ (.A_N(_05319_),
    .B(_11568_),
    .X(_11569_));
 sky130_fd_sc_hd__and2b_1 _39080_ (.A_N(_11568_),
    .B(_05319_),
    .X(_11571_));
 sky130_fd_sc_hd__nor2_1 _39081_ (.A(_11569_),
    .B(_11571_),
    .Y(_11572_));
 sky130_fd_sc_hd__o21ba_1 _39082_ (.A1(_03702_),
    .A2(_08253_),
    .B1_N(_09702_),
    .X(_11573_));
 sky130_fd_sc_hd__xnor2_2 _39083_ (.A(_11572_),
    .B(_11573_),
    .Y(_11574_));
 sky130_fd_sc_hd__nor2_1 _39084_ (.A(_09700_),
    .B(_09702_),
    .Y(_11575_));
 sky130_fd_sc_hd__o21ai_1 _39085_ (.A1(_08262_),
    .A2(_08265_),
    .B1(_11575_),
    .Y(_11576_));
 sky130_fd_sc_hd__xnor2_2 _39086_ (.A(_11574_),
    .B(_11576_),
    .Y(_11577_));
 sky130_fd_sc_hd__xnor2_2 _39087_ (.A(_11567_),
    .B(_11577_),
    .Y(_11578_));
 sky130_fd_sc_hd__a211o_1 _39088_ (.A1(_08237_),
    .A2(_08232_),
    .B1(_08231_),
    .C1(_11578_),
    .X(_11579_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39089_ (.A(_09686_),
    .X(_11580_));
 sky130_fd_sc_hd__nand2_1 _39090_ (.A(_11578_),
    .B(_11580_),
    .Y(_11582_));
 sky130_fd_sc_hd__inv_2 _39091_ (.A(_09686_),
    .Y(_11583_));
 sky130_fd_sc_hd__o21ai_1 _39092_ (.A1(_09708_),
    .A2(_11583_),
    .B1(_09707_),
    .Y(_11584_));
 sky130_fd_sc_hd__a21oi_1 _39093_ (.A1(_11579_),
    .A2(_11582_),
    .B1(_11584_),
    .Y(_11585_));
 sky130_fd_sc_hd__o21a_1 _39094_ (.A1(_09716_),
    .A2(_08202_),
    .B1(_09715_),
    .X(_11586_));
 sky130_fd_sc_hd__o21a_1 _39095_ (.A1(_05342_),
    .A2(_08193_),
    .B1(_08192_),
    .X(_11587_));
 sky130_fd_sc_hd__clkbuf_4 _39096_ (.A(_08192_),
    .X(_11588_));
 sky130_fd_sc_hd__o21a_1 _39097_ (.A1(_03663_),
    .A2(_05342_),
    .B1(_11588_),
    .X(_11589_));
 sky130_fd_sc_hd__a2bb2o_1 _39098_ (.A1_N(_06753_),
    .A2_N(_11587_),
    .B1(_11589_),
    .B2(_08193_),
    .X(_11590_));
 sky130_fd_sc_hd__xnor2_1 _39099_ (.A(_11586_),
    .B(_11590_),
    .Y(_11591_));
 sky130_fd_sc_hd__or3_1 _39100_ (.A(_08204_),
    .B(_06717_),
    .C(_05379_),
    .X(_11593_));
 sky130_fd_sc_hd__a21oi_1 _39101_ (.A1(_09721_),
    .A2(_11593_),
    .B1(_09727_),
    .Y(_11594_));
 sky130_fd_sc_hd__or3_1 _39102_ (.A(_05358_),
    .B(_08214_),
    .C(_08215_),
    .X(_11595_));
 sky130_fd_sc_hd__a21oi_2 _39103_ (.A1(_05362_),
    .A2(_11595_),
    .B1(_09733_),
    .Y(_11596_));
 sky130_fd_sc_hd__xnor2_1 _39104_ (.A(_11594_),
    .B(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__or2_1 _39105_ (.A(_11591_),
    .B(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__nand2_1 _39106_ (.A(_11591_),
    .B(_11597_),
    .Y(_11599_));
 sky130_fd_sc_hd__nand2_2 _39107_ (.A(_11598_),
    .B(_11599_),
    .Y(_11600_));
 sky130_fd_sc_hd__nor2_2 _39108_ (.A(_11585_),
    .B(_11600_),
    .Y(_11601_));
 sky130_fd_sc_hd__nand3_1 _39109_ (.A(_11584_),
    .B(_11579_),
    .C(_11582_),
    .Y(_11602_));
 sky130_fd_sc_hd__inv_2 _39110_ (.A(_11602_),
    .Y(_11604_));
 sky130_fd_sc_hd__o21a_1 _39111_ (.A1(_11585_),
    .A2(_11604_),
    .B1(_11600_),
    .X(_11605_));
 sky130_fd_sc_hd__a21o_1 _39112_ (.A1(_11601_),
    .A2(_11602_),
    .B1(_11605_),
    .X(_11606_));
 sky130_fd_sc_hd__a21bo_1 _39113_ (.A1(_11556_),
    .A2(_11558_),
    .B1_N(_11606_),
    .X(_11607_));
 sky130_fd_sc_hd__nand3b_1 _39114_ (.A_N(_11606_),
    .B(_11556_),
    .C(_11558_),
    .Y(_11608_));
 sky130_fd_sc_hd__inv_2 _39115_ (.A(_10127_),
    .Y(_11609_));
 sky130_fd_sc_hd__o21a_1 _39116_ (.A1(_11609_),
    .A2(_10269_),
    .B1(_10271_),
    .X(_11610_));
 sky130_fd_sc_hd__a21bo_1 _39117_ (.A1(_11607_),
    .A2(_11608_),
    .B1_N(_11610_),
    .X(_11611_));
 sky130_fd_sc_hd__nand3b_1 _39118_ (.A_N(_11610_),
    .B(_11607_),
    .C(_11608_),
    .Y(_11612_));
 sky130_fd_sc_hd__nand2_1 _39119_ (.A(_11611_),
    .B(_11612_),
    .Y(_11613_));
 sky130_fd_sc_hd__xor2_1 _39120_ (.A(_11474_),
    .B(_11613_),
    .X(_11615_));
 sky130_fd_sc_hd__or2_1 _39121_ (.A(_11472_),
    .B(_11615_),
    .X(_11616_));
 sky130_fd_sc_hd__nand2_1 _39122_ (.A(_11615_),
    .B(_11472_),
    .Y(_11617_));
 sky130_fd_sc_hd__nand2_1 _39123_ (.A(_11616_),
    .B(_11617_),
    .Y(_11618_));
 sky130_fd_sc_hd__xnor2_2 _39124_ (.A(_10970_),
    .B(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__nand3_1 _39125_ (.A(_10968_),
    .B(_10962_),
    .C(_10967_),
    .Y(_11620_));
 sky130_fd_sc_hd__nand2_1 _39126_ (.A(_11619_),
    .B(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__nor2_1 _39127_ (.A(_09570_),
    .B(_10283_),
    .Y(_11622_));
 sky130_fd_sc_hd__a21o_1 _39128_ (.A1(_10962_),
    .A2(_10967_),
    .B1(_10968_),
    .X(_11623_));
 sky130_fd_sc_hd__clkbuf_2 _39129_ (.A(_11620_),
    .X(_11624_));
 sky130_fd_sc_hd__a21o_1 _39130_ (.A1(_11623_),
    .A2(_11624_),
    .B1(_11619_),
    .X(_11626_));
 sky130_fd_sc_hd__o221ai_2 _39131_ (.A1(_10969_),
    .A2(_11621_),
    .B1(_10285_),
    .B2(_11622_),
    .C1(_11626_),
    .Y(_11627_));
 sky130_fd_sc_hd__clkbuf_2 _39132_ (.A(_11627_),
    .X(_11628_));
 sky130_fd_sc_hd__nor2_2 _39133_ (.A(_10969_),
    .B(_11621_),
    .Y(_11629_));
 sky130_fd_sc_hd__a21oi_1 _39134_ (.A1(_11623_),
    .A2(_11624_),
    .B1(_11619_),
    .Y(_11630_));
 sky130_fd_sc_hd__o22a_1 _39135_ (.A1(_09572_),
    .A2(_10280_),
    .B1(_09570_),
    .B2(_10283_),
    .X(_11631_));
 sky130_fd_sc_hd__o21ai_2 _39136_ (.A1(_11629_),
    .A2(_11630_),
    .B1(_11631_),
    .Y(_11632_));
 sky130_fd_sc_hd__nand3_1 _39137_ (.A(_10484_),
    .B(_11628_),
    .C(_11632_),
    .Y(_11633_));
 sky130_fd_sc_hd__a21o_1 _39138_ (.A1(_10475_),
    .A2(_10478_),
    .B1(_10479_),
    .X(_11634_));
 sky130_fd_sc_hd__o211ai_2 _39139_ (.A1(_10335_),
    .A2(_10482_),
    .B1(_10475_),
    .C1(_10478_),
    .Y(_11635_));
 sky130_fd_sc_hd__a22o_1 _39140_ (.A1(_11634_),
    .A2(_11635_),
    .B1(_11627_),
    .B2(_11632_),
    .X(_11637_));
 sky130_fd_sc_hd__o211ai_2 _39141_ (.A1(_10425_),
    .A2(_10397_),
    .B1(_11633_),
    .C1(_11637_),
    .Y(_11638_));
 sky130_fd_sc_hd__buf_1 _39142_ (.A(_11638_),
    .X(_11639_));
 sky130_fd_sc_hd__o21a_1 _39143_ (.A1(_10396_),
    .A2(_10355_),
    .B1(_10291_),
    .X(_11640_));
 sky130_fd_sc_hd__nand2_1 _39144_ (.A(_11634_),
    .B(_11635_),
    .Y(_11641_));
 sky130_fd_sc_hd__a21o_1 _39145_ (.A1(_11628_),
    .A2(_11632_),
    .B1(_11641_),
    .X(_11642_));
 sky130_fd_sc_hd__o211ai_1 _39146_ (.A1(_10480_),
    .A2(_10483_),
    .B1(_11628_),
    .C1(_11632_),
    .Y(_11643_));
 sky130_fd_sc_hd__nand3_2 _39147_ (.A(_11640_),
    .B(_11642_),
    .C(_11643_),
    .Y(_11644_));
 sky130_fd_sc_hd__o21ai_1 _39148_ (.A1(_10342_),
    .A2(_10351_),
    .B1(_10346_),
    .Y(_11645_));
 sky130_fd_sc_hd__or2_1 _39149_ (.A(_10378_),
    .B(_10380_),
    .X(_11646_));
 sky130_fd_sc_hd__o21bai_4 _39150_ (.A1(_09061_),
    .A2(_10374_),
    .B1_N(_10373_),
    .Y(_11648_));
 sky130_fd_sc_hd__nor2_1 _39151_ (.A(_04574_),
    .B(_23595_),
    .Y(_11649_));
 sky130_fd_sc_hd__o21a_1 _39152_ (.A1(_23593_),
    .A2(_23594_),
    .B1(_03001_),
    .X(_11650_));
 sky130_fd_sc_hd__a211oi_1 _39153_ (.A1(_20958_),
    .A2(_10367_),
    .B1(_11649_),
    .C1(_11650_),
    .Y(_11651_));
 sky130_fd_sc_hd__inv_2 _39154_ (.A(_11651_),
    .Y(_11652_));
 sky130_fd_sc_hd__o211ai_2 _39155_ (.A1(_11649_),
    .A2(_11650_),
    .B1(_20958_),
    .C1(_10367_),
    .Y(_11653_));
 sky130_fd_sc_hd__a32o_1 _39156_ (.A1(_08957_),
    .A2(_10297_),
    .A3(_08971_),
    .B1(_11652_),
    .B2(_11653_),
    .X(_11654_));
 sky130_fd_sc_hd__nand4_1 _39157_ (.A(_11652_),
    .B(_11653_),
    .C(_08961_),
    .D(_08971_),
    .Y(_11655_));
 sky130_fd_sc_hd__and3_1 _39158_ (.A(_11654_),
    .B(_11655_),
    .C(_10369_),
    .X(_11656_));
 sky130_fd_sc_hd__a21oi_1 _39159_ (.A1(_11654_),
    .A2(_11655_),
    .B1(_10369_),
    .Y(_11657_));
 sky130_fd_sc_hd__o211ai_1 _39160_ (.A1(_08986_),
    .A2(net166),
    .B1(_10312_),
    .C1(_10313_),
    .Y(_11659_));
 sky130_fd_sc_hd__or4_1 _39161_ (.A(_10298_),
    .B(_10299_),
    .C(_10314_),
    .D(_10315_),
    .X(_11660_));
 sky130_fd_sc_hd__o211ai_1 _39162_ (.A1(_11656_),
    .A2(_11657_),
    .B1(_11659_),
    .C1(_11660_),
    .Y(_11661_));
 sky130_fd_sc_hd__a211o_1 _39163_ (.A1(_11659_),
    .A2(_11660_),
    .B1(_11656_),
    .C1(_11657_),
    .X(_11662_));
 sky130_fd_sc_hd__and2_1 _39164_ (.A(_11661_),
    .B(_11662_),
    .X(_11663_));
 sky130_fd_sc_hd__xor2_4 _39165_ (.A(_11648_),
    .B(_11663_),
    .X(_11664_));
 sky130_fd_sc_hd__xnor2_2 _39166_ (.A(_11646_),
    .B(_11664_),
    .Y(_11665_));
 sky130_fd_sc_hd__a21oi_2 _39167_ (.A1(_10353_),
    .A2(_11645_),
    .B1(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__o211a_1 _39168_ (.A1(_10347_),
    .A2(_10343_),
    .B1(_10353_),
    .C1(_11665_),
    .X(_11667_));
 sky130_fd_sc_hd__nor2_1 _39169_ (.A(_11666_),
    .B(_11667_),
    .Y(_11668_));
 sky130_fd_sc_hd__xnor2_1 _39170_ (.A(_10386_),
    .B(_11668_),
    .Y(_11670_));
 sky130_fd_sc_hd__a21o_1 _39171_ (.A1(_11639_),
    .A2(_11644_),
    .B1(_11670_),
    .X(_11671_));
 sky130_fd_sc_hd__nand3_1 _39172_ (.A(_11670_),
    .B(_11639_),
    .C(_11644_),
    .Y(_11672_));
 sky130_fd_sc_hd__o21ai_2 _39173_ (.A1(_09077_),
    .A2(_10390_),
    .B1(_10387_),
    .Y(_11673_));
 sky130_fd_sc_hd__a31oi_2 _39174_ (.A1(_10424_),
    .A2(_11671_),
    .A3(_11672_),
    .B1(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__o21ai_2 _39175_ (.A1(_10391_),
    .A2(_10401_),
    .B1(_10358_),
    .Y(_11675_));
 sky130_fd_sc_hd__xor2_1 _39176_ (.A(_10386_),
    .B(_11668_),
    .X(_11676_));
 sky130_fd_sc_hd__nand3_2 _39177_ (.A(_11676_),
    .B(_11638_),
    .C(_11644_),
    .Y(_11677_));
 sky130_fd_sc_hd__a21o_1 _39178_ (.A1(_11639_),
    .A2(_11644_),
    .B1(_11676_),
    .X(_11678_));
 sky130_fd_sc_hd__nand3_4 _39179_ (.A(_11675_),
    .B(_11677_),
    .C(_11678_),
    .Y(_11679_));
 sky130_fd_sc_hd__o21ai_1 _39180_ (.A1(_09111_),
    .A2(_10412_),
    .B1(_10403_),
    .Y(_11681_));
 sky130_fd_sc_hd__nand3_1 _39181_ (.A(_10424_),
    .B(_11671_),
    .C(_11672_),
    .Y(_11682_));
 sky130_fd_sc_hd__inv_2 _39182_ (.A(_11673_),
    .Y(_11683_));
 sky130_fd_sc_hd__a21oi_1 _39183_ (.A1(_11679_),
    .A2(_11682_),
    .B1(_11683_),
    .Y(_11684_));
 sky130_fd_sc_hd__a221oi_2 _39184_ (.A1(_11674_),
    .A2(_11679_),
    .B1(_11681_),
    .B2(_10410_),
    .C1(_11684_),
    .Y(_11685_));
 sky130_fd_sc_hd__nand2_1 _39185_ (.A(_11674_),
    .B(_11679_),
    .Y(_11686_));
 sky130_fd_sc_hd__a21o_1 _39186_ (.A1(_11679_),
    .A2(_11682_),
    .B1(_11683_),
    .X(_11687_));
 sky130_fd_sc_hd__nand2_1 _39187_ (.A(_10410_),
    .B(_11681_),
    .Y(_11688_));
 sky130_fd_sc_hd__a21oi_1 _39188_ (.A1(_11686_),
    .A2(_11687_),
    .B1(_11688_),
    .Y(_11689_));
 sky130_fd_sc_hd__nor2_2 _39189_ (.A(_11685_),
    .B(_11689_),
    .Y(_11690_));
 sky130_fd_sc_hd__and3_1 _39190_ (.A(_09109_),
    .B(_10415_),
    .C(_10420_),
    .X(_11692_));
 sky130_fd_sc_hd__a21oi_1 _39191_ (.A1(_10417_),
    .A2(_10418_),
    .B1(_10419_),
    .Y(_11693_));
 sky130_fd_sc_hd__a21oi_1 _39192_ (.A1(_09107_),
    .A2(_10420_),
    .B1(_11693_),
    .Y(_11694_));
 sky130_fd_sc_hd__a21oi_2 _39193_ (.A1(_10422_),
    .A2(_11692_),
    .B1(_11694_),
    .Y(_11695_));
 sky130_fd_sc_hd__xnor2_4 _39194_ (.A(_11690_),
    .B(_11695_),
    .Y(_00012_));
 sky130_fd_sc_hd__o21ba_1 _39195_ (.A1(_11689_),
    .A2(_11695_),
    .B1_N(_11685_),
    .X(_11696_));
 sky130_fd_sc_hd__o211ai_4 _39196_ (.A1(_10347_),
    .A2(_10343_),
    .B1(_10353_),
    .C1(_11665_),
    .Y(_11697_));
 sky130_fd_sc_hd__nand2_1 _39197_ (.A(_11639_),
    .B(_11677_),
    .Y(_11698_));
 sky130_fd_sc_hd__inv_2 _39198_ (.A(_10960_),
    .Y(_11699_));
 sky130_fd_sc_hd__a311oi_4 _39199_ (.A1(_10485_),
    .A2(_10931_),
    .A3(_10936_),
    .B1(_10953_),
    .C1(_10955_),
    .Y(_11700_));
 sky130_fd_sc_hd__inv_2 _39200_ (.A(_10941_),
    .Y(_11702_));
 sky130_fd_sc_hd__a2bb2o_1 _39201_ (.A1_N(_10918_),
    .A2_N(_10919_),
    .B1(_10916_),
    .B2(_10939_),
    .X(_11703_));
 sky130_fd_sc_hd__o21ai_1 _39202_ (.A1(_08046_),
    .A2(_09455_),
    .B1(_10851_),
    .Y(_11704_));
 sky130_fd_sc_hd__or3_1 _39203_ (.A(_08046_),
    .B(_09455_),
    .C(_10851_),
    .X(_11705_));
 sky130_fd_sc_hd__o21ba_1 _39204_ (.A1(_10780_),
    .A2(_10776_),
    .B1_N(_10777_),
    .X(_11706_));
 sky130_fd_sc_hd__a21boi_1 _39205_ (.A1(_11704_),
    .A2(_11705_),
    .B1_N(_11706_),
    .Y(_11707_));
 sky130_fd_sc_hd__nand3b_1 _39206_ (.A_N(_11706_),
    .B(_11704_),
    .C(_11705_),
    .Y(_11708_));
 sky130_fd_sc_hd__nand2b_1 _39207_ (.A_N(_11707_),
    .B(_11708_),
    .Y(_11709_));
 sky130_fd_sc_hd__xnor2_1 _39208_ (.A(_10853_),
    .B(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__a21oi_1 _39209_ (.A1(_10782_),
    .A2(_10783_),
    .B1(_10770_),
    .Y(_11711_));
 sky130_fd_sc_hd__nor2_1 _39210_ (.A(_11710_),
    .B(_11711_),
    .Y(_11713_));
 sky130_fd_sc_hd__and2_1 _39211_ (.A(_11711_),
    .B(_11710_),
    .X(_11714_));
 sky130_fd_sc_hd__a21o_1 _39212_ (.A1(_09392_),
    .A2(_09390_),
    .B1(_09389_),
    .X(_11715_));
 sky130_fd_sc_hd__a21oi_1 _39213_ (.A1(_10854_),
    .A2(_11715_),
    .B1(_10858_),
    .Y(_11716_));
 sky130_fd_sc_hd__o21ai_1 _39214_ (.A1(_11713_),
    .A2(_11714_),
    .B1(_11716_),
    .Y(_11717_));
 sky130_fd_sc_hd__or3_2 _39215_ (.A(_11716_),
    .B(_11713_),
    .C(_11714_),
    .X(_11718_));
 sky130_fd_sc_hd__o221a_1 _39216_ (.A1(_10858_),
    .A2(_10859_),
    .B1(_09397_),
    .B2(_09425_),
    .C1(_10861_),
    .X(_11719_));
 sky130_fd_sc_hd__or3b_1 _39217_ (.A(_10858_),
    .B(_10859_),
    .C_N(_10862_),
    .X(_11720_));
 sky130_fd_sc_hd__o21ai_1 _39218_ (.A1(_10847_),
    .A2(_11719_),
    .B1(_11720_),
    .Y(_11721_));
 sky130_fd_sc_hd__a21oi_1 _39219_ (.A1(_11717_),
    .A2(_11718_),
    .B1(_11721_),
    .Y(_11722_));
 sky130_fd_sc_hd__and3_1 _39220_ (.A(_11721_),
    .B(_11717_),
    .C(_11718_),
    .X(_11724_));
 sky130_fd_sc_hd__buf_1 _39221_ (.A(_11724_),
    .X(_11725_));
 sky130_fd_sc_hd__or2_1 _39222_ (.A(_11722_),
    .B(_11725_),
    .X(_11726_));
 sky130_fd_sc_hd__a21oi_1 _39223_ (.A1(_10826_),
    .A2(_10830_),
    .B1(_11726_),
    .Y(_11727_));
 sky130_fd_sc_hd__buf_1 _39224_ (.A(_11727_),
    .X(_11728_));
 sky130_fd_sc_hd__and2_1 _39225_ (.A(_09471_),
    .B(_10845_),
    .X(_11729_));
 sky130_fd_sc_hd__a311o_1 _39226_ (.A1(_10826_),
    .A2(_10830_),
    .A3(_11726_),
    .B1(_10864_),
    .C1(_11729_),
    .X(_11730_));
 sky130_fd_sc_hd__o21a_1 _39227_ (.A1(_11728_),
    .A2(_11730_),
    .B1(_10865_),
    .X(_11731_));
 sky130_fd_sc_hd__inv_2 _39228_ (.A(_11727_),
    .Y(_11732_));
 sky130_fd_sc_hd__o211ai_2 _39229_ (.A1(_10825_),
    .A2(_10741_),
    .B1(_11726_),
    .C1(_10830_),
    .Y(_11733_));
 sky130_fd_sc_hd__and3_1 _39230_ (.A(_11732_),
    .B(_11733_),
    .C(_11730_),
    .X(_11735_));
 sky130_fd_sc_hd__a31o_1 _39231_ (.A1(_10498_),
    .A2(_10531_),
    .A3(_10532_),
    .B1(_10535_),
    .X(_11736_));
 sky130_fd_sc_hd__buf_1 _39232_ (.A(_01741_),
    .X(_11737_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39233_ (.A(_09139_),
    .X(_11738_));
 sky130_fd_sc_hd__nand2_1 _39234_ (.A(_11737_),
    .B(_11738_),
    .Y(_11739_));
 sky130_fd_sc_hd__a21oi_1 _39235_ (.A1(_11737_),
    .A2(_10687_),
    .B1(_09124_),
    .Y(_11740_));
 sky130_fd_sc_hd__and3_1 _39236_ (.A(_11737_),
    .B(_09124_),
    .C(_10687_),
    .X(_11741_));
 sky130_fd_sc_hd__nor3_1 _39237_ (.A(_10677_),
    .B(_11740_),
    .C(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__o21a_1 _39238_ (.A1(_11740_),
    .A2(_11741_),
    .B1(_09128_),
    .X(_11743_));
 sky130_fd_sc_hd__o22a_1 _39239_ (.A1(_09141_),
    .A2(_11739_),
    .B1(_11742_),
    .B2(_11743_),
    .X(_11744_));
 sky130_fd_sc_hd__nor4_1 _39240_ (.A(_09141_),
    .B(_11739_),
    .C(_11742_),
    .D(_11743_),
    .Y(_11746_));
 sky130_fd_sc_hd__or2_1 _39241_ (.A(_11744_),
    .B(net190),
    .X(_11747_));
 sky130_fd_sc_hd__clkbuf_2 _39242_ (.A(_09128_),
    .X(_11748_));
 sky130_fd_sc_hd__clkbuf_2 _39243_ (.A(_11748_),
    .X(_11749_));
 sky130_fd_sc_hd__or3b_1 _39244_ (.A(_25339_),
    .B(_01789_),
    .C_N(_11749_),
    .X(_11750_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39245_ (.A(_23974_),
    .X(_11751_));
 sky130_fd_sc_hd__buf_2 _39246_ (.A(_04646_),
    .X(_11752_));
 sky130_fd_sc_hd__clkbuf_2 _39247_ (.A(_10677_),
    .X(_11753_));
 sky130_fd_sc_hd__a21oi_1 _39248_ (.A1(_11751_),
    .A2(_11753_),
    .B1(_03322_),
    .Y(_11754_));
 sky130_fd_sc_hd__a311oi_2 _39249_ (.A1(_01793_),
    .A2(_11749_),
    .A3(_11751_),
    .B1(_11752_),
    .C1(_11754_),
    .Y(_11755_));
 sky130_fd_sc_hd__nand2_1 _39250_ (.A(_11751_),
    .B(_11753_),
    .Y(_11757_));
 sky130_fd_sc_hd__nand2_1 _39251_ (.A(_11757_),
    .B(_03322_),
    .Y(_11758_));
 sky130_fd_sc_hd__o211a_1 _39252_ (.A1(_01793_),
    .A2(_11757_),
    .B1(_11758_),
    .C1(_11752_),
    .X(_11759_));
 sky130_fd_sc_hd__a211o_1 _39253_ (.A1(_10683_),
    .A2(_11750_),
    .B1(_11755_),
    .C1(_11759_),
    .X(_11760_));
 sky130_fd_sc_hd__o211ai_1 _39254_ (.A1(_11755_),
    .A2(_11759_),
    .B1(_10683_),
    .C1(_11750_),
    .Y(_11761_));
 sky130_fd_sc_hd__nand2_1 _39255_ (.A(_11760_),
    .B(_11761_),
    .Y(_11762_));
 sky130_fd_sc_hd__xor2_2 _39256_ (.A(_11747_),
    .B(_11762_),
    .X(_11763_));
 sky130_fd_sc_hd__a2bb2o_1 _39257_ (.A1_N(_10707_),
    .A2_N(_10704_),
    .B1(_09155_),
    .B2(_10710_),
    .X(_11764_));
 sky130_fd_sc_hd__o21ai_2 _39258_ (.A1(_09196_),
    .A2(_10523_),
    .B1(_10529_),
    .Y(_11765_));
 sky130_fd_sc_hd__nand4_2 _39259_ (.A(_06341_),
    .B(_10513_),
    .C(_10515_),
    .D(_09154_),
    .Y(_11766_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39260_ (.A(_06445_),
    .X(_11768_));
 sky130_fd_sc_hd__nor2_1 _39261_ (.A(_11768_),
    .B(_09154_),
    .Y(_11769_));
 sky130_fd_sc_hd__and2_1 _39262_ (.A(_06445_),
    .B(_09153_),
    .X(_11770_));
 sky130_fd_sc_hd__a211o_1 _39263_ (.A1(_10513_),
    .A2(_11766_),
    .B1(_11769_),
    .C1(_11770_),
    .X(_11771_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39264_ (.A(_09154_),
    .X(_11772_));
 sky130_fd_sc_hd__o211ai_2 _39265_ (.A1(_11769_),
    .A2(_11770_),
    .B1(_10513_),
    .C1(_11766_),
    .Y(_11773_));
 sky130_fd_sc_hd__nand4_1 _39266_ (.A(_11771_),
    .B(_11772_),
    .C(_10705_),
    .D(_11773_),
    .Y(_11774_));
 sky130_fd_sc_hd__a22o_1 _39267_ (.A1(_10705_),
    .A2(_11772_),
    .B1(_11773_),
    .B2(_11771_),
    .X(_11775_));
 sky130_fd_sc_hd__and2_1 _39268_ (.A(_11774_),
    .B(_11775_),
    .X(_11776_));
 sky130_fd_sc_hd__xnor2_1 _39269_ (.A(_11765_),
    .B(_11776_),
    .Y(_11777_));
 sky130_fd_sc_hd__or2b_1 _39270_ (.A(_11764_),
    .B_N(_11777_),
    .X(_11779_));
 sky130_fd_sc_hd__or2b_1 _39271_ (.A(_11777_),
    .B_N(_11764_),
    .X(_11780_));
 sky130_fd_sc_hd__nand2_1 _39272_ (.A(_11779_),
    .B(_11780_),
    .Y(_11781_));
 sky130_fd_sc_hd__nand3_1 _39273_ (.A(_10714_),
    .B(_10717_),
    .C(_11781_),
    .Y(_11782_));
 sky130_fd_sc_hd__a21o_1 _39274_ (.A1(_10714_),
    .A2(_10717_),
    .B1(_11781_),
    .X(_11783_));
 sky130_fd_sc_hd__nand2_1 _39275_ (.A(_11782_),
    .B(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__xnor2_2 _39276_ (.A(_11763_),
    .B(_11784_),
    .Y(_11785_));
 sky130_fd_sc_hd__xnor2_2 _39277_ (.A(_11736_),
    .B(_11785_),
    .Y(_11786_));
 sky130_fd_sc_hd__a311oi_4 _39278_ (.A1(_10702_),
    .A2(_10716_),
    .A3(_10717_),
    .B1(_10722_),
    .C1(_11786_),
    .Y(_11787_));
 sky130_fd_sc_hd__and3_1 _39279_ (.A(_10702_),
    .B(_10716_),
    .C(_10717_),
    .X(_11788_));
 sky130_fd_sc_hd__o21a_1 _39280_ (.A1(_11788_),
    .A2(_10722_),
    .B1(_11786_),
    .X(_11790_));
 sky130_fd_sc_hd__a32o_2 _39281_ (.A1(_10538_),
    .A2(_10630_),
    .A3(_10632_),
    .B1(_10638_),
    .B2(_10656_),
    .X(_11791_));
 sky130_fd_sc_hd__a32o_2 _39282_ (.A1(_10539_),
    .A2(_10606_),
    .A3(_10615_),
    .B1(_10622_),
    .B2(_10631_),
    .X(_11792_));
 sky130_fd_sc_hd__and4b_2 _39283_ (.A_N(_04775_),
    .B(_06272_),
    .C(_10608_),
    .D(_04734_),
    .X(_11793_));
 sky130_fd_sc_hd__or2_1 _39284_ (.A(_04771_),
    .B(_10540_),
    .X(_11794_));
 sky130_fd_sc_hd__nand2_1 _39285_ (.A(_04775_),
    .B(_10608_),
    .Y(_11795_));
 sky130_fd_sc_hd__o2bb2a_1 _39286_ (.A1_N(_11794_),
    .A2_N(_11795_),
    .B1(_06266_),
    .B2(_09277_),
    .X(_11796_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39287_ (.A(_03148_),
    .X(_11797_));
 sky130_fd_sc_hd__and4bb_2 _39288_ (.A_N(_11793_),
    .B_N(_11796_),
    .C(_11797_),
    .D(_10541_),
    .X(_11798_));
 sky130_fd_sc_hd__o2bb2a_1 _39289_ (.A1_N(_11797_),
    .A2_N(_10628_),
    .B1(_11793_),
    .B2(_11796_),
    .X(_11799_));
 sky130_fd_sc_hd__clkbuf_2 _39290_ (.A(_07796_),
    .X(_11801_));
 sky130_fd_sc_hd__and3_2 _39291_ (.A(_11801_),
    .B(_10541_),
    .C(_10607_),
    .X(_11802_));
 sky130_fd_sc_hd__nand2_2 _39292_ (.A(_11801_),
    .B(_09278_),
    .Y(_11803_));
 sky130_fd_sc_hd__nand2_1 _39293_ (.A(_10598_),
    .B(_10608_),
    .Y(_11804_));
 sky130_fd_sc_hd__o2bb2a_1 _39294_ (.A1_N(_11803_),
    .A2_N(_11804_),
    .B1(_06272_),
    .B2(_10545_),
    .X(_11805_));
 sky130_fd_sc_hd__clkbuf_2 _39295_ (.A(_10578_),
    .X(_11806_));
 sky130_fd_sc_hd__inv_2 _39296_ (.A(_10554_),
    .Y(_11807_));
 sky130_fd_sc_hd__nand2_1 _39297_ (.A(_09243_),
    .B(_09244_),
    .Y(_11808_));
 sky130_fd_sc_hd__o211ai_4 _39298_ (.A1(_09237_),
    .A2(_09240_),
    .B1(_11807_),
    .C1(_11808_),
    .Y(_11809_));
 sky130_fd_sc_hd__o2bb2a_2 _39299_ (.A1_N(_10549_),
    .A2_N(_10552_),
    .B1(_10554_),
    .B2(_10559_),
    .X(_11810_));
 sky130_fd_sc_hd__or2_1 _39300_ (.A(_10549_),
    .B(_10556_),
    .X(_11812_));
 sky130_fd_sc_hd__nand2_1 _39301_ (.A(_10557_),
    .B(_10549_),
    .Y(_11813_));
 sky130_fd_sc_hd__a31oi_2 _39302_ (.A1(_10551_),
    .A2(_07767_),
    .A3(\delay_line[4][14] ),
    .B1(_10548_),
    .Y(_11814_));
 sky130_fd_sc_hd__a21oi_2 _39303_ (.A1(_11812_),
    .A2(_11813_),
    .B1(_11814_),
    .Y(_11815_));
 sky130_fd_sc_hd__and3_1 _39304_ (.A(_11814_),
    .B(_11813_),
    .C(_11812_),
    .X(_11816_));
 sky130_fd_sc_hd__or2_1 _39305_ (.A(_11815_),
    .B(_11816_),
    .X(_11817_));
 sky130_fd_sc_hd__a21oi_2 _39306_ (.A1(_11809_),
    .A2(_11810_),
    .B1(_11817_),
    .Y(_11818_));
 sky130_fd_sc_hd__inv_2 _39307_ (.A(_10572_),
    .Y(_11819_));
 sky130_fd_sc_hd__and4b_2 _39308_ (.A_N(_06233_),
    .B(_11819_),
    .C(_09247_),
    .D(net409),
    .X(_11820_));
 sky130_fd_sc_hd__inv_2 _39309_ (.A(_11820_),
    .Y(_11821_));
 sky130_fd_sc_hd__clkbuf_2 _39310_ (.A(\delay_line[11][12] ),
    .X(_11823_));
 sky130_fd_sc_hd__clkbuf_2 _39311_ (.A(net408),
    .X(_11824_));
 sky130_fd_sc_hd__clkbuf_2 _39312_ (.A(\delay_line[11][13] ),
    .X(_11825_));
 sky130_fd_sc_hd__a31oi_4 _39313_ (.A1(_10567_),
    .A2(_11823_),
    .A3(_11824_),
    .B1(_11825_),
    .Y(_11826_));
 sky130_fd_sc_hd__and2_1 _39314_ (.A(_11823_),
    .B(_11825_),
    .X(_11827_));
 sky130_fd_sc_hd__and3_1 _39315_ (.A(_10567_),
    .B(_11824_),
    .C(_11827_),
    .X(_11828_));
 sky130_fd_sc_hd__nor2_1 _39316_ (.A(_11826_),
    .B(_11828_),
    .Y(_11829_));
 sky130_fd_sc_hd__a21oi_1 _39317_ (.A1(_10586_),
    .A2(_11821_),
    .B1(_11829_),
    .Y(_11830_));
 sky130_fd_sc_hd__and3_1 _39318_ (.A(_10586_),
    .B(_11829_),
    .C(_11821_),
    .X(_11831_));
 sky130_fd_sc_hd__o211ai_4 _39319_ (.A1(_11815_),
    .A2(_11816_),
    .B1(_11810_),
    .C1(_11809_),
    .Y(_11832_));
 sky130_fd_sc_hd__o21ai_2 _39320_ (.A1(_11830_),
    .A2(_11831_),
    .B1(_11832_),
    .Y(_11834_));
 sky130_fd_sc_hd__clkbuf_2 _39321_ (.A(_10549_),
    .X(_11835_));
 sky130_fd_sc_hd__a22o_1 _39322_ (.A1(_11835_),
    .A2(_10552_),
    .B1(_11807_),
    .B2(_10561_),
    .X(_11836_));
 sky130_fd_sc_hd__a211oi_4 _39323_ (.A1(_09243_),
    .A2(_09244_),
    .B1(_10555_),
    .C1(_09256_),
    .Y(_11837_));
 sky130_fd_sc_hd__o21ai_1 _39324_ (.A1(_11836_),
    .A2(_11837_),
    .B1(_11817_),
    .Y(_11838_));
 sky130_fd_sc_hd__nand3b_1 _39325_ (.A_N(_11817_),
    .B(_11809_),
    .C(_11810_),
    .Y(_11839_));
 sky130_fd_sc_hd__a311o_1 _39326_ (.A1(_10567_),
    .A2(_11824_),
    .A3(_11827_),
    .B1(_11820_),
    .C1(_11826_),
    .X(_11840_));
 sky130_fd_sc_hd__o22ai_4 _39327_ (.A1(_11826_),
    .A2(_11828_),
    .B1(_11820_),
    .B2(_10576_),
    .Y(_11841_));
 sky130_fd_sc_hd__o21a_1 _39328_ (.A1(_10576_),
    .A2(_11840_),
    .B1(_11841_),
    .X(_11842_));
 sky130_fd_sc_hd__nand3_1 _39329_ (.A(_11838_),
    .B(_11839_),
    .C(_11842_),
    .Y(_11843_));
 sky130_fd_sc_hd__o21ai_1 _39330_ (.A1(_11818_),
    .A2(_11834_),
    .B1(_11843_),
    .Y(_11845_));
 sky130_fd_sc_hd__o21ai_2 _39331_ (.A1(_10594_),
    .A2(_10596_),
    .B1(_11801_),
    .Y(_11846_));
 sky130_fd_sc_hd__nand3_2 _39332_ (.A(_11806_),
    .B(_11845_),
    .C(_11846_),
    .Y(_11847_));
 sky130_fd_sc_hd__a21oi_2 _39333_ (.A1(_10588_),
    .A2(_10562_),
    .B1(_10598_),
    .Y(_11848_));
 sky130_fd_sc_hd__o21ai_4 _39334_ (.A1(_10576_),
    .A2(_11840_),
    .B1(_11841_),
    .Y(_11849_));
 sky130_fd_sc_hd__o21bai_2 _39335_ (.A1(_11836_),
    .A2(_11837_),
    .B1_N(_11817_),
    .Y(_11850_));
 sky130_fd_sc_hd__nand3_2 _39336_ (.A(_11849_),
    .B(_11850_),
    .C(_11832_),
    .Y(_11851_));
 sky130_fd_sc_hd__buf_2 _39337_ (.A(_11843_),
    .X(_11852_));
 sky130_fd_sc_hd__o211ai_4 _39338_ (.A1(_10604_),
    .A2(_11848_),
    .B1(_11851_),
    .C1(_11852_),
    .Y(_11853_));
 sky130_fd_sc_hd__o21ai_1 _39339_ (.A1(_10594_),
    .A2(_10596_),
    .B1(_11806_),
    .Y(_11854_));
 sky130_fd_sc_hd__o2bb2ai_1 _39340_ (.A1_N(_11801_),
    .A2_N(_11854_),
    .B1(_10603_),
    .B2(_10604_),
    .Y(_11856_));
 sky130_fd_sc_hd__a21oi_2 _39341_ (.A1(_11847_),
    .A2(_11853_),
    .B1(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__buf_2 _39342_ (.A(_10598_),
    .X(_11858_));
 sky130_fd_sc_hd__a21oi_1 _39343_ (.A1(_11806_),
    .A2(_10589_),
    .B1(_11858_),
    .Y(_11859_));
 sky130_fd_sc_hd__o211a_1 _39344_ (.A1(_10611_),
    .A2(_11859_),
    .B1(_11853_),
    .C1(_11847_),
    .X(_11860_));
 sky130_fd_sc_hd__o22ai_4 _39345_ (.A1(_11802_),
    .A2(_11805_),
    .B1(_11857_),
    .B2(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__a21o_1 _39346_ (.A1(_11847_),
    .A2(_11853_),
    .B1(_11856_),
    .X(_11862_));
 sky130_fd_sc_hd__o211ai_2 _39347_ (.A1(_10611_),
    .A2(_11859_),
    .B1(_11853_),
    .C1(_11847_),
    .Y(_11863_));
 sky130_fd_sc_hd__nor2_1 _39348_ (.A(_11802_),
    .B(_11805_),
    .Y(_11864_));
 sky130_fd_sc_hd__nand3_2 _39349_ (.A(_11862_),
    .B(_11863_),
    .C(_11864_),
    .Y(_11865_));
 sky130_fd_sc_hd__a21o_1 _39350_ (.A1(_10617_),
    .A2(_10614_),
    .B1(_10601_),
    .X(_11867_));
 sky130_fd_sc_hd__a21oi_2 _39351_ (.A1(_11861_),
    .A2(_11865_),
    .B1(_11867_),
    .Y(_11868_));
 sky130_fd_sc_hd__o211a_1 _39352_ (.A1(_10607_),
    .A2(_09277_),
    .B1(_10609_),
    .C1(_10614_),
    .X(_11869_));
 sky130_fd_sc_hd__o211a_1 _39353_ (.A1(_10601_),
    .A2(_11869_),
    .B1(_11865_),
    .C1(_11861_),
    .X(_11870_));
 sky130_fd_sc_hd__o22ai_4 _39354_ (.A1(_11798_),
    .A2(_11799_),
    .B1(_11868_),
    .B2(_11870_),
    .Y(_11871_));
 sky130_fd_sc_hd__or2_1 _39355_ (.A(_11798_),
    .B(_11799_),
    .X(_11872_));
 sky130_fd_sc_hd__a21o_1 _39356_ (.A1(_11861_),
    .A2(_11865_),
    .B1(_11867_),
    .X(_11873_));
 sky130_fd_sc_hd__o211ai_4 _39357_ (.A1(_10601_),
    .A2(_11869_),
    .B1(_11865_),
    .C1(_11861_),
    .Y(_11874_));
 sky130_fd_sc_hd__nand3b_4 _39358_ (.A_N(_11872_),
    .B(_11873_),
    .C(_11874_),
    .Y(_11875_));
 sky130_fd_sc_hd__nand3_4 _39359_ (.A(_11792_),
    .B(_11871_),
    .C(_11875_),
    .Y(_11876_));
 sky130_fd_sc_hd__o21bai_1 _39360_ (.A1(_11868_),
    .A2(_11870_),
    .B1_N(_11872_),
    .Y(_11878_));
 sky130_fd_sc_hd__a32oi_1 _39361_ (.A1(_10539_),
    .A2(_10606_),
    .A3(_10615_),
    .B1(_10622_),
    .B2(_10631_),
    .Y(_11879_));
 sky130_fd_sc_hd__nand3_1 _39362_ (.A(_11872_),
    .B(_11873_),
    .C(_11874_),
    .Y(_11880_));
 sky130_fd_sc_hd__nand3_1 _39363_ (.A(_11878_),
    .B(_11879_),
    .C(_11880_),
    .Y(_11881_));
 sky130_fd_sc_hd__buf_2 _39364_ (.A(_11881_),
    .X(_11882_));
 sky130_fd_sc_hd__clkbuf_2 _39365_ (.A(_06198_),
    .X(_11883_));
 sky130_fd_sc_hd__nand2_1 _39366_ (.A(_04786_),
    .B(_11883_),
    .Y(_11884_));
 sky130_fd_sc_hd__or2_1 _39367_ (.A(_04786_),
    .B(_11883_),
    .X(_11885_));
 sky130_fd_sc_hd__a211oi_2 _39368_ (.A1(_11884_),
    .A2(_11885_),
    .B1(_10625_),
    .C1(_10627_),
    .Y(_11886_));
 sky130_fd_sc_hd__o211a_2 _39369_ (.A1(_10625_),
    .A2(_10627_),
    .B1(_11884_),
    .C1(_11885_),
    .X(_11887_));
 sky130_fd_sc_hd__nor2_1 _39370_ (.A(_11886_),
    .B(_11887_),
    .Y(_11889_));
 sky130_fd_sc_hd__o211a_2 _39371_ (.A1(_10648_),
    .A2(_10645_),
    .B1(_11889_),
    .C1(_10641_),
    .X(_11890_));
 sky130_fd_sc_hd__nor2_1 _39372_ (.A(_10647_),
    .B(_11889_),
    .Y(_11891_));
 sky130_fd_sc_hd__o2bb2ai_4 _39373_ (.A1_N(_11876_),
    .A2_N(_11882_),
    .B1(_11890_),
    .B2(_11891_),
    .Y(_11892_));
 sky130_fd_sc_hd__nor3_2 _39374_ (.A(_10647_),
    .B(_11886_),
    .C(_11887_),
    .Y(_11893_));
 sky130_fd_sc_hd__o221a_2 _39375_ (.A1(_10648_),
    .A2(_10645_),
    .B1(_11886_),
    .B2(_11887_),
    .C1(_10641_),
    .X(_11894_));
 sky130_fd_sc_hd__o211ai_4 _39376_ (.A1(_11893_),
    .A2(_11894_),
    .B1(_11876_),
    .C1(_11882_),
    .Y(_11895_));
 sky130_fd_sc_hd__nand3_4 _39377_ (.A(_11791_),
    .B(_11892_),
    .C(_11895_),
    .Y(_11896_));
 sky130_fd_sc_hd__o2bb2ai_1 _39378_ (.A1_N(_11876_),
    .A2_N(_11881_),
    .B1(_11893_),
    .B2(_11894_),
    .Y(_11897_));
 sky130_fd_sc_hd__a32oi_2 _39379_ (.A1(_10538_),
    .A2(_10630_),
    .A3(_10632_),
    .B1(_10638_),
    .B2(_10656_),
    .Y(_11898_));
 sky130_fd_sc_hd__o211ai_1 _39380_ (.A1(_11890_),
    .A2(_11891_),
    .B1(_11876_),
    .C1(_11882_),
    .Y(_11900_));
 sky130_fd_sc_hd__nand3_2 _39381_ (.A(_11897_),
    .B(_11898_),
    .C(_11900_),
    .Y(_11901_));
 sky130_fd_sc_hd__buf_2 _39382_ (.A(_11901_),
    .X(_11902_));
 sky130_fd_sc_hd__or2b_1 _39383_ (.A(_10509_),
    .B_N(_10531_),
    .X(_11903_));
 sky130_fd_sc_hd__o211ai_2 _39384_ (.A1(_09222_),
    .A2(_09223_),
    .B1(_01537_),
    .C1(_10651_),
    .Y(_11904_));
 sky130_fd_sc_hd__buf_1 _39385_ (.A(_10507_),
    .X(_11905_));
 sky130_fd_sc_hd__o2111a_1 _39386_ (.A1(_10644_),
    .A2(_10643_),
    .B1(_11905_),
    .C1(_07891_),
    .D1(_09204_),
    .X(_11906_));
 sky130_fd_sc_hd__nor2_1 _39387_ (.A(_01527_),
    .B(_09204_),
    .Y(_11907_));
 sky130_fd_sc_hd__o22a_1 _39388_ (.A1(_10643_),
    .A2(_10644_),
    .B1(_01527_),
    .B2(_10505_),
    .X(_11908_));
 sky130_fd_sc_hd__and3_1 _39389_ (.A(_07888_),
    .B(_09204_),
    .C(_11905_),
    .X(_11909_));
 sky130_fd_sc_hd__o22a_1 _39390_ (.A1(_11907_),
    .A2(_10508_),
    .B1(_11908_),
    .B2(_11909_),
    .X(_11911_));
 sky130_fd_sc_hd__nor2_1 _39391_ (.A(_11906_),
    .B(_11911_),
    .Y(_11912_));
 sky130_fd_sc_hd__or2_1 _39392_ (.A(_25370_),
    .B(_07869_),
    .X(_11913_));
 sky130_fd_sc_hd__nand2_1 _39393_ (.A(_07869_),
    .B(_25376_),
    .Y(_11914_));
 sky130_fd_sc_hd__a22o_1 _39394_ (.A1(_03283_),
    .A2(_07861_),
    .B1(_11913_),
    .B2(_11914_),
    .X(_11915_));
 sky130_fd_sc_hd__nand4_1 _39395_ (.A(_11913_),
    .B(_11914_),
    .C(_03283_),
    .D(_06363_),
    .Y(_11916_));
 sky130_fd_sc_hd__and3_1 _39396_ (.A(_11915_),
    .B(_10511_),
    .C(_11916_),
    .X(_11917_));
 sky130_fd_sc_hd__o2bb2a_1 _39397_ (.A1_N(_11916_),
    .A2_N(_11915_),
    .B1(_04844_),
    .B2(_07878_),
    .X(_11918_));
 sky130_fd_sc_hd__and2b_1 _39398_ (.A_N(_06363_),
    .B(_06364_),
    .X(_11919_));
 sky130_fd_sc_hd__and2b_1 _39399_ (.A_N(_06364_),
    .B(_06363_),
    .X(_11920_));
 sky130_fd_sc_hd__o21ai_1 _39400_ (.A1(_10518_),
    .A2(_10519_),
    .B1(_09202_),
    .Y(_11922_));
 sky130_fd_sc_hd__or3_1 _39401_ (.A(_11919_),
    .B(_11920_),
    .C(_11922_),
    .X(_11923_));
 sky130_fd_sc_hd__o21ai_1 _39402_ (.A1(_11919_),
    .A2(_11920_),
    .B1(_11922_),
    .Y(_11924_));
 sky130_fd_sc_hd__o211a_1 _39403_ (.A1(_11917_),
    .A2(_11918_),
    .B1(_11923_),
    .C1(_11924_),
    .X(_11925_));
 sky130_fd_sc_hd__a211oi_1 _39404_ (.A1(_11923_),
    .A2(_11924_),
    .B1(_11917_),
    .C1(_11918_),
    .Y(_11926_));
 sky130_fd_sc_hd__nor2_1 _39405_ (.A(_11925_),
    .B(_11926_),
    .Y(_11927_));
 sky130_fd_sc_hd__xnor2_1 _39406_ (.A(_11912_),
    .B(_11927_),
    .Y(_11928_));
 sky130_fd_sc_hd__nand3_1 _39407_ (.A(_10650_),
    .B(_11904_),
    .C(_11928_),
    .Y(_11929_));
 sky130_fd_sc_hd__a21o_1 _39408_ (.A1(_10650_),
    .A2(_11904_),
    .B1(_11928_),
    .X(_11930_));
 sky130_fd_sc_hd__nand2_1 _39409_ (.A(_11929_),
    .B(_11930_),
    .Y(_11931_));
 sky130_fd_sc_hd__nor2_1 _39410_ (.A(_11903_),
    .B(_11931_),
    .Y(_11933_));
 sky130_fd_sc_hd__and2_1 _39411_ (.A(_11903_),
    .B(_11931_),
    .X(_11934_));
 sky130_fd_sc_hd__or2_4 _39412_ (.A(_11933_),
    .B(_11934_),
    .X(_11935_));
 sky130_fd_sc_hd__a21oi_4 _39413_ (.A1(_11896_),
    .A2(_11902_),
    .B1(_11935_),
    .Y(_11936_));
 sky130_fd_sc_hd__nand2_1 _39414_ (.A(_10655_),
    .B(_10658_),
    .Y(_11937_));
 sky130_fd_sc_hd__inv_2 _39415_ (.A(_10659_),
    .Y(_11938_));
 sky130_fd_sc_hd__a21oi_2 _39416_ (.A1(_11937_),
    .A2(_11938_),
    .B1(_10665_),
    .Y(_11939_));
 sky130_fd_sc_hd__nand3_4 _39417_ (.A(_11896_),
    .B(_11901_),
    .C(_11935_),
    .Y(_11940_));
 sky130_fd_sc_hd__o21ai_2 _39418_ (.A1(_10663_),
    .A2(_11939_),
    .B1(_11940_),
    .Y(_11941_));
 sky130_fd_sc_hd__nor2_1 _39419_ (.A(_11936_),
    .B(_11941_),
    .Y(_11942_));
 sky130_fd_sc_hd__or2b_1 _39420_ (.A(_11931_),
    .B_N(_11903_),
    .X(_11944_));
 sky130_fd_sc_hd__inv_2 _39421_ (.A(_11944_),
    .Y(_11945_));
 sky130_fd_sc_hd__and3b_1 _39422_ (.A_N(_10509_),
    .B(_10531_),
    .C(_11931_),
    .X(_11946_));
 sky130_fd_sc_hd__o2bb2ai_4 _39423_ (.A1_N(_11896_),
    .A2_N(_11902_),
    .B1(_11945_),
    .B2(_11946_),
    .Y(_11947_));
 sky130_fd_sc_hd__o21ai_2 _39424_ (.A1(_10665_),
    .A2(_10660_),
    .B1(_10667_),
    .Y(_11948_));
 sky130_fd_sc_hd__a21oi_4 _39425_ (.A1(_11940_),
    .A2(_11947_),
    .B1(_11948_),
    .Y(_11949_));
 sky130_fd_sc_hd__o22ai_2 _39426_ (.A1(_11787_),
    .A2(_11790_),
    .B1(_11942_),
    .B2(_11949_),
    .Y(_11950_));
 sky130_fd_sc_hd__a21oi_1 _39427_ (.A1(_10674_),
    .A2(_10730_),
    .B1(_10737_),
    .Y(_11951_));
 sky130_fd_sc_hd__nor2_1 _39428_ (.A(_11787_),
    .B(_11790_),
    .Y(_11952_));
 sky130_fd_sc_hd__o211a_1 _39429_ (.A1(_11933_),
    .A2(_11934_),
    .B1(_11896_),
    .C1(_11902_),
    .X(_11953_));
 sky130_fd_sc_hd__o21bai_2 _39430_ (.A1(_11953_),
    .A2(_11936_),
    .B1_N(_11948_),
    .Y(_11955_));
 sky130_fd_sc_hd__o211ai_2 _39431_ (.A1(_11941_),
    .A2(_11936_),
    .B1(_11952_),
    .C1(_11955_),
    .Y(_11956_));
 sky130_fd_sc_hd__nand3_4 _39432_ (.A(_11950_),
    .B(_11951_),
    .C(_11956_),
    .Y(_11957_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39433_ (.A(_11957_),
    .X(_11958_));
 sky130_fd_sc_hd__o22ai_4 _39434_ (.A1(_11787_),
    .A2(_11790_),
    .B1(_11936_),
    .B2(_11941_),
    .Y(_11959_));
 sky130_fd_sc_hd__a32o_1 _39435_ (.A1(_10496_),
    .A2(_10664_),
    .A3(_10669_),
    .B1(_10674_),
    .B2(_10730_),
    .X(_11960_));
 sky130_fd_sc_hd__o21ba_1 _39436_ (.A1(_11788_),
    .A2(_10722_),
    .B1_N(_11786_),
    .X(_11961_));
 sky130_fd_sc_hd__nor3b_2 _39437_ (.A(_11788_),
    .B(_10722_),
    .C_N(_11786_),
    .Y(_11962_));
 sky130_fd_sc_hd__o22ai_2 _39438_ (.A1(_11961_),
    .A2(_11962_),
    .B1(_11942_),
    .B2(_11949_),
    .Y(_11963_));
 sky130_fd_sc_hd__o211ai_4 _39439_ (.A1(_11959_),
    .A2(_11949_),
    .B1(_11960_),
    .C1(_11963_),
    .Y(_11964_));
 sky130_fd_sc_hd__o21a_1 _39440_ (.A1(_10787_),
    .A2(_10824_),
    .B1(_10821_),
    .X(_11966_));
 sky130_fd_sc_hd__inv_2 _39441_ (.A(_10819_),
    .Y(_11967_));
 sky130_fd_sc_hd__or2b_1 _39442_ (.A(\delay_line[7][14] ),
    .B_N(\delay_line[7][15] ),
    .X(_11968_));
 sky130_fd_sc_hd__or2b_1 _39443_ (.A(\delay_line[7][15] ),
    .B_N(_04659_),
    .X(_11969_));
 sky130_fd_sc_hd__nand2_1 _39444_ (.A(_11968_),
    .B(_11969_),
    .Y(_11970_));
 sky130_fd_sc_hd__nor2_1 _39445_ (.A(_10802_),
    .B(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__and2_1 _39446_ (.A(_11970_),
    .B(_03338_),
    .X(_11972_));
 sky130_fd_sc_hd__or2_1 _39447_ (.A(_25296_),
    .B(_06088_),
    .X(_11973_));
 sky130_fd_sc_hd__nand2_1 _39448_ (.A(_25297_),
    .B(_06088_),
    .Y(_11974_));
 sky130_fd_sc_hd__and4_1 _39449_ (.A(_10806_),
    .B(_10807_),
    .C(_11973_),
    .D(_11974_),
    .X(_11975_));
 sky130_fd_sc_hd__a22oi_4 _39450_ (.A1(_10806_),
    .A2(_10807_),
    .B1(_11973_),
    .B2(_11974_),
    .Y(_11977_));
 sky130_fd_sc_hd__nor4_1 _39451_ (.A(_00268_),
    .B(_09355_),
    .C(_11975_),
    .D(_11977_),
    .Y(_11978_));
 sky130_fd_sc_hd__o22a_1 _39452_ (.A1(_10797_),
    .A2(_00268_),
    .B1(_11977_),
    .B2(_11975_),
    .X(_11979_));
 sky130_fd_sc_hd__nor4_1 _39453_ (.A(_11971_),
    .B(_11972_),
    .C(_11978_),
    .D(_11979_),
    .Y(_11980_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39454_ (.A(_11980_),
    .X(_11981_));
 sky130_fd_sc_hd__o22a_1 _39455_ (.A1(_11971_),
    .A2(_11972_),
    .B1(_11978_),
    .B2(_11979_),
    .X(_11982_));
 sky130_fd_sc_hd__a211oi_1 _39456_ (.A1(_10694_),
    .A2(_10695_),
    .B1(_11981_),
    .C1(_11982_),
    .Y(_11983_));
 sky130_fd_sc_hd__o211a_1 _39457_ (.A1(_11980_),
    .A2(_11982_),
    .B1(_10694_),
    .C1(_10695_),
    .X(_11984_));
 sky130_fd_sc_hd__nor3_1 _39458_ (.A(_11983_),
    .B(_10810_),
    .C(_11984_),
    .Y(_11985_));
 sky130_fd_sc_hd__o21ai_1 _39459_ (.A1(_11984_),
    .A2(_11983_),
    .B1(_10810_),
    .Y(_11986_));
 sky130_fd_sc_hd__and2b_1 _39460_ (.A_N(_11985_),
    .B(_11986_),
    .X(_11988_));
 sky130_fd_sc_hd__o21bai_1 _39461_ (.A1(_10686_),
    .A2(_10697_),
    .B1_N(_10685_),
    .Y(_11989_));
 sky130_fd_sc_hd__nand2_1 _39462_ (.A(_11988_),
    .B(_11989_),
    .Y(_11990_));
 sky130_fd_sc_hd__or2_1 _39463_ (.A(_11989_),
    .B(_11988_),
    .X(_11991_));
 sky130_fd_sc_hd__nand2_1 _39464_ (.A(_11990_),
    .B(_11991_),
    .Y(_11992_));
 sky130_fd_sc_hd__and2b_1 _39465_ (.A_N(_10814_),
    .B(_10816_),
    .X(_11993_));
 sky130_fd_sc_hd__nand2_1 _39466_ (.A(_11992_),
    .B(_11993_),
    .Y(_11994_));
 sky130_fd_sc_hd__or2_1 _39467_ (.A(_11993_),
    .B(_11992_),
    .X(_11995_));
 sky130_fd_sc_hd__nand2_1 _39468_ (.A(_11994_),
    .B(_11995_),
    .Y(_11996_));
 sky130_fd_sc_hd__a21oi_1 _39469_ (.A1(_10817_),
    .A2(_11967_),
    .B1(_11996_),
    .Y(_11997_));
 sky130_fd_sc_hd__nand3_1 _39470_ (.A(_10817_),
    .B(_11967_),
    .C(_11996_),
    .Y(_11999_));
 sky130_fd_sc_hd__inv_2 _39471_ (.A(_11999_),
    .Y(_12000_));
 sky130_fd_sc_hd__a21o_1 _39472_ (.A1(_03457_),
    .A2(_10849_),
    .B1(_10773_),
    .X(_12001_));
 sky130_fd_sc_hd__buf_1 _39473_ (.A(_10746_),
    .X(_12002_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39474_ (.A(_12002_),
    .X(_12003_));
 sky130_fd_sc_hd__a21oi_1 _39475_ (.A1(_12003_),
    .A2(_10749_),
    .B1(_10747_),
    .Y(_12004_));
 sky130_fd_sc_hd__xor2_1 _39476_ (.A(_12001_),
    .B(_12004_),
    .X(_12005_));
 sky130_fd_sc_hd__buf_1 _39477_ (.A(_04933_),
    .X(_12006_));
 sky130_fd_sc_hd__o2bb2a_1 _39478_ (.A1_N(_12006_),
    .A2_N(_10751_),
    .B1(_10753_),
    .B2(_10750_),
    .X(_12007_));
 sky130_fd_sc_hd__or2_2 _39479_ (.A(_12005_),
    .B(_12007_),
    .X(_12008_));
 sky130_fd_sc_hd__nand2_1 _39480_ (.A(_12007_),
    .B(_12005_),
    .Y(_12010_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39481_ (.A(_10746_),
    .X(_12011_));
 sky130_fd_sc_hd__clkbuf_2 _39482_ (.A(_12011_),
    .X(_12012_));
 sky130_fd_sc_hd__clkbuf_2 _39483_ (.A(_10773_),
    .X(_12013_));
 sky130_fd_sc_hd__or2_1 _39484_ (.A(_10849_),
    .B(_12013_),
    .X(_12014_));
 sky130_fd_sc_hd__clkbuf_2 _39485_ (.A(_07996_),
    .X(_12015_));
 sky130_fd_sc_hd__nand2_1 _39486_ (.A(_12015_),
    .B(_10849_),
    .Y(_12016_));
 sky130_fd_sc_hd__a2111oi_1 _39487_ (.A1(_01865_),
    .A2(_04941_),
    .B1(_09400_),
    .C1(_12016_),
    .D1(_09405_),
    .Y(_12017_));
 sky130_fd_sc_hd__a31oi_1 _39488_ (.A1(_12012_),
    .A2(_09402_),
    .A3(_12014_),
    .B1(net245),
    .Y(_12018_));
 sky130_fd_sc_hd__a21boi_1 _39489_ (.A1(_12008_),
    .A2(_12010_),
    .B1_N(_12018_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand3b_2 _39490_ (.A_N(_12018_),
    .B(_12008_),
    .C(_12010_),
    .Y(_12021_));
 sky130_fd_sc_hd__or2b_1 _39491_ (.A(_12019_),
    .B_N(_12021_),
    .X(_12022_));
 sky130_fd_sc_hd__o21ai_1 _39492_ (.A1(_09414_),
    .A2(_09421_),
    .B1(_09420_),
    .Y(_12023_));
 sky130_fd_sc_hd__nor2_1 _39493_ (.A(_10762_),
    .B(_10764_),
    .Y(_12024_));
 sky130_fd_sc_hd__buf_1 _39494_ (.A(_06097_),
    .X(_12025_));
 sky130_fd_sc_hd__buf_1 _39495_ (.A(_10797_),
    .X(_12026_));
 sky130_fd_sc_hd__and3_1 _39496_ (.A(_12025_),
    .B(_09361_),
    .C(_12026_),
    .X(_12027_));
 sky130_fd_sc_hd__a211o_1 _39497_ (.A1(_12025_),
    .A2(_10758_),
    .B1(_10796_),
    .C1(net223),
    .X(_12028_));
 sky130_fd_sc_hd__clkbuf_2 _39498_ (.A(_10758_),
    .X(_12029_));
 sky130_fd_sc_hd__o211ai_2 _39499_ (.A1(_10796_),
    .A2(net223),
    .B1(_12025_),
    .C1(_12029_),
    .Y(_12030_));
 sky130_fd_sc_hd__o211a_1 _39500_ (.A1(_12027_),
    .A2(_10762_),
    .B1(_12028_),
    .C1(_12030_),
    .X(_12032_));
 sky130_fd_sc_hd__buf_1 _39501_ (.A(_04928_),
    .X(_12033_));
 sky130_fd_sc_hd__a21oi_1 _39502_ (.A1(_12006_),
    .A2(_12002_),
    .B1(_12033_),
    .Y(_12034_));
 sky130_fd_sc_hd__and3_1 _39503_ (.A(_12006_),
    .B(_12033_),
    .C(_10746_),
    .X(_12035_));
 sky130_fd_sc_hd__or2_2 _39504_ (.A(_06151_),
    .B(_10773_),
    .X(_12036_));
 sky130_fd_sc_hd__nand2_1 _39505_ (.A(_10773_),
    .B(_06151_),
    .Y(_12037_));
 sky130_fd_sc_hd__nand3_2 _39506_ (.A(_12036_),
    .B(_12002_),
    .C(_12037_),
    .Y(_12038_));
 sky130_fd_sc_hd__a21o_1 _39507_ (.A1(_12037_),
    .A2(_12036_),
    .B1(_10746_),
    .X(_12039_));
 sky130_fd_sc_hd__o211ai_2 _39508_ (.A1(_12034_),
    .A2(_12035_),
    .B1(_12038_),
    .C1(_12039_),
    .Y(_12040_));
 sky130_fd_sc_hd__a211o_1 _39509_ (.A1(_12038_),
    .A2(_12039_),
    .B1(_12034_),
    .C1(_12035_),
    .X(_12041_));
 sky130_fd_sc_hd__nand2_1 _39510_ (.A(_12040_),
    .B(_12041_),
    .Y(_12043_));
 sky130_fd_sc_hd__a221o_1 _39511_ (.A1(_10760_),
    .A2(_10761_),
    .B1(_12028_),
    .B2(_12030_),
    .C1(_12027_),
    .X(_12044_));
 sky130_fd_sc_hd__inv_2 _39512_ (.A(_12044_),
    .Y(_12045_));
 sky130_fd_sc_hd__or3_2 _39513_ (.A(_12032_),
    .B(_12043_),
    .C(_12045_),
    .X(_12046_));
 sky130_fd_sc_hd__o21ai_2 _39514_ (.A1(_12045_),
    .A2(_12032_),
    .B1(_12043_),
    .Y(_12047_));
 sky130_fd_sc_hd__and2b_1 _39515_ (.A_N(_10755_),
    .B(_10768_),
    .X(_12048_));
 sky130_fd_sc_hd__a221o_1 _39516_ (.A1(_12023_),
    .A2(_12024_),
    .B1(_12046_),
    .B2(_12047_),
    .C1(_12048_),
    .X(_12049_));
 sky130_fd_sc_hd__o211ai_4 _39517_ (.A1(_10765_),
    .A2(_12048_),
    .B1(_12047_),
    .C1(_12046_),
    .Y(_12050_));
 sky130_fd_sc_hd__nand2_1 _39518_ (.A(_12049_),
    .B(_12050_),
    .Y(_12051_));
 sky130_fd_sc_hd__xnor2_1 _39519_ (.A(_12022_),
    .B(_12051_),
    .Y(_12052_));
 sky130_fd_sc_hd__o21a_1 _39520_ (.A1(_11997_),
    .A2(_12000_),
    .B1(_12052_),
    .X(_12054_));
 sky130_fd_sc_hd__inv_2 _39521_ (.A(_12054_),
    .Y(_12055_));
 sky130_fd_sc_hd__or3_1 _39522_ (.A(_12052_),
    .B(_11997_),
    .C(_12000_),
    .X(_12056_));
 sky130_fd_sc_hd__a211o_1 _39523_ (.A1(_12055_),
    .A2(_12056_),
    .B1(_10724_),
    .C1(_10727_),
    .X(_12057_));
 sky130_fd_sc_hd__o211ai_2 _39524_ (.A1(_10724_),
    .A2(_10727_),
    .B1(_12055_),
    .C1(_12056_),
    .Y(_12058_));
 sky130_fd_sc_hd__nand2_1 _39525_ (.A(_12057_),
    .B(_12058_),
    .Y(_12059_));
 sky130_fd_sc_hd__xor2_1 _39526_ (.A(_11966_),
    .B(_12059_),
    .X(_12060_));
 sky130_fd_sc_hd__clkbuf_2 _39527_ (.A(_12060_),
    .X(_12061_));
 sky130_fd_sc_hd__a21oi_4 _39528_ (.A1(_11958_),
    .A2(_11964_),
    .B1(_12061_),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_1 _39529_ (.A(_10729_),
    .B(_10731_),
    .Y(_12063_));
 sky130_fd_sc_hd__o21a_1 _39530_ (.A1(_09334_),
    .A2(_09335_),
    .B1(_09328_),
    .X(_12065_));
 sky130_fd_sc_hd__a21oi_1 _39531_ (.A1(_12063_),
    .A2(_12065_),
    .B1(_10832_),
    .Y(_12066_));
 sky130_fd_sc_hd__a31oi_2 _39532_ (.A1(_10671_),
    .A2(_10672_),
    .A3(_10673_),
    .B1(_10735_),
    .Y(_12067_));
 sky130_fd_sc_hd__o22ai_4 _39533_ (.A1(_10737_),
    .A2(_12067_),
    .B1(_11959_),
    .B2(_11949_),
    .Y(_12068_));
 sky130_fd_sc_hd__o211ai_4 _39534_ (.A1(_10663_),
    .A2(_11939_),
    .B1(_11940_),
    .C1(_11947_),
    .Y(_12069_));
 sky130_fd_sc_hd__a2bb2oi_4 _39535_ (.A1_N(_11961_),
    .A2_N(_11962_),
    .B1(_12069_),
    .B2(_11955_),
    .Y(_12070_));
 sky130_fd_sc_hd__o211ai_2 _39536_ (.A1(_12068_),
    .A2(_12070_),
    .B1(_12060_),
    .C1(_11957_),
    .Y(_12071_));
 sky130_fd_sc_hd__o21ai_2 _39537_ (.A1(_10738_),
    .A2(_12066_),
    .B1(_12071_),
    .Y(_12072_));
 sky130_fd_sc_hd__nor2_2 _39538_ (.A(_12062_),
    .B(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__o21ai_1 _39539_ (.A1(_12070_),
    .A2(_12068_),
    .B1(_11958_),
    .Y(_12074_));
 sky130_fd_sc_hd__inv_2 _39540_ (.A(_12061_),
    .Y(_12076_));
 sky130_fd_sc_hd__nand2_1 _39541_ (.A(_12074_),
    .B(_12076_),
    .Y(_12077_));
 sky130_fd_sc_hd__o21ai_1 _39542_ (.A1(_10832_),
    .A2(_10733_),
    .B1(_10836_),
    .Y(_12078_));
 sky130_fd_sc_hd__a21oi_2 _39543_ (.A1(_12077_),
    .A2(_12071_),
    .B1(_12078_),
    .Y(_12079_));
 sky130_fd_sc_hd__o22ai_1 _39544_ (.A1(_11731_),
    .A2(_11735_),
    .B1(_12073_),
    .B2(_12079_),
    .Y(_12080_));
 sky130_fd_sc_hd__a32oi_2 _39545_ (.A1(_10494_),
    .A2(_10834_),
    .A3(_10837_),
    .B1(_10885_),
    .B2(_10876_),
    .Y(_12081_));
 sky130_fd_sc_hd__and3_1 _39546_ (.A(_11732_),
    .B(_11733_),
    .C(_10865_),
    .X(_12082_));
 sky130_fd_sc_hd__a21oi_2 _39547_ (.A1(_11732_),
    .A2(_11733_),
    .B1(_10865_),
    .Y(_12083_));
 sky130_fd_sc_hd__and3_1 _39548_ (.A(_11958_),
    .B(_11964_),
    .C(_12061_),
    .X(_12084_));
 sky130_fd_sc_hd__o21bai_2 _39549_ (.A1(_12062_),
    .A2(_12084_),
    .B1_N(_12078_),
    .Y(_12085_));
 sky130_fd_sc_hd__o221ai_2 _39550_ (.A1(_12082_),
    .A2(_12083_),
    .B1(_12062_),
    .B2(_12072_),
    .C1(_12085_),
    .Y(_12087_));
 sky130_fd_sc_hd__nand3_2 _39551_ (.A(_12080_),
    .B(_12081_),
    .C(_12087_),
    .Y(_12088_));
 sky130_fd_sc_hd__a32o_1 _39552_ (.A1(_10494_),
    .A2(_10834_),
    .A3(_10837_),
    .B1(_10885_),
    .B2(_10876_),
    .X(_12089_));
 sky130_fd_sc_hd__o22ai_2 _39553_ (.A1(_12082_),
    .A2(_12083_),
    .B1(_12073_),
    .B2(_12079_),
    .Y(_12090_));
 sky130_fd_sc_hd__inv_2 _39554_ (.A(_11730_),
    .Y(_12091_));
 sky130_fd_sc_hd__a21o_1 _39555_ (.A1(_12091_),
    .A2(_11732_),
    .B1(_12083_),
    .X(_12092_));
 sky130_fd_sc_hd__inv_2 _39556_ (.A(_12092_),
    .Y(_12093_));
 sky130_fd_sc_hd__o211ai_2 _39557_ (.A1(_12072_),
    .A2(_12062_),
    .B1(_12093_),
    .C1(_12085_),
    .Y(_12094_));
 sky130_fd_sc_hd__nand3_2 _39558_ (.A(_12089_),
    .B(_12090_),
    .C(_12094_),
    .Y(_12095_));
 sky130_fd_sc_hd__a21oi_2 _39559_ (.A1(_10870_),
    .A2(_10869_),
    .B1(_10872_),
    .Y(_12096_));
 sky130_fd_sc_hd__nand3_1 _39560_ (.A(_12088_),
    .B(_12095_),
    .C(_12096_),
    .Y(_12098_));
 sky130_fd_sc_hd__clkbuf_2 _39561_ (.A(_12098_),
    .X(_12099_));
 sky130_fd_sc_hd__o21ai_2 _39562_ (.A1(_09477_),
    .A2(net89),
    .B1(_10889_),
    .Y(_12100_));
 sky130_fd_sc_hd__nand2_1 _39563_ (.A(_12088_),
    .B(_12095_),
    .Y(_12101_));
 sky130_fd_sc_hd__inv_2 _39564_ (.A(_12096_),
    .Y(_12102_));
 sky130_fd_sc_hd__a22oi_4 _39565_ (.A1(_10896_),
    .A2(_12100_),
    .B1(_12101_),
    .B2(_12102_),
    .Y(_12103_));
 sky130_fd_sc_hd__o21a_1 _39566_ (.A1(_09453_),
    .A2(_09475_),
    .B1(_10869_),
    .X(_12104_));
 sky130_fd_sc_hd__o2bb2ai_2 _39567_ (.A1_N(_12088_),
    .A2_N(_12095_),
    .B1(_12104_),
    .B2(_10872_),
    .Y(_12105_));
 sky130_fd_sc_hd__nand2_1 _39568_ (.A(_10896_),
    .B(_12100_),
    .Y(_12106_));
 sky130_fd_sc_hd__a21oi_2 _39569_ (.A1(_12098_),
    .A2(_12105_),
    .B1(_12106_),
    .Y(_12107_));
 sky130_fd_sc_hd__a21oi_4 _39570_ (.A1(_12099_),
    .A2(_12103_),
    .B1(_12107_),
    .Y(_12109_));
 sky130_fd_sc_hd__o211a_1 _39571_ (.A1(_10905_),
    .A2(_10900_),
    .B1(_09489_),
    .C1(_09501_),
    .X(_12110_));
 sky130_fd_sc_hd__nand2_1 _39572_ (.A(_08114_),
    .B(_09507_),
    .Y(_12111_));
 sky130_fd_sc_hd__a22oi_4 _39573_ (.A1(_09505_),
    .A2(_12111_),
    .B1(_08127_),
    .B2(_10908_),
    .Y(_12112_));
 sky130_fd_sc_hd__o22ai_4 _39574_ (.A1(_10898_),
    .A2(_10905_),
    .B1(_12110_),
    .B2(_12112_),
    .Y(_12113_));
 sky130_fd_sc_hd__o21a_2 _39575_ (.A1(_11594_),
    .A2(_11596_),
    .B1(_11598_),
    .X(_12114_));
 sky130_fd_sc_hd__inv_2 _39576_ (.A(_12114_),
    .Y(_12115_));
 sky130_fd_sc_hd__a21o_1 _39577_ (.A1(_10889_),
    .A2(_10896_),
    .B1(_10894_),
    .X(_12116_));
 sky130_fd_sc_hd__a31oi_2 _39578_ (.A1(_10894_),
    .A2(_10889_),
    .A3(_10893_),
    .B1(_10897_),
    .Y(_12117_));
 sky130_fd_sc_hd__a21o_1 _39579_ (.A1(_12116_),
    .A2(_12117_),
    .B1(_12109_),
    .X(_12118_));
 sky130_fd_sc_hd__o21bai_2 _39580_ (.A1(_10906_),
    .A2(_12112_),
    .B1_N(_12118_),
    .Y(_12120_));
 sky130_fd_sc_hd__nand2_1 _39581_ (.A(_12115_),
    .B(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__a21oi_4 _39582_ (.A1(_12109_),
    .A2(_12113_),
    .B1(_12121_),
    .Y(_12122_));
 sky130_fd_sc_hd__nand2_1 _39583_ (.A(_12113_),
    .B(_12109_),
    .Y(_12123_));
 sky130_fd_sc_hd__a21oi_2 _39584_ (.A1(_12120_),
    .A2(_12123_),
    .B1(_12115_),
    .Y(_12124_));
 sky130_fd_sc_hd__o21bai_4 _39585_ (.A1(_12122_),
    .A2(_12124_),
    .B1_N(_10939_),
    .Y(_12125_));
 sky130_fd_sc_hd__a21o_1 _39586_ (.A1(_12120_),
    .A2(_12123_),
    .B1(_12115_),
    .X(_12126_));
 sky130_fd_sc_hd__clkbuf_2 _39587_ (.A(_09521_),
    .X(_12127_));
 sky130_fd_sc_hd__a21o_1 _39588_ (.A1(_12109_),
    .A2(_12113_),
    .B1(_12121_),
    .X(_12128_));
 sky130_fd_sc_hd__nand3_2 _39589_ (.A(_12126_),
    .B(_12127_),
    .C(_12128_),
    .Y(_12129_));
 sky130_fd_sc_hd__a31o_1 _39590_ (.A1(_11584_),
    .A2(_11579_),
    .A3(_11582_),
    .B1(_11601_),
    .X(_12131_));
 sky130_fd_sc_hd__a21o_1 _39591_ (.A1(_12125_),
    .A2(_12129_),
    .B1(_12131_),
    .X(_12132_));
 sky130_fd_sc_hd__o211ai_4 _39592_ (.A1(_11604_),
    .A2(_11601_),
    .B1(_12125_),
    .C1(_12129_),
    .Y(_12133_));
 sky130_fd_sc_hd__nand3_1 _39593_ (.A(_11703_),
    .B(_12132_),
    .C(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__a21oi_2 _39594_ (.A1(_12125_),
    .A2(_12129_),
    .B1(_12131_),
    .Y(_12135_));
 sky130_fd_sc_hd__o211a_1 _39595_ (.A1(_11604_),
    .A2(_11601_),
    .B1(_12125_),
    .C1(_12129_),
    .X(_12136_));
 sky130_fd_sc_hd__inv_2 _39596_ (.A(_11703_),
    .Y(_12137_));
 sky130_fd_sc_hd__o21ai_1 _39597_ (.A1(_12135_),
    .A2(_12136_),
    .B1(_12137_),
    .Y(_12138_));
 sky130_fd_sc_hd__o211ai_2 _39598_ (.A1(_10938_),
    .A2(_11702_),
    .B1(_12134_),
    .C1(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__o21ai_1 _39599_ (.A1(_12135_),
    .A2(_12136_),
    .B1(_11703_),
    .Y(_12140_));
 sky130_fd_sc_hd__o31a_1 _39600_ (.A1(_10924_),
    .A2(_10928_),
    .A3(_10929_),
    .B1(_10941_),
    .X(_12142_));
 sky130_fd_sc_hd__nand3_1 _39601_ (.A(_12132_),
    .B(_12133_),
    .C(_12137_),
    .Y(_12143_));
 sky130_fd_sc_hd__nand3_2 _39602_ (.A(_12140_),
    .B(_12142_),
    .C(_12143_),
    .Y(_12144_));
 sky130_fd_sc_hd__nand2_1 _39603_ (.A(_12139_),
    .B(_12144_),
    .Y(_12145_));
 sky130_fd_sc_hd__nor2_1 _39604_ (.A(_24252_),
    .B(_02015_),
    .Y(_12146_));
 sky130_fd_sc_hd__nand2_2 _39605_ (.A(_24252_),
    .B(_02019_),
    .Y(_12147_));
 sky130_fd_sc_hd__and2b_1 _39606_ (.A_N(_12146_),
    .B(_12147_),
    .X(_12148_));
 sky130_fd_sc_hd__and3_1 _39607_ (.A(_24238_),
    .B(_06644_),
    .C(_24251_),
    .X(_12149_));
 sky130_fd_sc_hd__o21ba_1 _39608_ (.A1(_24256_),
    .A2(_12148_),
    .B1_N(_12149_),
    .X(_12150_));
 sky130_fd_sc_hd__clkbuf_2 _39609_ (.A(_08132_),
    .X(_12151_));
 sky130_fd_sc_hd__clkbuf_2 _39610_ (.A(_08163_),
    .X(_12153_));
 sky130_fd_sc_hd__and3_1 _39611_ (.A(_12151_),
    .B(_09526_),
    .C(_12153_),
    .X(_12154_));
 sky130_fd_sc_hd__nand2_2 _39612_ (.A(_12151_),
    .B(_10933_),
    .Y(_12155_));
 sky130_fd_sc_hd__or3_1 _39613_ (.A(_08163_),
    .B(_08132_),
    .C(_10933_),
    .X(_12156_));
 sky130_fd_sc_hd__and3b_1 _39614_ (.A_N(_12154_),
    .B(_12155_),
    .C(_12156_),
    .X(_12157_));
 sky130_fd_sc_hd__xor2_2 _39615_ (.A(_12150_),
    .B(_12157_),
    .X(_12158_));
 sky130_fd_sc_hd__nand2_1 _39616_ (.A(_12145_),
    .B(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__inv_2 _39617_ (.A(_12158_),
    .Y(_12160_));
 sky130_fd_sc_hd__nand3_2 _39618_ (.A(_12139_),
    .B(_12144_),
    .C(_12160_),
    .Y(_12161_));
 sky130_fd_sc_hd__a21boi_4 _39619_ (.A1(_11611_),
    .A2(_11474_),
    .B1_N(_11612_),
    .Y(_12162_));
 sky130_fd_sc_hd__nand3_2 _39620_ (.A(_12159_),
    .B(_12161_),
    .C(_12162_),
    .Y(_12164_));
 sky130_fd_sc_hd__nand2_1 _39621_ (.A(_12144_),
    .B(_12158_),
    .Y(_12165_));
 sky130_fd_sc_hd__o211a_1 _39622_ (.A1(_10938_),
    .A2(_11702_),
    .B1(_12134_),
    .C1(_12138_),
    .X(_12166_));
 sky130_fd_sc_hd__inv_2 _39623_ (.A(_12162_),
    .Y(_12167_));
 sky130_fd_sc_hd__nand2_1 _39624_ (.A(_12145_),
    .B(_12160_),
    .Y(_12168_));
 sky130_fd_sc_hd__o211ai_4 _39625_ (.A1(_12165_),
    .A2(_12166_),
    .B1(_12167_),
    .C1(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__o211a_1 _39626_ (.A1(_11699_),
    .A2(_11700_),
    .B1(_12164_),
    .C1(_12169_),
    .X(_12170_));
 sky130_fd_sc_hd__a21oi_2 _39627_ (.A1(_10959_),
    .A2(_10956_),
    .B1(_11699_),
    .Y(_12171_));
 sky130_fd_sc_hd__a21boi_1 _39628_ (.A1(_12164_),
    .A2(_12169_),
    .B1_N(_12171_),
    .Y(_12172_));
 sky130_fd_sc_hd__a32o_1 _39629_ (.A1(_11320_),
    .A2(_11313_),
    .A3(_11316_),
    .B1(_11321_),
    .B2(_11466_),
    .X(_12173_));
 sky130_fd_sc_hd__a21boi_1 _39630_ (.A1(_11194_),
    .A2(_11192_),
    .B1_N(_11191_),
    .Y(_12175_));
 sky130_fd_sc_hd__o21ai_1 _39631_ (.A1(_09796_),
    .A2(_09832_),
    .B1(_11004_),
    .Y(_12176_));
 sky130_fd_sc_hd__o21bai_2 _39632_ (.A1(_09836_),
    .A2(_09839_),
    .B1_N(_12176_),
    .Y(_12177_));
 sky130_fd_sc_hd__o2bb2a_1 _39633_ (.A1_N(_10999_),
    .A2_N(_10975_),
    .B1(_10974_),
    .B2(_11000_),
    .X(_12178_));
 sky130_fd_sc_hd__clkbuf_2 _39634_ (.A(_09797_),
    .X(_12179_));
 sky130_fd_sc_hd__and3_1 _39635_ (.A(_07425_),
    .B(_12179_),
    .C(_05698_),
    .X(_12180_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39636_ (.A(_05698_),
    .X(_12181_));
 sky130_fd_sc_hd__clkbuf_2 _39637_ (.A(_07418_),
    .X(_12182_));
 sky130_fd_sc_hd__nand2_2 _39638_ (.A(_12182_),
    .B(_09797_),
    .Y(_12183_));
 sky130_fd_sc_hd__or2_1 _39639_ (.A(_07418_),
    .B(_09797_),
    .X(_12184_));
 sky130_fd_sc_hd__a22oi_2 _39640_ (.A1(_12181_),
    .A2(_12179_),
    .B1(_12183_),
    .B2(_12184_),
    .Y(_12186_));
 sky130_fd_sc_hd__or3b_1 _39641_ (.A(_04047_),
    .B(_05691_),
    .C_N(_09803_),
    .X(_12187_));
 sky130_fd_sc_hd__nor2_2 _39642_ (.A(_04047_),
    .B(_05691_),
    .Y(_12188_));
 sky130_fd_sc_hd__or2_1 _39643_ (.A(_09803_),
    .B(_12188_),
    .X(_12189_));
 sky130_fd_sc_hd__o21ai_1 _39644_ (.A1(_10980_),
    .A2(_10979_),
    .B1(_05697_),
    .Y(_12190_));
 sky130_fd_sc_hd__a21oi_1 _39645_ (.A1(_12187_),
    .A2(_12189_),
    .B1(_12190_),
    .Y(_12191_));
 sky130_fd_sc_hd__and3_1 _39646_ (.A(_12187_),
    .B(_12189_),
    .C(_12190_),
    .X(_12192_));
 sky130_fd_sc_hd__o22a_1 _39647_ (.A1(_12180_),
    .A2(_12186_),
    .B1(_12191_),
    .B2(_12192_),
    .X(_12193_));
 sky130_fd_sc_hd__nor4_1 _39648_ (.A(_12180_),
    .B(_12186_),
    .C(_12191_),
    .D(_12192_),
    .Y(_12194_));
 sky130_fd_sc_hd__o211a_1 _39649_ (.A1(_12193_),
    .A2(_12194_),
    .B1(_10985_),
    .C1(_10988_),
    .X(_12195_));
 sky130_fd_sc_hd__a211o_1 _39650_ (.A1(_10985_),
    .A2(_10988_),
    .B1(_12193_),
    .C1(_12194_),
    .X(_12197_));
 sky130_fd_sc_hd__inv_2 _39651_ (.A(_12197_),
    .Y(_12198_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39652_ (.A(_09803_),
    .X(_12199_));
 sky130_fd_sc_hd__a21o_1 _39653_ (.A1(_07427_),
    .A2(_12199_),
    .B1(_07423_),
    .X(_12200_));
 sky130_fd_sc_hd__o21ai_1 _39654_ (.A1(_10979_),
    .A2(_02589_),
    .B1(_10977_),
    .Y(_12201_));
 sky130_fd_sc_hd__nand2_1 _39655_ (.A(_12200_),
    .B(_12201_),
    .Y(_12202_));
 sky130_fd_sc_hd__o21ai_1 _39656_ (.A1(_12195_),
    .A2(_12198_),
    .B1(_12202_),
    .Y(_12203_));
 sky130_fd_sc_hd__or3_1 _39657_ (.A(_12202_),
    .B(_12195_),
    .C(_12198_),
    .X(_12204_));
 sky130_fd_sc_hd__a211oi_1 _39658_ (.A1(_12203_),
    .A2(_12204_),
    .B1(_10992_),
    .C1(_10996_),
    .Y(_12205_));
 sky130_fd_sc_hd__o211ai_2 _39659_ (.A1(_10992_),
    .A2(_10996_),
    .B1(_12203_),
    .C1(_12204_),
    .Y(_12206_));
 sky130_fd_sc_hd__or2b_1 _39660_ (.A(_12205_),
    .B_N(_12206_),
    .X(_12208_));
 sky130_fd_sc_hd__a211o_1 _39661_ (.A1(_22944_),
    .A2(_10980_),
    .B1(_10973_),
    .C1(_09807_),
    .X(_12209_));
 sky130_fd_sc_hd__xor2_1 _39662_ (.A(_12208_),
    .B(_12209_),
    .X(_12210_));
 sky130_fd_sc_hd__and2b_1 _39663_ (.A_N(_12178_),
    .B(_12210_),
    .X(_12211_));
 sky130_fd_sc_hd__and2b_1 _39664_ (.A_N(_12210_),
    .B(_12178_),
    .X(_12212_));
 sky130_fd_sc_hd__nor2_1 _39665_ (.A(_12211_),
    .B(_12212_),
    .Y(_12213_));
 sky130_fd_sc_hd__a21oi_1 _39666_ (.A1(_11002_),
    .A2(_12177_),
    .B1(_12213_),
    .Y(_12214_));
 sky130_fd_sc_hd__o311a_1 _39667_ (.A1(_09834_),
    .A2(_09840_),
    .A3(_11003_),
    .B1(_12213_),
    .C1(_11002_),
    .X(_12215_));
 sky130_fd_sc_hd__nor2_1 _39668_ (.A(_12214_),
    .B(_12215_),
    .Y(_12216_));
 sky130_fd_sc_hd__o21a_1 _39669_ (.A1(_11008_),
    .A2(_11032_),
    .B1(_11033_),
    .X(_12217_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39670_ (.A(_11012_),
    .X(_12219_));
 sky130_fd_sc_hd__and3_1 _39671_ (.A(_11012_),
    .B(_09755_),
    .C(_09753_),
    .X(_12220_));
 sky130_fd_sc_hd__and4bb_1 _39672_ (.A_N(_12220_),
    .B_N(_11027_),
    .C(_11028_),
    .D(_09755_),
    .X(_12221_));
 sky130_fd_sc_hd__clkbuf_2 _39673_ (.A(_08695_),
    .X(_12222_));
 sky130_fd_sc_hd__o21ai_4 _39674_ (.A1(_12222_),
    .A2(_11013_),
    .B1(_11011_),
    .Y(_12223_));
 sky130_fd_sc_hd__clkbuf_2 _39675_ (.A(_11024_),
    .X(_12224_));
 sky130_fd_sc_hd__buf_1 _39676_ (.A(_11016_),
    .X(_12225_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39677_ (.A(_09761_),
    .X(_12226_));
 sky130_fd_sc_hd__buf_1 _39678_ (.A(_02638_),
    .X(_12227_));
 sky130_fd_sc_hd__buf_1 _39679_ (.A(_02635_),
    .X(_12228_));
 sky130_fd_sc_hd__o21a_1 _39680_ (.A1(_11011_),
    .A2(_12227_),
    .B1(_12228_),
    .X(_12230_));
 sky130_fd_sc_hd__nor3_1 _39681_ (.A(_11011_),
    .B(_12228_),
    .C(_12227_),
    .Y(_12231_));
 sky130_fd_sc_hd__buf_1 _39682_ (.A(_07381_),
    .X(_12232_));
 sky130_fd_sc_hd__or3b_2 _39683_ (.A(_12232_),
    .B(_12226_),
    .C_N(_11016_),
    .X(_12233_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39684_ (.A(_09758_),
    .X(_12234_));
 sky130_fd_sc_hd__nor2_1 _39685_ (.A(_12232_),
    .B(_12234_),
    .Y(_12235_));
 sky130_fd_sc_hd__inv_2 _39686_ (.A(_07381_),
    .Y(_12236_));
 sky130_fd_sc_hd__nor2_1 _39687_ (.A(_12236_),
    .B(_12226_),
    .Y(_12237_));
 sky130_fd_sc_hd__a2bb2o_1 _39688_ (.A1_N(_12235_),
    .A2_N(_12237_),
    .B1(_11016_),
    .B2(_12234_),
    .X(_12238_));
 sky130_fd_sc_hd__o211ai_2 _39689_ (.A1(_12230_),
    .A2(_12231_),
    .B1(_12233_),
    .C1(_12238_),
    .Y(_12239_));
 sky130_fd_sc_hd__a211o_1 _39690_ (.A1(_12233_),
    .A2(_12238_),
    .B1(_12230_),
    .C1(_12231_),
    .X(_12241_));
 sky130_fd_sc_hd__nand2_1 _39691_ (.A(_12239_),
    .B(_12241_),
    .Y(_12242_));
 sky130_fd_sc_hd__o311a_1 _39692_ (.A1(_12224_),
    .A2(_12225_),
    .A3(_12226_),
    .B1(_11023_),
    .C1(_12242_),
    .X(_12243_));
 sky130_fd_sc_hd__a21o_1 _39693_ (.A1(_11025_),
    .A2(_11023_),
    .B1(_12242_),
    .X(_12244_));
 sky130_fd_sc_hd__and2b_1 _39694_ (.A_N(_12243_),
    .B(_12244_),
    .X(_12245_));
 sky130_fd_sc_hd__xnor2_2 _39695_ (.A(_12223_),
    .B(_12245_),
    .Y(_12246_));
 sky130_fd_sc_hd__or3_1 _39696_ (.A(_11027_),
    .B(_12221_),
    .C(_12246_),
    .X(_12247_));
 sky130_fd_sc_hd__o21ai_2 _39697_ (.A1(_11027_),
    .A2(_12221_),
    .B1(_12246_),
    .Y(_12248_));
 sky130_fd_sc_hd__a32o_1 _39698_ (.A1(_09753_),
    .A2(_09755_),
    .A3(_12219_),
    .B1(_12247_),
    .B2(_12248_),
    .X(_12249_));
 sky130_fd_sc_hd__o211ai_2 _39699_ (.A1(_11027_),
    .A2(_12246_),
    .B1(_12220_),
    .C1(_12248_),
    .Y(_12250_));
 sky130_fd_sc_hd__and3b_1 _39700_ (.A_N(_12217_),
    .B(_12249_),
    .C(_12250_),
    .X(_12252_));
 sky130_fd_sc_hd__a21boi_1 _39701_ (.A1(_12249_),
    .A2(_12250_),
    .B1_N(_12217_),
    .Y(_12253_));
 sky130_fd_sc_hd__or2_1 _39702_ (.A(_12252_),
    .B(_12253_),
    .X(_12254_));
 sky130_fd_sc_hd__a21oi_1 _39703_ (.A1(_11036_),
    .A2(_11043_),
    .B1(_12254_),
    .Y(_12255_));
 sky130_fd_sc_hd__nand3_1 _39704_ (.A(_11036_),
    .B(_11043_),
    .C(_12254_),
    .Y(_12256_));
 sky130_fd_sc_hd__and2b_1 _39705_ (.A_N(_12255_),
    .B(_12256_),
    .X(_12257_));
 sky130_fd_sc_hd__a21boi_1 _39706_ (.A1(_11079_),
    .A2(_11077_),
    .B1_N(_11078_),
    .Y(_12258_));
 sky130_fd_sc_hd__or3b_1 _39707_ (.A(_04099_),
    .B(_07350_),
    .C_N(_02550_),
    .X(_12259_));
 sky130_fd_sc_hd__nor2_1 _39708_ (.A(_04099_),
    .B(_07350_),
    .Y(_12260_));
 sky130_fd_sc_hd__or2_1 _39709_ (.A(_09849_),
    .B(_12260_),
    .X(_12261_));
 sky130_fd_sc_hd__nand2_1 _39710_ (.A(_12259_),
    .B(_12261_),
    .Y(_12263_));
 sky130_fd_sc_hd__a21oi_1 _39711_ (.A1(_11059_),
    .A2(_11061_),
    .B1(_11058_),
    .Y(_12264_));
 sky130_fd_sc_hd__xor2_1 _39712_ (.A(_12263_),
    .B(_12264_),
    .X(_12265_));
 sky130_fd_sc_hd__or2_1 _39713_ (.A(_05602_),
    .B(_05603_),
    .X(_12266_));
 sky130_fd_sc_hd__mux2_1 _39714_ (.A0(_07336_),
    .A1(_12266_),
    .S(_09845_),
    .X(_12267_));
 sky130_fd_sc_hd__or2_1 _39715_ (.A(_12265_),
    .B(_12267_),
    .X(_12268_));
 sky130_fd_sc_hd__nand2_1 _39716_ (.A(_12265_),
    .B(_12267_),
    .Y(_12269_));
 sky130_fd_sc_hd__a211oi_1 _39717_ (.A1(_12268_),
    .A2(_12269_),
    .B1(_11051_),
    .C1(_11066_),
    .Y(_12270_));
 sky130_fd_sc_hd__o211ai_2 _39718_ (.A1(_11051_),
    .A2(_11066_),
    .B1(_12268_),
    .C1(_12269_),
    .Y(_12271_));
 sky130_fd_sc_hd__inv_2 _39719_ (.A(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__a21o_1 _39720_ (.A1(_09865_),
    .A2(_09849_),
    .B1(_11069_),
    .X(_12274_));
 sky130_fd_sc_hd__o21ai_1 _39721_ (.A1(_11057_),
    .A2(_11058_),
    .B1(_11056_),
    .Y(_12275_));
 sky130_fd_sc_hd__nand2_1 _39722_ (.A(_12274_),
    .B(_12275_),
    .Y(_12276_));
 sky130_fd_sc_hd__o21ai_1 _39723_ (.A1(_12270_),
    .A2(_12272_),
    .B1(_12276_),
    .Y(_12277_));
 sky130_fd_sc_hd__or3_2 _39724_ (.A(_12276_),
    .B(_12270_),
    .C(_12272_),
    .X(_12278_));
 sky130_fd_sc_hd__a211oi_1 _39725_ (.A1(_12277_),
    .A2(_12278_),
    .B1(_11068_),
    .C1(_11074_),
    .Y(_12279_));
 sky130_fd_sc_hd__o211ai_2 _39726_ (.A1(_11068_),
    .A2(_11074_),
    .B1(_12277_),
    .C1(_12278_),
    .Y(_12280_));
 sky130_fd_sc_hd__or2b_1 _39727_ (.A(_12279_),
    .B_N(_12280_),
    .X(_12281_));
 sky130_fd_sc_hd__o221a_1 _39728_ (.A1(_09867_),
    .A2(_11069_),
    .B1(_00614_),
    .B2(_09853_),
    .C1(_09865_),
    .X(_12282_));
 sky130_fd_sc_hd__xnor2_1 _39729_ (.A(_12281_),
    .B(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__and2b_1 _39730_ (.A_N(_12258_),
    .B(_12283_),
    .X(_12285_));
 sky130_fd_sc_hd__and2b_1 _39731_ (.A_N(_12283_),
    .B(_12258_),
    .X(_12286_));
 sky130_fd_sc_hd__nor2_1 _39732_ (.A(_12285_),
    .B(_12286_),
    .Y(_12287_));
 sky130_fd_sc_hd__a31o_1 _39733_ (.A1(_09871_),
    .A2(_09873_),
    .A3(_09876_),
    .B1(_09881_),
    .X(_12288_));
 sky130_fd_sc_hd__a21oi_1 _39734_ (.A1(_12288_),
    .A2(_11082_),
    .B1(_09885_),
    .Y(_12289_));
 sky130_fd_sc_hd__o21ai_2 _39735_ (.A1(_09887_),
    .A2(_09889_),
    .B1(_12289_),
    .Y(_12290_));
 sky130_fd_sc_hd__o311a_1 _39736_ (.A1(_09879_),
    .A2(_09881_),
    .A3(_11082_),
    .B1(_12287_),
    .C1(_12290_),
    .X(_12291_));
 sky130_fd_sc_hd__a21oi_1 _39737_ (.A1(_11083_),
    .A2(_12290_),
    .B1(_12287_),
    .Y(_12292_));
 sky130_fd_sc_hd__nor2_1 _39738_ (.A(_12291_),
    .B(_12292_),
    .Y(_12293_));
 sky130_fd_sc_hd__o21ai_2 _39739_ (.A1(_12216_),
    .A2(_12257_),
    .B1(_12293_),
    .Y(_12294_));
 sky130_fd_sc_hd__a21o_1 _39740_ (.A1(_12216_),
    .A2(_12257_),
    .B1(_12294_),
    .X(_12296_));
 sky130_fd_sc_hd__or3b_4 _39741_ (.A(_12214_),
    .B(_12215_),
    .C_N(_12257_),
    .X(_12297_));
 sky130_fd_sc_hd__or2_1 _39742_ (.A(_12216_),
    .B(_12257_),
    .X(_12298_));
 sky130_fd_sc_hd__a21o_1 _39743_ (.A1(_12297_),
    .A2(_12298_),
    .B1(_12293_),
    .X(_12299_));
 sky130_fd_sc_hd__nor2_1 _39744_ (.A(_11188_),
    .B(_11189_),
    .Y(_12300_));
 sky130_fd_sc_hd__a32o_1 _39745_ (.A1(_11092_),
    .A2(_11116_),
    .A3(_11117_),
    .B1(_11120_),
    .B2(_09955_),
    .X(_12301_));
 sky130_fd_sc_hd__o21a_1 _39746_ (.A1(_07210_),
    .A2(_09962_),
    .B1(_05739_),
    .X(_12302_));
 sky130_fd_sc_hd__o211a_1 _39747_ (.A1(_11093_),
    .A2(_11096_),
    .B1(_05754_),
    .C1(_09969_),
    .X(_12303_));
 sky130_fd_sc_hd__nor2_1 _39748_ (.A(_12302_),
    .B(_12303_),
    .Y(_12304_));
 sky130_fd_sc_hd__a21oi_1 _39749_ (.A1(_11096_),
    .A2(_07214_),
    .B1(_09970_),
    .Y(_12305_));
 sky130_fd_sc_hd__o21a_1 _39750_ (.A1(_05747_),
    .A2(_07214_),
    .B1(_03885_),
    .X(_12307_));
 sky130_fd_sc_hd__o2bb2a_1 _39751_ (.A1_N(_09970_),
    .A2_N(_09958_),
    .B1(_12305_),
    .B2(_12307_),
    .X(_12308_));
 sky130_fd_sc_hd__o31a_1 _39752_ (.A1(_09958_),
    .A2(_11099_),
    .A3(_11100_),
    .B1(_12308_),
    .X(_12309_));
 sky130_fd_sc_hd__a31o_1 _39753_ (.A1(_09970_),
    .A2(_11110_),
    .A3(_11099_),
    .B1(_12309_),
    .X(_12310_));
 sky130_fd_sc_hd__buf_1 _39754_ (.A(_08539_),
    .X(_12311_));
 sky130_fd_sc_hd__o31a_1 _39755_ (.A1(_12311_),
    .A2(_09966_),
    .A3(_11103_),
    .B1(_11109_),
    .X(_12312_));
 sky130_fd_sc_hd__xor2_1 _39756_ (.A(_12310_),
    .B(_12312_),
    .X(_12313_));
 sky130_fd_sc_hd__xnor2_1 _39757_ (.A(_12304_),
    .B(_12313_),
    .Y(_12314_));
 sky130_fd_sc_hd__a21o_1 _39758_ (.A1(_11113_),
    .A2(_11116_),
    .B1(_12314_),
    .X(_12315_));
 sky130_fd_sc_hd__inv_2 _39759_ (.A(_12315_),
    .Y(_12316_));
 sky130_fd_sc_hd__o311a_1 _39760_ (.A1(_11094_),
    .A2(_11095_),
    .A3(_11114_),
    .B1(_12314_),
    .C1(_11113_),
    .X(_12318_));
 sky130_fd_sc_hd__nor2_1 _39761_ (.A(_12316_),
    .B(_12318_),
    .Y(_12319_));
 sky130_fd_sc_hd__xor2_1 _39762_ (.A(_11094_),
    .B(_12319_),
    .X(_12320_));
 sky130_fd_sc_hd__xnor2_1 _39763_ (.A(_12301_),
    .B(_12320_),
    .Y(_12321_));
 sky130_fd_sc_hd__a21oi_1 _39764_ (.A1(_11091_),
    .A2(_11126_),
    .B1(_11124_),
    .Y(_12322_));
 sky130_fd_sc_hd__xnor2_1 _39765_ (.A(_12321_),
    .B(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39766_ (.A(_08597_),
    .X(_12324_));
 sky130_fd_sc_hd__o21ai_2 _39767_ (.A1(_12324_),
    .A2(_24740_),
    .B1(_11131_),
    .Y(_12325_));
 sky130_fd_sc_hd__o21a_1 _39768_ (.A1(_02430_),
    .A2(_02435_),
    .B1(_08597_),
    .X(_12326_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39769_ (.A(_07254_),
    .X(_12327_));
 sky130_fd_sc_hd__nor2_1 _39770_ (.A(_12324_),
    .B(_12327_),
    .Y(_12329_));
 sky130_fd_sc_hd__o21ai_2 _39771_ (.A1(_12326_),
    .A2(_12329_),
    .B1(_08601_),
    .Y(_12330_));
 sky130_fd_sc_hd__or3_1 _39772_ (.A(_08601_),
    .B(_12326_),
    .C(_12329_),
    .X(_12331_));
 sky130_fd_sc_hd__a2111oi_1 _39773_ (.A1(_09930_),
    .A2(_11135_),
    .B1(_11133_),
    .C1(_11134_),
    .D1(_11136_),
    .Y(_12332_));
 sky130_fd_sc_hd__a221oi_2 _39774_ (.A1(_08606_),
    .A2(_09928_),
    .B1(_12330_),
    .B2(_12331_),
    .C1(net218),
    .Y(_12333_));
 sky130_fd_sc_hd__o211ai_2 _39775_ (.A1(_11134_),
    .A2(net219),
    .B1(_12330_),
    .C1(_12331_),
    .Y(_12334_));
 sky130_fd_sc_hd__and2b_1 _39776_ (.A_N(_12333_),
    .B(_12334_),
    .X(_12335_));
 sky130_fd_sc_hd__xnor2_2 _39777_ (.A(_12325_),
    .B(_12335_),
    .Y(_12336_));
 sky130_fd_sc_hd__o21ai_2 _39778_ (.A1(_11144_),
    .A2(_11143_),
    .B1(_12336_),
    .Y(_12337_));
 sky130_fd_sc_hd__or3_1 _39779_ (.A(_11144_),
    .B(_11143_),
    .C(_12336_),
    .X(_12338_));
 sky130_fd_sc_hd__a21o_1 _39780_ (.A1(_12337_),
    .A2(_12338_),
    .B1(_11132_),
    .X(_12340_));
 sky130_fd_sc_hd__o211ai_1 _39781_ (.A1(_11144_),
    .A2(_12336_),
    .B1(_11132_),
    .C1(_12337_),
    .Y(_12341_));
 sky130_fd_sc_hd__a211o_1 _39782_ (.A1(_12340_),
    .A2(_12341_),
    .B1(_11146_),
    .C1(_11148_),
    .X(_12342_));
 sky130_fd_sc_hd__o211ai_1 _39783_ (.A1(_11146_),
    .A2(_11148_),
    .B1(_12340_),
    .C1(_12341_),
    .Y(_12343_));
 sky130_fd_sc_hd__and2_1 _39784_ (.A(_12342_),
    .B(_12343_),
    .X(_12344_));
 sky130_fd_sc_hd__inv_2 _39785_ (.A(_12344_),
    .Y(_12345_));
 sky130_fd_sc_hd__a21o_1 _39786_ (.A1(_11151_),
    .A2(_11156_),
    .B1(_12345_),
    .X(_12346_));
 sky130_fd_sc_hd__nand3_1 _39787_ (.A(_11151_),
    .B(_11156_),
    .C(_12345_),
    .Y(_12347_));
 sky130_fd_sc_hd__and3_1 _39788_ (.A(_11176_),
    .B(_11177_),
    .C(_11179_),
    .X(_12348_));
 sky130_fd_sc_hd__xnor2_1 _39789_ (.A(_11162_),
    .B(_07293_),
    .Y(_12349_));
 sky130_fd_sc_hd__xnor2_1 _39790_ (.A(_07293_),
    .B(net389),
    .Y(_12351_));
 sky130_fd_sc_hd__and3_1 _39791_ (.A(_12349_),
    .B(_12351_),
    .C(\delay_line[14][15] ),
    .X(_12352_));
 sky130_fd_sc_hd__a21oi_1 _39792_ (.A1(_12349_),
    .A2(net388),
    .B1(_12351_),
    .Y(_12353_));
 sky130_fd_sc_hd__a21o_1 _39793_ (.A1(_11162_),
    .A2(_11164_),
    .B1(_08570_),
    .X(_12354_));
 sky130_fd_sc_hd__nand3_2 _39794_ (.A(_08570_),
    .B(_11162_),
    .C(_11164_),
    .Y(_12355_));
 sky130_fd_sc_hd__o211a_1 _39795_ (.A1(_12352_),
    .A2(_12353_),
    .B1(_12354_),
    .C1(_12355_),
    .X(_12356_));
 sky130_fd_sc_hd__a211o_1 _39796_ (.A1(_12354_),
    .A2(_12355_),
    .B1(_12352_),
    .C1(_12353_),
    .X(_12357_));
 sky130_fd_sc_hd__and2b_1 _39797_ (.A_N(_12356_),
    .B(_12357_),
    .X(_12358_));
 sky130_fd_sc_hd__o211a_1 _39798_ (.A1(_11166_),
    .A2(_11167_),
    .B1(_11169_),
    .C1(_11170_),
    .X(_12359_));
 sky130_fd_sc_hd__a31o_1 _39799_ (.A1(_11160_),
    .A2(_11159_),
    .A3(_12349_),
    .B1(_12359_),
    .X(_12360_));
 sky130_fd_sc_hd__nand2_1 _39800_ (.A(_12358_),
    .B(_12360_),
    .Y(_12362_));
 sky130_fd_sc_hd__a311o_1 _39801_ (.A1(_11160_),
    .A2(_11159_),
    .A3(_12349_),
    .B1(_12359_),
    .C1(_12358_),
    .X(_12363_));
 sky130_fd_sc_hd__a32o_1 _39802_ (.A1(_08568_),
    .A2(_11158_),
    .A3(_11168_),
    .B1(_12362_),
    .B2(_12363_),
    .X(_12364_));
 sky130_fd_sc_hd__nand4_1 _39803_ (.A(_12363_),
    .B(_11168_),
    .C(_11158_),
    .D(_08568_),
    .Y(_12365_));
 sky130_fd_sc_hd__nand2_1 _39804_ (.A(_12364_),
    .B(_12365_),
    .Y(_12366_));
 sky130_fd_sc_hd__a21oi_1 _39805_ (.A1(_11173_),
    .A2(_11177_),
    .B1(_12366_),
    .Y(_12367_));
 sky130_fd_sc_hd__and3_1 _39806_ (.A(_11173_),
    .B(_11177_),
    .C(_12366_),
    .X(_12368_));
 sky130_fd_sc_hd__or2_1 _39807_ (.A(_12367_),
    .B(_12368_),
    .X(_12369_));
 sky130_fd_sc_hd__o21ba_1 _39808_ (.A1(_12348_),
    .A2(_11184_),
    .B1_N(_12369_),
    .X(_12370_));
 sky130_fd_sc_hd__or3b_1 _39809_ (.A(_12348_),
    .B(_11184_),
    .C_N(_12369_),
    .X(_12371_));
 sky130_fd_sc_hd__nand2b_4 _39810_ (.A_N(_12370_),
    .B(_12371_),
    .Y(_12373_));
 sky130_fd_sc_hd__a21o_1 _39811_ (.A1(_12346_),
    .A2(_12347_),
    .B1(_12373_),
    .X(_12374_));
 sky130_fd_sc_hd__nand3_1 _39812_ (.A(_12373_),
    .B(_12346_),
    .C(_12347_),
    .Y(_12375_));
 sky130_fd_sc_hd__and3_1 _39813_ (.A(_12323_),
    .B(_12374_),
    .C(_12375_),
    .X(_12376_));
 sky130_fd_sc_hd__nand2_1 _39814_ (.A(_12346_),
    .B(_12347_),
    .Y(_12377_));
 sky130_fd_sc_hd__a21o_1 _39815_ (.A1(_12377_),
    .A2(_12373_),
    .B1(_12323_),
    .X(_12378_));
 sky130_fd_sc_hd__o21ba_1 _39816_ (.A1(_12373_),
    .A2(_12377_),
    .B1_N(_12378_),
    .X(_12379_));
 sky130_fd_sc_hd__or3_4 _39817_ (.A(_12300_),
    .B(_12376_),
    .C(_12379_),
    .X(_12380_));
 sky130_fd_sc_hd__o21ai_4 _39818_ (.A1(_12376_),
    .A2(_12379_),
    .B1(_12300_),
    .Y(_12381_));
 sky130_fd_sc_hd__nand4_4 _39819_ (.A(_12296_),
    .B(_12299_),
    .C(_12380_),
    .D(_12381_),
    .Y(_12382_));
 sky130_fd_sc_hd__a22o_2 _39820_ (.A1(_12296_),
    .A2(_12299_),
    .B1(_12380_),
    .B2(_12381_),
    .X(_12384_));
 sky130_fd_sc_hd__nand3b_4 _39821_ (.A_N(_12175_),
    .B(_12382_),
    .C(_12384_),
    .Y(_12385_));
 sky130_fd_sc_hd__inv_2 _39822_ (.A(_12385_),
    .Y(_12386_));
 sky130_fd_sc_hd__inv_2 _39823_ (.A(_11301_),
    .Y(_12387_));
 sky130_fd_sc_hd__o21a_1 _39824_ (.A1(_11266_),
    .A2(_12387_),
    .B1(_11304_),
    .X(_12388_));
 sky130_fd_sc_hd__nand2_4 _39825_ (.A(_11045_),
    .B(_11089_),
    .Y(_12389_));
 sky130_fd_sc_hd__or3_1 _39826_ (.A(_11219_),
    .B(_11202_),
    .C(_08406_),
    .X(_12390_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39827_ (.A(_11204_),
    .X(_12391_));
 sky130_fd_sc_hd__o21ai_1 _39828_ (.A1(_12391_),
    .A2(_11202_),
    .B1(_11219_),
    .Y(_12392_));
 sky130_fd_sc_hd__nand3b_2 _39829_ (.A_N(_10010_),
    .B(_05867_),
    .C(_07088_),
    .Y(_12393_));
 sky130_fd_sc_hd__nand3b_1 _39830_ (.A_N(_07088_),
    .B(_11204_),
    .C(_10010_),
    .Y(_12395_));
 sky130_fd_sc_hd__o211a_1 _39831_ (.A1(_11204_),
    .A2(_11205_),
    .B1(_12393_),
    .C1(_12395_),
    .X(_12396_));
 sky130_fd_sc_hd__and3_1 _39832_ (.A(_08418_),
    .B(_08414_),
    .C(_12396_),
    .X(_12397_));
 sky130_fd_sc_hd__a21oi_1 _39833_ (.A1(_08418_),
    .A2(_08414_),
    .B1(_12396_),
    .Y(_12398_));
 sky130_fd_sc_hd__o211a_1 _39834_ (.A1(_12397_),
    .A2(_12398_),
    .B1(_11210_),
    .C1(_11212_),
    .X(_12399_));
 sky130_fd_sc_hd__a211o_1 _39835_ (.A1(_11210_),
    .A2(_11212_),
    .B1(_12397_),
    .C1(_12398_),
    .X(_12400_));
 sky130_fd_sc_hd__and2b_1 _39836_ (.A_N(_12399_),
    .B(_12400_),
    .X(_12401_));
 sky130_fd_sc_hd__xnor2_1 _39837_ (.A(_12392_),
    .B(_12401_),
    .Y(_12402_));
 sky130_fd_sc_hd__a311o_1 _39838_ (.A1(_11216_),
    .A2(_10005_),
    .A3(_12390_),
    .B1(_12402_),
    .C1(_11215_),
    .X(_12403_));
 sky130_fd_sc_hd__and3_1 _39839_ (.A(_10005_),
    .B(_11217_),
    .C(_12390_),
    .X(_12404_));
 sky130_fd_sc_hd__o21a_1 _39840_ (.A1(_11215_),
    .A2(_12404_),
    .B1(_12402_),
    .X(_12406_));
 sky130_fd_sc_hd__nor2_1 _39841_ (.A(_12390_),
    .B(_12406_),
    .Y(_12407_));
 sky130_fd_sc_hd__or2b_1 _39842_ (.A(_12406_),
    .B_N(_12403_),
    .X(_12408_));
 sky130_fd_sc_hd__a22o_1 _39843_ (.A1(_12403_),
    .A2(_12407_),
    .B1(_12408_),
    .B2(_12390_),
    .X(_12409_));
 sky130_fd_sc_hd__a41o_1 _39844_ (.A1(_11202_),
    .A2(_11224_),
    .A3(_08402_),
    .A4(_08408_),
    .B1(_11223_),
    .X(_12410_));
 sky130_fd_sc_hd__and2b_1 _39845_ (.A_N(_12409_),
    .B(_12410_),
    .X(_12411_));
 sky130_fd_sc_hd__and2b_1 _39846_ (.A_N(_12410_),
    .B(_12409_),
    .X(_12412_));
 sky130_fd_sc_hd__nor2_1 _39847_ (.A(_12411_),
    .B(_12412_),
    .Y(_12413_));
 sky130_fd_sc_hd__a21oi_1 _39848_ (.A1(_10000_),
    .A2(_10028_),
    .B1(_11200_),
    .Y(_12414_));
 sky130_fd_sc_hd__o21ai_1 _39849_ (.A1(_11226_),
    .A2(_12414_),
    .B1(_11227_),
    .Y(_12415_));
 sky130_fd_sc_hd__xnor2_1 _39850_ (.A(_12413_),
    .B(_12415_),
    .Y(_12417_));
 sky130_fd_sc_hd__nand2_1 _39851_ (.A(_11294_),
    .B(_11296_),
    .Y(_12418_));
 sky130_fd_sc_hd__clkbuf_2 _39852_ (.A(_10074_),
    .X(_12419_));
 sky130_fd_sc_hd__buf_1 _39853_ (.A(_11268_),
    .X(_12420_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39854_ (.A(_12420_),
    .X(_12421_));
 sky130_fd_sc_hd__nor2_1 _39855_ (.A(_07166_),
    .B(_10080_),
    .Y(_12422_));
 sky130_fd_sc_hd__o211a_1 _39856_ (.A1(_11268_),
    .A2(_07164_),
    .B1(_07166_),
    .C1(_10074_),
    .X(_12423_));
 sky130_fd_sc_hd__nor2_1 _39857_ (.A(_12422_),
    .B(_12423_),
    .Y(_12424_));
 sky130_fd_sc_hd__buf_1 _39858_ (.A(_08488_),
    .X(_12425_));
 sky130_fd_sc_hd__a21oi_1 _39859_ (.A1(_07164_),
    .A2(_07159_),
    .B1(_10087_),
    .Y(_12426_));
 sky130_fd_sc_hd__o21a_1 _39860_ (.A1(_05948_),
    .A2(_07159_),
    .B1(_10087_),
    .X(_12428_));
 sky130_fd_sc_hd__o2bb2a_1 _39861_ (.A1_N(_11268_),
    .A2_N(_12425_),
    .B1(_12426_),
    .B2(_12428_),
    .X(_12429_));
 sky130_fd_sc_hd__o31a_1 _39862_ (.A1(_12425_),
    .A2(_11274_),
    .A3(_11275_),
    .B1(_12429_),
    .X(_12430_));
 sky130_fd_sc_hd__a31o_1 _39863_ (.A1(_11268_),
    .A2(_12425_),
    .A3(_11274_),
    .B1(_12430_),
    .X(_12431_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39864_ (.A(_08482_),
    .X(_12432_));
 sky130_fd_sc_hd__o31a_1 _39865_ (.A1(_12432_),
    .A2(_10083_),
    .A3(_11278_),
    .B1(_11283_),
    .X(_12433_));
 sky130_fd_sc_hd__xor2_1 _39866_ (.A(_12431_),
    .B(_12433_),
    .X(_12434_));
 sky130_fd_sc_hd__xnor2_1 _39867_ (.A(_12424_),
    .B(_12434_),
    .Y(_12435_));
 sky130_fd_sc_hd__a21o_1 _39868_ (.A1(_11287_),
    .A2(_11290_),
    .B1(_12435_),
    .X(_12436_));
 sky130_fd_sc_hd__inv_2 _39869_ (.A(_12436_),
    .Y(_12437_));
 sky130_fd_sc_hd__o311a_1 _39870_ (.A1(_11270_),
    .A2(_11271_),
    .A3(_11289_),
    .B1(_12435_),
    .C1(_11287_),
    .X(_12439_));
 sky130_fd_sc_hd__nor2_1 _39871_ (.A(_12437_),
    .B(_12439_),
    .Y(_12440_));
 sky130_fd_sc_hd__o2111a_1 _39872_ (.A1(_12419_),
    .A2(_12421_),
    .B1(_12440_),
    .C1(_11269_),
    .D1(_07171_),
    .X(_12441_));
 sky130_fd_sc_hd__nor2_1 _39873_ (.A(_11270_),
    .B(_12440_),
    .Y(_12442_));
 sky130_fd_sc_hd__nor2_1 _39874_ (.A(_12441_),
    .B(_12442_),
    .Y(_12443_));
 sky130_fd_sc_hd__nor2_1 _39875_ (.A(_12418_),
    .B(_12443_),
    .Y(_12444_));
 sky130_fd_sc_hd__nand2_1 _39876_ (.A(_12443_),
    .B(_12418_),
    .Y(_12445_));
 sky130_fd_sc_hd__or2b_1 _39877_ (.A(_12444_),
    .B_N(_12445_),
    .X(_12446_));
 sky130_fd_sc_hd__a21o_1 _39878_ (.A1(_10098_),
    .A2(_10100_),
    .B1(_11298_),
    .X(_12447_));
 sky130_fd_sc_hd__a21boi_1 _39879_ (.A1(_11300_),
    .A2(_11299_),
    .B1_N(_12447_),
    .Y(_12448_));
 sky130_fd_sc_hd__or2_1 _39880_ (.A(_12446_),
    .B(_12448_),
    .X(_12450_));
 sky130_fd_sc_hd__nand2_1 _39881_ (.A(_12448_),
    .B(_12446_),
    .Y(_12451_));
 sky130_fd_sc_hd__o21bai_2 _39882_ (.A1(_11265_),
    .A2(_11232_),
    .B1_N(_11263_),
    .Y(_12452_));
 sky130_fd_sc_hd__buf_1 _39883_ (.A(_00514_),
    .X(_12453_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _39884_ (.A(_02367_),
    .X(_12454_));
 sky130_fd_sc_hd__o21a_1 _39885_ (.A1(_12453_),
    .A2(_12454_),
    .B1(_08453_),
    .X(_12455_));
 sky130_fd_sc_hd__nor3_1 _39886_ (.A(_12453_),
    .B(_08453_),
    .C(_12454_),
    .Y(_12456_));
 sky130_fd_sc_hd__or3b_2 _39887_ (.A(_08456_),
    .B(_10044_),
    .C_N(_07121_),
    .X(_12457_));
 sky130_fd_sc_hd__nor2_1 _39888_ (.A(\delay_line[22][14] ),
    .B(_10037_),
    .Y(_12458_));
 sky130_fd_sc_hd__nor2_1 _39889_ (.A(_07119_),
    .B(_10044_),
    .Y(_12459_));
 sky130_fd_sc_hd__a2bb2o_1 _39890_ (.A1_N(_12458_),
    .A2_N(_12459_),
    .B1(_11236_),
    .B2(_10037_),
    .X(_12461_));
 sky130_fd_sc_hd__o211ai_2 _39891_ (.A1(_12455_),
    .A2(_12456_),
    .B1(_12457_),
    .C1(_12461_),
    .Y(_12462_));
 sky130_fd_sc_hd__a211o_1 _39892_ (.A1(_12457_),
    .A2(_12461_),
    .B1(_12455_),
    .C1(_12456_),
    .X(_12463_));
 sky130_fd_sc_hd__nand2_1 _39893_ (.A(_12462_),
    .B(_12463_),
    .Y(_12464_));
 sky130_fd_sc_hd__a21oi_1 _39894_ (.A1(_11245_),
    .A2(_11244_),
    .B1(_12464_),
    .Y(_12465_));
 sky130_fd_sc_hd__a21o_1 _39895_ (.A1(_12454_),
    .A2(_10034_),
    .B1(_10047_),
    .X(_12466_));
 sky130_fd_sc_hd__and3_1 _39896_ (.A(_11245_),
    .B(_11244_),
    .C(_12464_),
    .X(_12467_));
 sky130_fd_sc_hd__or3_1 _39897_ (.A(_12465_),
    .B(_12466_),
    .C(_12467_),
    .X(_12468_));
 sky130_fd_sc_hd__buf_1 _39898_ (.A(_12454_),
    .X(_12469_));
 sky130_fd_sc_hd__nand2_1 _39899_ (.A(_12469_),
    .B(_10034_),
    .Y(_12470_));
 sky130_fd_sc_hd__a2bb2o_1 _39900_ (.A1_N(_12467_),
    .A2_N(_12465_),
    .B1(_12453_),
    .B2(_12470_),
    .X(_12472_));
 sky130_fd_sc_hd__and2_1 _39901_ (.A(_12468_),
    .B(_12472_),
    .X(_12473_));
 sky130_fd_sc_hd__nor3_1 _39902_ (.A(_11247_),
    .B(_11252_),
    .C(_12473_),
    .Y(_12474_));
 sky130_fd_sc_hd__o21ai_1 _39903_ (.A1(_11247_),
    .A2(_11252_),
    .B1(_12473_),
    .Y(_12475_));
 sky130_fd_sc_hd__and2b_1 _39904_ (.A_N(_12474_),
    .B(_12475_),
    .X(_12476_));
 sky130_fd_sc_hd__xnor2_1 _39905_ (.A(_11234_),
    .B(_12476_),
    .Y(_12477_));
 sky130_fd_sc_hd__a21boi_1 _39906_ (.A1(_11253_),
    .A2(_11258_),
    .B1_N(_12477_),
    .Y(_12478_));
 sky130_fd_sc_hd__a211oi_1 _39907_ (.A1(_11256_),
    .A2(_11255_),
    .B1(_11259_),
    .C1(_12477_),
    .Y(_12479_));
 sky130_fd_sc_hd__or2_1 _39908_ (.A(_12478_),
    .B(_12479_),
    .X(_12480_));
 sky130_fd_sc_hd__xnor2_2 _39909_ (.A(_12452_),
    .B(_12480_),
    .Y(_12481_));
 sky130_fd_sc_hd__a21o_1 _39910_ (.A1(_12450_),
    .A2(_12451_),
    .B1(_12481_),
    .X(_12483_));
 sky130_fd_sc_hd__nand3_2 _39911_ (.A(_12450_),
    .B(_12451_),
    .C(_12481_),
    .Y(_12484_));
 sky130_fd_sc_hd__nand2_1 _39912_ (.A(_12483_),
    .B(_12484_),
    .Y(_12485_));
 sky130_fd_sc_hd__nand2_1 _39913_ (.A(_12417_),
    .B(_12485_),
    .Y(_12486_));
 sky130_fd_sc_hd__or2_1 _39914_ (.A(_12417_),
    .B(_12485_),
    .X(_12487_));
 sky130_fd_sc_hd__and2_1 _39915_ (.A(_12486_),
    .B(_12487_),
    .X(_12488_));
 sky130_fd_sc_hd__nor2_1 _39916_ (.A(_12389_),
    .B(_12488_),
    .Y(_12489_));
 sky130_fd_sc_hd__nand2_1 _39917_ (.A(_12488_),
    .B(_12389_),
    .Y(_12490_));
 sky130_fd_sc_hd__and2b_1 _39918_ (.A_N(_12489_),
    .B(_12490_),
    .X(_12491_));
 sky130_fd_sc_hd__xor2_1 _39919_ (.A(_12388_),
    .B(_12491_),
    .X(_12492_));
 sky130_fd_sc_hd__a21boi_4 _39920_ (.A1(_12382_),
    .A2(_12384_),
    .B1_N(_12175_),
    .Y(_12494_));
 sky130_fd_sc_hd__or2_1 _39921_ (.A(_12492_),
    .B(_12494_),
    .X(_12495_));
 sky130_fd_sc_hd__o21ai_1 _39922_ (.A1(_12494_),
    .A2(_12386_),
    .B1(_12492_),
    .Y(_12496_));
 sky130_fd_sc_hd__o21ai_1 _39923_ (.A1(_12386_),
    .A2(_12495_),
    .B1(_12496_),
    .Y(_12497_));
 sky130_fd_sc_hd__a21oi_1 _39924_ (.A1(_11314_),
    .A2(_11312_),
    .B1(_12497_),
    .Y(_12498_));
 sky130_fd_sc_hd__o211ai_1 _39925_ (.A1(_11197_),
    .A2(_11311_),
    .B1(_11314_),
    .C1(_12497_),
    .Y(_12499_));
 sky130_fd_sc_hd__or2b_1 _39926_ (.A(_12498_),
    .B_N(_12499_),
    .X(_12500_));
 sky130_fd_sc_hd__and2b_1 _39927_ (.A_N(_11324_),
    .B(_11378_),
    .X(_12501_));
 sky130_fd_sc_hd__a21oi_2 _39928_ (.A1(_11458_),
    .A2(_11379_),
    .B1(_12501_),
    .Y(_12502_));
 sky130_fd_sc_hd__a21o_1 _39929_ (.A1(_11308_),
    .A2(_11310_),
    .B1(_11307_),
    .X(_12503_));
 sky130_fd_sc_hd__and3_1 _39930_ (.A(_04409_),
    .B(_11442_),
    .C(_11443_),
    .X(_12505_));
 sky130_fd_sc_hd__and3_1 _39931_ (.A(_11442_),
    .B(_06941_),
    .C(_11443_),
    .X(_12506_));
 sky130_fd_sc_hd__a2bb2o_1 _39932_ (.A1_N(_06941_),
    .A2_N(_12505_),
    .B1(_12506_),
    .B2(_04409_),
    .X(_12507_));
 sky130_fd_sc_hd__o211a_1 _39933_ (.A1(_11444_),
    .A2(_11445_),
    .B1(_08886_),
    .C1(_10186_),
    .X(_12508_));
 sky130_fd_sc_hd__or3_2 _39934_ (.A(_12507_),
    .B(_12508_),
    .C(_11452_),
    .X(_12509_));
 sky130_fd_sc_hd__o21ai_2 _39935_ (.A1(_11452_),
    .A2(_12508_),
    .B1(_12507_),
    .Y(_12510_));
 sky130_fd_sc_hd__o21ai_2 _39936_ (.A1(_10225_),
    .A2(_11434_),
    .B1(_11440_),
    .Y(_12511_));
 sky130_fd_sc_hd__nor2_1 _39937_ (.A(_11412_),
    .B(_11417_),
    .Y(_12512_));
 sky130_fd_sc_hd__buf_1 _39938_ (.A(_08896_),
    .X(_12513_));
 sky130_fd_sc_hd__and3_1 _39939_ (.A(_12513_),
    .B(_10204_),
    .C(_10217_),
    .X(_12514_));
 sky130_fd_sc_hd__a21oi_1 _39940_ (.A1(_12513_),
    .A2(_10217_),
    .B1(_10204_),
    .Y(_12516_));
 sky130_fd_sc_hd__a21oi_1 _39941_ (.A1(_10199_),
    .A2(_10211_),
    .B1(_10213_),
    .Y(_12517_));
 sky130_fd_sc_hd__a2111oi_1 _39942_ (.A1(_10217_),
    .A2(_10203_),
    .B1(_11413_),
    .C1(_12517_),
    .D1(_06925_),
    .Y(_12518_));
 sky130_fd_sc_hd__and3_1 _39943_ (.A(_02110_),
    .B(_10199_),
    .C(_10211_),
    .X(_12519_));
 sky130_fd_sc_hd__o22a_1 _39944_ (.A1(_06925_),
    .A2(_11413_),
    .B1(_12519_),
    .B2(_12517_),
    .X(_12520_));
 sky130_fd_sc_hd__nor4_1 _39945_ (.A(_12514_),
    .B(_12516_),
    .C(net188),
    .D(_12520_),
    .Y(_12521_));
 sky130_fd_sc_hd__o22a_1 _39946_ (.A1(_12514_),
    .A2(_12516_),
    .B1(net188),
    .B2(_12520_),
    .X(_12522_));
 sky130_fd_sc_hd__a32o_1 _39947_ (.A1(_11410_),
    .A2(_11423_),
    .A3(_10210_),
    .B1(_11420_),
    .B2(_11421_),
    .X(_12523_));
 sky130_fd_sc_hd__nor3b_1 _39948_ (.A(_12521_),
    .B(_12522_),
    .C_N(_12523_),
    .Y(_12524_));
 sky130_fd_sc_hd__o21ba_1 _39949_ (.A1(_12521_),
    .A2(_12522_),
    .B1_N(_12523_),
    .X(_12525_));
 sky130_fd_sc_hd__or3_1 _39950_ (.A(_12512_),
    .B(_12524_),
    .C(_12525_),
    .X(_12527_));
 sky130_fd_sc_hd__inv_2 _39951_ (.A(_12527_),
    .Y(_12528_));
 sky130_fd_sc_hd__o21a_1 _39952_ (.A1(net164),
    .A2(_12525_),
    .B1(_12512_),
    .X(_12529_));
 sky130_fd_sc_hd__a21boi_1 _39953_ (.A1(_11408_),
    .A2(_11425_),
    .B1_N(_11426_),
    .Y(_12530_));
 sky130_fd_sc_hd__nor3_1 _39954_ (.A(_12528_),
    .B(_12529_),
    .C(_12530_),
    .Y(_12531_));
 sky130_fd_sc_hd__o21a_1 _39955_ (.A1(_12528_),
    .A2(_12529_),
    .B1(_12530_),
    .X(_12532_));
 sky130_fd_sc_hd__nor2_1 _39956_ (.A(_12531_),
    .B(_12532_),
    .Y(_12533_));
 sky130_fd_sc_hd__o31a_1 _39957_ (.A1(_11428_),
    .A2(_11429_),
    .A3(_11430_),
    .B1(_12533_),
    .X(_12534_));
 sky130_fd_sc_hd__nor2_1 _39958_ (.A(_11431_),
    .B(_12533_),
    .Y(_12535_));
 sky130_fd_sc_hd__nor2_1 _39959_ (.A(_12534_),
    .B(_12535_),
    .Y(_12536_));
 sky130_fd_sc_hd__nand3_2 _39960_ (.A(_11437_),
    .B(_12511_),
    .C(_12536_),
    .Y(_12538_));
 sky130_fd_sc_hd__o2bb2ai_4 _39961_ (.A1_N(_11437_),
    .A2_N(_12511_),
    .B1(_12534_),
    .B2(_12535_),
    .Y(_12539_));
 sky130_fd_sc_hd__a22oi_4 _39962_ (.A1(_12509_),
    .A2(_12510_),
    .B1(_12538_),
    .B2(_12539_),
    .Y(_12540_));
 sky130_fd_sc_hd__nand4_4 _39963_ (.A(_12509_),
    .B(_12510_),
    .C(_12538_),
    .D(_12539_),
    .Y(_12541_));
 sky130_fd_sc_hd__inv_2 _39964_ (.A(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__xnor2_1 _39965_ (.A(_10237_),
    .B(_08857_),
    .Y(_12543_));
 sky130_fd_sc_hd__xnor2_1 _39966_ (.A(_12543_),
    .B(_11384_),
    .Y(_12544_));
 sky130_fd_sc_hd__xnor2_1 _39967_ (.A(_11391_),
    .B(_12544_),
    .Y(_12545_));
 sky130_fd_sc_hd__xor2_2 _39968_ (.A(_11387_),
    .B(_12545_),
    .X(_12546_));
 sky130_fd_sc_hd__o21ai_1 _39969_ (.A1(_11393_),
    .A2(_11398_),
    .B1(_12546_),
    .Y(_12547_));
 sky130_fd_sc_hd__or3_1 _39970_ (.A(_11393_),
    .B(_11398_),
    .C(_12546_),
    .X(_12549_));
 sky130_fd_sc_hd__nand2_1 _39971_ (.A(_12547_),
    .B(_12549_),
    .Y(_12550_));
 sky130_fd_sc_hd__inv_2 _39972_ (.A(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__a21oi_2 _39973_ (.A1(_10256_),
    .A2(_11399_),
    .B1(_11403_),
    .Y(_12552_));
 sky130_fd_sc_hd__xor2_4 _39974_ (.A(_12551_),
    .B(_12552_),
    .X(_12553_));
 sky130_fd_sc_hd__o21a_1 _39975_ (.A1(_12540_),
    .A2(_12542_),
    .B1(_12553_),
    .X(_12554_));
 sky130_fd_sc_hd__nor3_1 _39976_ (.A(_12540_),
    .B(_12542_),
    .C(_12553_),
    .Y(_12555_));
 sky130_fd_sc_hd__o21bai_4 _39977_ (.A1(_11335_),
    .A2(_11377_),
    .B1_N(_11375_),
    .Y(_12556_));
 sky130_fd_sc_hd__nor2_1 _39978_ (.A(_11332_),
    .B(_11334_),
    .Y(_12557_));
 sky130_fd_sc_hd__buf_1 _39979_ (.A(_06999_),
    .X(_12558_));
 sky130_fd_sc_hd__a2bb2o_1 _39980_ (.A1_N(_12558_),
    .A2_N(_10168_),
    .B1(_08784_),
    .B2(_05559_),
    .X(_12560_));
 sky130_fd_sc_hd__o21ba_1 _39981_ (.A1(_06990_),
    .A2(_12560_),
    .B1_N(_06994_),
    .X(_12561_));
 sky130_fd_sc_hd__nand2_1 _39982_ (.A(_11329_),
    .B(_12561_),
    .Y(_12562_));
 sky130_fd_sc_hd__a2111o_2 _39983_ (.A1(_08785_),
    .A2(_10172_),
    .B1(_11325_),
    .C1(_11326_),
    .D1(_12561_),
    .X(_12563_));
 sky130_fd_sc_hd__o211ai_4 _39984_ (.A1(_11330_),
    .A2(_12557_),
    .B1(_12562_),
    .C1(_12563_),
    .Y(_12564_));
 sky130_fd_sc_hd__a211o_1 _39985_ (.A1(_12562_),
    .A2(_12563_),
    .B1(_11330_),
    .C1(_12557_),
    .X(_12565_));
 sky130_fd_sc_hd__nand2_2 _39986_ (.A(_12564_),
    .B(_12565_),
    .Y(_12566_));
 sky130_fd_sc_hd__nor2_1 _39987_ (.A(_11370_),
    .B(_11373_),
    .Y(_12567_));
 sky130_fd_sc_hd__nand2_1 _39988_ (.A(_04320_),
    .B(_04321_),
    .Y(_12568_));
 sky130_fd_sc_hd__xor2_1 _39989_ (.A(_12568_),
    .B(_11358_),
    .X(_12569_));
 sky130_fd_sc_hd__o31a_1 _39990_ (.A1(_00966_),
    .A2(_02215_),
    .A3(_02220_),
    .B1(_12569_),
    .X(_12571_));
 sky130_fd_sc_hd__nor2_1 _39991_ (.A(_05509_),
    .B(_12569_),
    .Y(_12572_));
 sky130_fd_sc_hd__or2_1 _39992_ (.A(_12571_),
    .B(_12572_),
    .X(_12573_));
 sky130_fd_sc_hd__inv_2 _39993_ (.A(_11363_),
    .Y(_12574_));
 sky130_fd_sc_hd__o21ai_1 _39994_ (.A1(_11362_),
    .A2(net191),
    .B1(_12574_),
    .Y(_12575_));
 sky130_fd_sc_hd__xnor2_1 _39995_ (.A(_12573_),
    .B(_12575_),
    .Y(_12576_));
 sky130_fd_sc_hd__or3_1 _39996_ (.A(_11367_),
    .B(_12567_),
    .C(_12576_),
    .X(_12577_));
 sky130_fd_sc_hd__o21ai_2 _39997_ (.A1(_11367_),
    .A2(_12567_),
    .B1(_12576_),
    .Y(_12578_));
 sky130_fd_sc_hd__buf_1 _39998_ (.A(_11343_),
    .X(_12579_));
 sky130_fd_sc_hd__a2111o_1 _39999_ (.A1(_08804_),
    .A2(_07018_),
    .B1(_08809_),
    .C1(_10154_),
    .D1(_10155_),
    .X(_12580_));
 sky130_fd_sc_hd__o32a_1 _40000_ (.A1(_12579_),
    .A2(_11344_),
    .A3(_12580_),
    .B1(_11336_),
    .B2(_11347_),
    .X(_12582_));
 sky130_fd_sc_hd__nand2_1 _40001_ (.A(_11337_),
    .B(_07013_),
    .Y(_12583_));
 sky130_fd_sc_hd__buf_1 _40002_ (.A(net334),
    .X(_12584_));
 sky130_fd_sc_hd__o21ai_1 _40003_ (.A1(net335),
    .A2(net334),
    .B1(_00995_),
    .Y(_12585_));
 sky130_fd_sc_hd__a21oi_1 _40004_ (.A1(_05531_),
    .A2(_12584_),
    .B1(_12585_),
    .Y(_12586_));
 sky130_fd_sc_hd__and2_1 _40005_ (.A(net335),
    .B(net334),
    .X(_12587_));
 sky130_fd_sc_hd__nor2_1 _40006_ (.A(_05531_),
    .B(_12584_),
    .Y(_12588_));
 sky130_fd_sc_hd__o21ba_1 _40007_ (.A1(_12587_),
    .A2(_12588_),
    .B1_N(_00995_),
    .X(_12589_));
 sky130_fd_sc_hd__a211oi_2 _40008_ (.A1(_12583_),
    .A2(_11341_),
    .B1(_12586_),
    .C1(_12589_),
    .Y(_12590_));
 sky130_fd_sc_hd__o211a_1 _40009_ (.A1(_12586_),
    .A2(_12589_),
    .B1(_12583_),
    .C1(_11341_),
    .X(_12591_));
 sky130_fd_sc_hd__a2111oi_1 _40010_ (.A1(_10154_),
    .A2(_11345_),
    .B1(_12590_),
    .C1(_12591_),
    .D1(_12579_),
    .Y(_12593_));
 sky130_fd_sc_hd__a2111oi_1 _40011_ (.A1(_10147_),
    .A2(_08807_),
    .B1(_10153_),
    .C1(_11343_),
    .D1(_11344_),
    .Y(_12594_));
 sky130_fd_sc_hd__o22a_1 _40012_ (.A1(_12590_),
    .A2(_12591_),
    .B1(net244),
    .B2(_12579_),
    .X(_12595_));
 sky130_fd_sc_hd__nor3_1 _40013_ (.A(_11349_),
    .B(net217),
    .C(_12595_),
    .Y(_12596_));
 sky130_fd_sc_hd__o21a_1 _40014_ (.A1(net216),
    .A2(_12595_),
    .B1(_11349_),
    .X(_12597_));
 sky130_fd_sc_hd__nor2_1 _40015_ (.A(_12596_),
    .B(_12597_),
    .Y(_12598_));
 sky130_fd_sc_hd__xnor2_1 _40016_ (.A(_12582_),
    .B(_12598_),
    .Y(_12599_));
 sky130_fd_sc_hd__nand3_1 _40017_ (.A(_10160_),
    .B(_10162_),
    .C(_11352_),
    .Y(_12600_));
 sky130_fd_sc_hd__o21ai_1 _40018_ (.A1(_11351_),
    .A2(_11348_),
    .B1(_12600_),
    .Y(_12601_));
 sky130_fd_sc_hd__xnor2_1 _40019_ (.A(_12599_),
    .B(_12601_),
    .Y(_12602_));
 sky130_fd_sc_hd__and3_1 _40020_ (.A(_12577_),
    .B(_12578_),
    .C(_12602_),
    .X(_12604_));
 sky130_fd_sc_hd__a21oi_1 _40021_ (.A1(_12577_),
    .A2(_12578_),
    .B1(_12602_),
    .Y(_12605_));
 sky130_fd_sc_hd__nor2_2 _40022_ (.A(_12604_),
    .B(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__xnor2_4 _40023_ (.A(_12566_),
    .B(_12606_),
    .Y(_12607_));
 sky130_fd_sc_hd__xnor2_1 _40024_ (.A(_12556_),
    .B(_12607_),
    .Y(_12608_));
 sky130_fd_sc_hd__o21ai_1 _40025_ (.A1(_12554_),
    .A2(net80),
    .B1(_12608_),
    .Y(_12609_));
 sky130_fd_sc_hd__or3_1 _40026_ (.A(_12554_),
    .B(net80),
    .C(_12608_),
    .X(_12610_));
 sky130_fd_sc_hd__nand2_1 _40027_ (.A(_12609_),
    .B(_12610_),
    .Y(_12611_));
 sky130_fd_sc_hd__xnor2_1 _40028_ (.A(_12503_),
    .B(_12611_),
    .Y(_12612_));
 sky130_fd_sc_hd__xor2_1 _40029_ (.A(_12502_),
    .B(_12612_),
    .X(_12613_));
 sky130_fd_sc_hd__inv_2 _40030_ (.A(_12613_),
    .Y(_12615_));
 sky130_fd_sc_hd__xnor2_1 _40031_ (.A(_12500_),
    .B(_12615_),
    .Y(_12616_));
 sky130_fd_sc_hd__xnor2_1 _40032_ (.A(_12173_),
    .B(_12616_),
    .Y(_12617_));
 sky130_fd_sc_hd__and2_1 _40033_ (.A(_11558_),
    .B(_11608_),
    .X(_12618_));
 sky130_fd_sc_hd__o21bai_4 _40034_ (.A1(_11553_),
    .A2(_11552_),
    .B1_N(_11551_),
    .Y(_12619_));
 sky130_fd_sc_hd__inv_2 _40035_ (.A(_11545_),
    .Y(_12620_));
 sky130_fd_sc_hd__o21ai_2 _40036_ (.A1(_11490_),
    .A2(_12620_),
    .B1(_11544_),
    .Y(_12621_));
 sky130_fd_sc_hd__and2_1 _40037_ (.A(_11486_),
    .B(_11485_),
    .X(_12622_));
 sky130_fd_sc_hd__or3b_1 _40038_ (.A(_06786_),
    .B(_08295_),
    .C_N(_08286_),
    .X(_12623_));
 sky130_fd_sc_hd__a21bo_1 _40039_ (.A1(_12623_),
    .A2(_11476_),
    .B1_N(_08284_),
    .X(_12624_));
 sky130_fd_sc_hd__nand2_1 _40040_ (.A(_12623_),
    .B(_06785_),
    .Y(_12626_));
 sky130_fd_sc_hd__a211o_1 _40041_ (.A1(_12624_),
    .A2(_12626_),
    .B1(_11480_),
    .C1(net177),
    .X(_12627_));
 sky130_fd_sc_hd__o211ai_2 _40042_ (.A1(_11480_),
    .A2(net177),
    .B1(_12624_),
    .C1(_12626_),
    .Y(_12628_));
 sky130_fd_sc_hd__and2_1 _40043_ (.A(_12627_),
    .B(_12628_),
    .X(_12629_));
 sky130_fd_sc_hd__o21ai_2 _40044_ (.A1(_12622_),
    .A2(_11488_),
    .B1(_12629_),
    .Y(_12630_));
 sky130_fd_sc_hd__or3_1 _40045_ (.A(_12622_),
    .B(_11488_),
    .C(_12629_),
    .X(_12631_));
 sky130_fd_sc_hd__nand2_1 _40046_ (.A(_12630_),
    .B(_12631_),
    .Y(_12632_));
 sky130_fd_sc_hd__clkbuf_2 _40047_ (.A(_03812_),
    .X(_12633_));
 sky130_fd_sc_hd__xnor2_1 _40048_ (.A(_05207_),
    .B(_12633_),
    .Y(_12634_));
 sky130_fd_sc_hd__and2b_1 _40049_ (.A_N(_09588_),
    .B(_11524_),
    .X(_12635_));
 sky130_fd_sc_hd__nand2_1 _40050_ (.A(_12634_),
    .B(_12635_),
    .Y(_12637_));
 sky130_fd_sc_hd__or2_1 _40051_ (.A(_12634_),
    .B(_12635_),
    .X(_12638_));
 sky130_fd_sc_hd__a21o_1 _40052_ (.A1(_12637_),
    .A2(_12638_),
    .B1(_06847_),
    .X(_12639_));
 sky130_fd_sc_hd__clkbuf_2 _40053_ (.A(_06847_),
    .X(_12640_));
 sky130_fd_sc_hd__nand3_2 _40054_ (.A(_12638_),
    .B(_12640_),
    .C(_12637_),
    .Y(_12641_));
 sky130_fd_sc_hd__nand3_1 _40055_ (.A(_12639_),
    .B(_11530_),
    .C(_12641_),
    .Y(_12642_));
 sky130_fd_sc_hd__a32o_1 _40056_ (.A1(_11529_),
    .A2(_11525_),
    .A3(_11527_),
    .B1(_12641_),
    .B2(_12639_),
    .X(_12643_));
 sky130_fd_sc_hd__nand2_1 _40057_ (.A(_12642_),
    .B(_12643_),
    .Y(_12644_));
 sky130_fd_sc_hd__o21ba_1 _40058_ (.A1(_09589_),
    .A2(_11531_),
    .B1_N(_11532_),
    .X(_12645_));
 sky130_fd_sc_hd__nor2_1 _40059_ (.A(_12644_),
    .B(_12645_),
    .Y(_12646_));
 sky130_fd_sc_hd__and3b_1 _40060_ (.A_N(_11532_),
    .B(_11533_),
    .C(_12644_),
    .X(_12648_));
 sky130_fd_sc_hd__nand2_1 _40061_ (.A(_11542_),
    .B(_11540_),
    .Y(_12649_));
 sky130_fd_sc_hd__and2_1 _40062_ (.A(_11538_),
    .B(_12649_),
    .X(_12650_));
 sky130_fd_sc_hd__o21ai_1 _40063_ (.A1(_12646_),
    .A2(_12648_),
    .B1(_12650_),
    .Y(_12651_));
 sky130_fd_sc_hd__or2_2 _40064_ (.A(_12646_),
    .B(_12648_),
    .X(_12652_));
 sky130_fd_sc_hd__a21o_1 _40065_ (.A1(_11538_),
    .A2(_12649_),
    .B1(_12652_),
    .X(_12653_));
 sky130_fd_sc_hd__a21o_1 _40066_ (.A1(_12651_),
    .A2(_12653_),
    .B1(_11536_),
    .X(_12654_));
 sky130_fd_sc_hd__a21bo_2 _40067_ (.A1(_12649_),
    .A2(_12652_),
    .B1_N(_11536_),
    .X(_12655_));
 sky130_fd_sc_hd__a21bo_1 _40068_ (.A1(_08322_),
    .A2(_09614_),
    .B1_N(_11498_),
    .X(_12656_));
 sky130_fd_sc_hd__or2_1 _40069_ (.A(_11496_),
    .B(_11501_),
    .X(_12657_));
 sky130_fd_sc_hd__buf_1 _40070_ (.A(\delay_line[33][14] ),
    .X(_12659_));
 sky130_fd_sc_hd__buf_1 _40071_ (.A(_11494_),
    .X(_12660_));
 sky130_fd_sc_hd__or3b_1 _40072_ (.A(_09633_),
    .B(_12659_),
    .C_N(_12660_),
    .X(_12661_));
 sky130_fd_sc_hd__nand4_1 _40073_ (.A(_06812_),
    .B(_12657_),
    .C(_12661_),
    .D(_09619_),
    .Y(_12662_));
 sky130_fd_sc_hd__a22o_1 _40074_ (.A1(_06812_),
    .A2(_09619_),
    .B1(_12657_),
    .B2(_12661_),
    .X(_12663_));
 sky130_fd_sc_hd__clkbuf_2 _40075_ (.A(_09617_),
    .X(_12664_));
 sky130_fd_sc_hd__mux2_1 _40076_ (.A0(_12659_),
    .A1(_12660_),
    .S(_12664_),
    .X(_12665_));
 sky130_fd_sc_hd__and3_1 _40077_ (.A(_12662_),
    .B(_12663_),
    .C(_12665_),
    .X(_12666_));
 sky130_fd_sc_hd__a21oi_1 _40078_ (.A1(_12662_),
    .A2(_12663_),
    .B1(_12665_),
    .Y(_12667_));
 sky130_fd_sc_hd__nor2_1 _40079_ (.A(_12666_),
    .B(_12667_),
    .Y(_12668_));
 sky130_fd_sc_hd__o41a_1 _40080_ (.A1(_09610_),
    .A2(_09615_),
    .A3(_11501_),
    .A4(_11500_),
    .B1(_11505_),
    .X(_12670_));
 sky130_fd_sc_hd__xnor2_1 _40081_ (.A(_12668_),
    .B(_12670_),
    .Y(_12671_));
 sky130_fd_sc_hd__xnor2_1 _40082_ (.A(_12656_),
    .B(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__a21oi_2 _40083_ (.A1(_11509_),
    .A2(_11510_),
    .B1(_12672_),
    .Y(_12673_));
 sky130_fd_sc_hd__and3_1 _40084_ (.A(_11509_),
    .B(_11510_),
    .C(_12672_),
    .X(_12674_));
 sky130_fd_sc_hd__a2111oi_1 _40085_ (.A1(_09631_),
    .A2(_11491_),
    .B1(_12673_),
    .C1(_11513_),
    .D1(_12674_),
    .Y(_12675_));
 sky130_fd_sc_hd__nor2_1 _40086_ (.A(_12674_),
    .B(_12673_),
    .Y(_12676_));
 sky130_fd_sc_hd__nor2_1 _40087_ (.A(_11516_),
    .B(_12676_),
    .Y(_12677_));
 sky130_fd_sc_hd__nor2_1 _40088_ (.A(net126),
    .B(_12677_),
    .Y(_12678_));
 sky130_fd_sc_hd__o21a_1 _40089_ (.A1(_11518_),
    .A2(_11521_),
    .B1(_12678_),
    .X(_12679_));
 sky130_fd_sc_hd__a211oi_1 _40090_ (.A1(_09639_),
    .A2(_11517_),
    .B1(_11521_),
    .C1(_12678_),
    .Y(_12681_));
 sky130_fd_sc_hd__nor2_1 _40091_ (.A(_12679_),
    .B(_12681_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand3_1 _40092_ (.A(_12654_),
    .B(_12655_),
    .C(_12682_),
    .Y(_12683_));
 sky130_fd_sc_hd__a21o_1 _40093_ (.A1(_12654_),
    .A2(_12655_),
    .B1(_12682_),
    .X(_12684_));
 sky130_fd_sc_hd__nand2_2 _40094_ (.A(_12683_),
    .B(_12684_),
    .Y(_12685_));
 sky130_fd_sc_hd__o21ai_1 _40095_ (.A1(_11435_),
    .A2(_11441_),
    .B1(_11453_),
    .Y(_12686_));
 sky130_fd_sc_hd__a21oi_4 _40096_ (.A1(_12686_),
    .A2(_11406_),
    .B1(_11455_),
    .Y(_12687_));
 sky130_fd_sc_hd__a21oi_1 _40097_ (.A1(_12632_),
    .A2(_12685_),
    .B1(_12687_),
    .Y(_12688_));
 sky130_fd_sc_hd__o21ai_2 _40098_ (.A1(_12632_),
    .A2(_12685_),
    .B1(_12688_),
    .Y(_12689_));
 sky130_fd_sc_hd__xnor2_1 _40099_ (.A(_12632_),
    .B(_12685_),
    .Y(_12690_));
 sky130_fd_sc_hd__nand2_1 _40100_ (.A(_12690_),
    .B(_12687_),
    .Y(_12692_));
 sky130_fd_sc_hd__nand3_4 _40101_ (.A(_12621_),
    .B(_12689_),
    .C(_12692_),
    .Y(_12693_));
 sky130_fd_sc_hd__a21o_2 _40102_ (.A1(_12689_),
    .A2(_12692_),
    .B1(_12621_),
    .X(_12694_));
 sky130_fd_sc_hd__a21oi_1 _40103_ (.A1(_12693_),
    .A2(_12694_),
    .B1(_12619_),
    .Y(_12695_));
 sky130_fd_sc_hd__buf_1 _40104_ (.A(_09686_),
    .X(_12696_));
 sky130_fd_sc_hd__and2b_1 _40105_ (.A_N(_11567_),
    .B(_11577_),
    .X(_12697_));
 sky130_fd_sc_hd__a21oi_1 _40106_ (.A1(_11578_),
    .A2(_12696_),
    .B1(_12697_),
    .Y(_12698_));
 sky130_fd_sc_hd__and2b_1 _40107_ (.A_N(net294),
    .B(net295),
    .X(_12699_));
 sky130_fd_sc_hd__or2b_1 _40108_ (.A(\delay_line[36][14] ),
    .B_N(\delay_line[36][15] ),
    .X(_12700_));
 sky130_fd_sc_hd__or2b_1 _40109_ (.A(_12699_),
    .B_N(_12700_),
    .X(_12701_));
 sky130_fd_sc_hd__o211a_1 _40110_ (.A1(_09687_),
    .A2(_11562_),
    .B1(_11561_),
    .C1(_11560_),
    .X(_12703_));
 sky130_fd_sc_hd__a221oi_4 _40111_ (.A1(net294),
    .A2(_09691_),
    .B1(_11566_),
    .B2(_11563_),
    .C1(_12703_),
    .Y(_12704_));
 sky130_fd_sc_hd__xor2_1 _40112_ (.A(_12701_),
    .B(_12704_),
    .X(_12705_));
 sky130_fd_sc_hd__o211ai_2 _40113_ (.A1(_08262_),
    .A2(_08265_),
    .B1(_11575_),
    .C1(_11574_),
    .Y(_12706_));
 sky130_fd_sc_hd__xor2_1 _40114_ (.A(_08248_),
    .B(_11568_),
    .X(_12707_));
 sky130_fd_sc_hd__o21ba_1 _40115_ (.A1(_11571_),
    .A2(_09698_),
    .B1_N(_11569_),
    .X(_12708_));
 sky130_fd_sc_hd__xnor2_1 _40116_ (.A(_12707_),
    .B(_12708_),
    .Y(_12709_));
 sky130_fd_sc_hd__or3b_1 _40117_ (.A(_11569_),
    .B(_11571_),
    .C_N(_09702_),
    .X(_12710_));
 sky130_fd_sc_hd__nand3_1 _40118_ (.A(_12706_),
    .B(_12709_),
    .C(_12710_),
    .Y(_12711_));
 sky130_fd_sc_hd__a21o_1 _40119_ (.A1(_12706_),
    .A2(_12710_),
    .B1(_12709_),
    .X(_12712_));
 sky130_fd_sc_hd__nand3_2 _40120_ (.A(_12705_),
    .B(_12711_),
    .C(_12712_),
    .Y(_12714_));
 sky130_fd_sc_hd__a21o_1 _40121_ (.A1(_12711_),
    .A2(_12712_),
    .B1(_12705_),
    .X(_12715_));
 sky130_fd_sc_hd__a21oi_1 _40122_ (.A1(_12714_),
    .A2(_12715_),
    .B1(_12696_),
    .Y(_12716_));
 sky130_fd_sc_hd__and3_1 _40123_ (.A(_09686_),
    .B(_12714_),
    .C(_12715_),
    .X(_12717_));
 sky130_fd_sc_hd__nor3_1 _40124_ (.A(_12698_),
    .B(_12716_),
    .C(_12717_),
    .Y(_12718_));
 sky130_fd_sc_hd__o21ai_1 _40125_ (.A1(_12716_),
    .A2(_12717_),
    .B1(_12698_),
    .Y(_12719_));
 sky130_fd_sc_hd__and2b_1 _40126_ (.A_N(_12718_),
    .B(_12719_),
    .X(_12720_));
 sky130_fd_sc_hd__a21o_2 _40127_ (.A1(_11586_),
    .A2(_11590_),
    .B1(_11587_),
    .X(_12721_));
 sky130_fd_sc_hd__nor2_1 _40128_ (.A(_09721_),
    .B(_08215_),
    .Y(_12722_));
 sky130_fd_sc_hd__and2_1 _40129_ (.A(_09721_),
    .B(_08215_),
    .X(_12723_));
 sky130_fd_sc_hd__nor2_1 _40130_ (.A(_12722_),
    .B(_12723_),
    .Y(_12725_));
 sky130_fd_sc_hd__and2_1 _40131_ (.A(_12721_),
    .B(_12725_),
    .X(_12726_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40132_ (.A(_12725_),
    .X(_12727_));
 sky130_fd_sc_hd__nor2_1 _40133_ (.A(_12727_),
    .B(_12721_),
    .Y(_12728_));
 sky130_fd_sc_hd__or2_1 _40134_ (.A(_12726_),
    .B(_12728_),
    .X(_12729_));
 sky130_fd_sc_hd__xnor2_2 _40135_ (.A(_12720_),
    .B(_12729_),
    .Y(_12730_));
 sky130_fd_sc_hd__or2b_1 _40136_ (.A(_12695_),
    .B_N(_12730_),
    .X(_12731_));
 sky130_fd_sc_hd__a31o_1 _40137_ (.A1(_12619_),
    .A2(_12693_),
    .A3(_12694_),
    .B1(_12731_),
    .X(_12732_));
 sky130_fd_sc_hd__and3_1 _40138_ (.A(_12619_),
    .B(_12693_),
    .C(_12694_),
    .X(_12733_));
 sky130_fd_sc_hd__o21bai_1 _40139_ (.A1(_12733_),
    .A2(_12695_),
    .B1_N(_12730_),
    .Y(_12734_));
 sky130_fd_sc_hd__inv_2 _40140_ (.A(_11462_),
    .Y(_12736_));
 sky130_fd_sc_hd__o21ai_2 _40141_ (.A1(_11464_),
    .A2(_12736_),
    .B1(_11461_),
    .Y(_12737_));
 sky130_fd_sc_hd__a21oi_1 _40142_ (.A1(_12732_),
    .A2(_12734_),
    .B1(_12737_),
    .Y(_12738_));
 sky130_fd_sc_hd__o211ai_2 _40143_ (.A1(_12733_),
    .A2(_12731_),
    .B1(_12734_),
    .C1(_12737_),
    .Y(_12739_));
 sky130_fd_sc_hd__and2b_1 _40144_ (.A_N(_12738_),
    .B(_12739_),
    .X(_12740_));
 sky130_fd_sc_hd__xor2_1 _40145_ (.A(_12618_),
    .B(_12740_),
    .X(_12741_));
 sky130_fd_sc_hd__nand2_1 _40146_ (.A(_12617_),
    .B(_12741_),
    .Y(_12742_));
 sky130_fd_sc_hd__or2_1 _40147_ (.A(_12617_),
    .B(_12741_),
    .X(_12743_));
 sky130_fd_sc_hd__o21ai_1 _40148_ (.A1(_10971_),
    .A2(_11470_),
    .B1(_11616_),
    .Y(_12744_));
 sky130_fd_sc_hd__a21oi_2 _40149_ (.A1(_12742_),
    .A2(_12743_),
    .B1(_12744_),
    .Y(_12745_));
 sky130_fd_sc_hd__and3_1 _40150_ (.A(_12744_),
    .B(_12742_),
    .C(_12743_),
    .X(_12747_));
 sky130_fd_sc_hd__nor2_1 _40151_ (.A(_12745_),
    .B(_12747_),
    .Y(_12748_));
 sky130_fd_sc_hd__o21ai_1 _40152_ (.A1(_12170_),
    .A2(_12172_),
    .B1(_12748_),
    .Y(_12749_));
 sky130_fd_sc_hd__o211ai_4 _40153_ (.A1(_11699_),
    .A2(_11700_),
    .B1(_12164_),
    .C1(_12169_),
    .Y(_12750_));
 sky130_fd_sc_hd__a21bo_1 _40154_ (.A1(_12164_),
    .A2(_12169_),
    .B1_N(_12171_),
    .X(_12751_));
 sky130_fd_sc_hd__o211ai_1 _40155_ (.A1(_12745_),
    .A2(_12747_),
    .B1(_12750_),
    .C1(_12751_),
    .Y(_12752_));
 sky130_fd_sc_hd__and3_1 _40156_ (.A(_10970_),
    .B(_11616_),
    .C(_11617_),
    .X(_12753_));
 sky130_fd_sc_hd__a31oi_1 _40157_ (.A1(_11623_),
    .A2(_11624_),
    .A3(_11619_),
    .B1(_12753_),
    .Y(_12754_));
 sky130_fd_sc_hd__nand3_2 _40158_ (.A(_12749_),
    .B(_12752_),
    .C(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__o21ai_1 _40159_ (.A1(_10963_),
    .A2(_09751_),
    .B1(_10966_),
    .Y(_12756_));
 sky130_fd_sc_hd__and3_1 _40160_ (.A(_10959_),
    .B(_10960_),
    .C(_10956_),
    .X(_12758_));
 sky130_fd_sc_hd__o2bb2ai_1 _40161_ (.A1_N(_10968_),
    .A2_N(_10962_),
    .B1(_12756_),
    .B2(_12758_),
    .Y(_12759_));
 sky130_fd_sc_hd__or3b_1 _40162_ (.A(_07520_),
    .B(_01452_),
    .C_N(_10296_),
    .X(_12760_));
 sky130_fd_sc_hd__or2_1 _40163_ (.A(_10467_),
    .B(_10461_),
    .X(_12761_));
 sky130_fd_sc_hd__nor2_2 _40164_ (.A(_08982_),
    .B(_08975_),
    .Y(_12762_));
 sky130_fd_sc_hd__and2_1 _40165_ (.A(_08975_),
    .B(_08982_),
    .X(_12763_));
 sky130_fd_sc_hd__clkbuf_2 _40166_ (.A(_08979_),
    .X(_12764_));
 sky130_fd_sc_hd__or3b_2 _40167_ (.A(_09001_),
    .B(_09003_),
    .C_N(net362),
    .X(_12765_));
 sky130_fd_sc_hd__or2_1 _40168_ (.A(_08999_),
    .B(_09007_),
    .X(_12766_));
 sky130_fd_sc_hd__and3_1 _40169_ (.A(_12764_),
    .B(_12765_),
    .C(_12766_),
    .X(_12767_));
 sky130_fd_sc_hd__a21oi_2 _40170_ (.A1(_12765_),
    .A2(_12766_),
    .B1(_12764_),
    .Y(_12769_));
 sky130_fd_sc_hd__o221a_1 _40171_ (.A1(_07550_),
    .A2(_10451_),
    .B1(_12767_),
    .B2(_12769_),
    .C1(_10454_),
    .X(_12770_));
 sky130_fd_sc_hd__a211oi_4 _40172_ (.A1(_10452_),
    .A2(_10454_),
    .B1(_12767_),
    .C1(_12769_),
    .Y(_12771_));
 sky130_fd_sc_hd__nor4_2 _40173_ (.A(_12762_),
    .B(_12763_),
    .C(_12770_),
    .D(_12771_),
    .Y(_12772_));
 sky130_fd_sc_hd__o22a_1 _40174_ (.A1(_12762_),
    .A2(_12763_),
    .B1(_12770_),
    .B2(_12771_),
    .X(_12773_));
 sky130_fd_sc_hd__or3_1 _40175_ (.A(_10461_),
    .B(_10450_),
    .C(_10462_),
    .X(_12774_));
 sky130_fd_sc_hd__o211ai_1 _40176_ (.A1(_12772_),
    .A2(_12773_),
    .B1(_10458_),
    .C1(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__a211o_1 _40177_ (.A1(_10458_),
    .A2(_12774_),
    .B1(_12772_),
    .C1(_12773_),
    .X(_12776_));
 sky130_fd_sc_hd__and4_1 _40178_ (.A(_12760_),
    .B(_12761_),
    .C(_12775_),
    .D(_12776_),
    .X(_12777_));
 sky130_fd_sc_hd__a22oi_1 _40179_ (.A1(_12760_),
    .A2(_12761_),
    .B1(_12775_),
    .B2(_12776_),
    .Y(_12778_));
 sky130_fd_sc_hd__nor2_2 _40180_ (.A(_12777_),
    .B(_12778_),
    .Y(_12780_));
 sky130_fd_sc_hd__or3b_1 _40181_ (.A(_12153_),
    .B(_10934_),
    .C_N(_03565_),
    .X(_12781_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40182_ (.A(_10436_),
    .X(_12782_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40183_ (.A(_06644_),
    .X(_12783_));
 sky130_fd_sc_hd__o2bb2a_1 _40184_ (.A1_N(_09006_),
    .A2_N(_12782_),
    .B1(_12783_),
    .B2(_10947_),
    .X(_12784_));
 sky130_fd_sc_hd__and3_1 _40185_ (.A(_09006_),
    .B(_12782_),
    .C(_10948_),
    .X(_12785_));
 sky130_fd_sc_hd__a211o_1 _40186_ (.A1(_10952_),
    .A2(_12781_),
    .B1(_12784_),
    .C1(_12785_),
    .X(_12786_));
 sky130_fd_sc_hd__o211ai_2 _40187_ (.A1(_12785_),
    .A2(_12784_),
    .B1(_12781_),
    .C1(_10952_),
    .Y(_12787_));
 sky130_fd_sc_hd__o21ai_2 _40188_ (.A1(_07549_),
    .A2(_09541_),
    .B1(_10434_),
    .Y(_12788_));
 sky130_fd_sc_hd__a21oi_1 _40189_ (.A1(_12786_),
    .A2(_12787_),
    .B1(_12788_),
    .Y(_12789_));
 sky130_fd_sc_hd__and3_1 _40190_ (.A(_12788_),
    .B(_12786_),
    .C(_12787_),
    .X(_12791_));
 sky130_fd_sc_hd__o211ai_2 _40191_ (.A1(_12789_),
    .A2(_12791_),
    .B1(_10439_),
    .C1(_10443_),
    .Y(_12792_));
 sky130_fd_sc_hd__a211o_1 _40192_ (.A1(_10439_),
    .A2(_10443_),
    .B1(_12789_),
    .C1(_12791_),
    .X(_12793_));
 sky130_fd_sc_hd__and3_1 _40193_ (.A(_12780_),
    .B(_12792_),
    .C(_12793_),
    .X(_12794_));
 sky130_fd_sc_hd__a21oi_1 _40194_ (.A1(_12793_),
    .A2(_12792_),
    .B1(_12780_),
    .Y(_12795_));
 sky130_fd_sc_hd__or2_1 _40195_ (.A(_12794_),
    .B(_12795_),
    .X(_12796_));
 sky130_fd_sc_hd__inv_2 _40196_ (.A(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__nand2_1 _40197_ (.A(_12759_),
    .B(_12797_),
    .Y(_12798_));
 sky130_fd_sc_hd__o211ai_2 _40198_ (.A1(_12756_),
    .A2(_12758_),
    .B1(_12796_),
    .C1(_11624_),
    .Y(_12799_));
 sky130_fd_sc_hd__a21bo_1 _40199_ (.A1(_10447_),
    .A2(_10473_),
    .B1_N(_10446_),
    .X(_12800_));
 sky130_fd_sc_hd__a21oi_2 _40200_ (.A1(_12798_),
    .A2(_12799_),
    .B1(_12800_),
    .Y(_12802_));
 sky130_fd_sc_hd__and3_1 _40201_ (.A(_12800_),
    .B(_12798_),
    .C(_12799_),
    .X(_12803_));
 sky130_fd_sc_hd__nor2_1 _40202_ (.A(_12802_),
    .B(_12803_),
    .Y(_12804_));
 sky130_fd_sc_hd__nand2_1 _40203_ (.A(_12755_),
    .B(_12804_),
    .Y(_12805_));
 sky130_fd_sc_hd__nand3_2 _40204_ (.A(_12751_),
    .B(_12748_),
    .C(_12750_),
    .Y(_12806_));
 sky130_fd_sc_hd__o22ai_2 _40205_ (.A1(_12745_),
    .A2(_12747_),
    .B1(_12170_),
    .B2(_12172_),
    .Y(_12807_));
 sky130_fd_sc_hd__o211a_1 _40206_ (.A1(_12753_),
    .A2(_11629_),
    .B1(_12806_),
    .C1(_12807_),
    .X(_12808_));
 sky130_fd_sc_hd__nand2_1 _40207_ (.A(_11628_),
    .B(_11633_),
    .Y(_12809_));
 sky130_fd_sc_hd__o211ai_4 _40208_ (.A1(_12753_),
    .A2(_11629_),
    .B1(_12806_),
    .C1(_12807_),
    .Y(_12810_));
 sky130_fd_sc_hd__nand2_1 _40209_ (.A(_12810_),
    .B(_12755_),
    .Y(_12811_));
 sky130_fd_sc_hd__o21ai_1 _40210_ (.A1(_12802_),
    .A2(_12803_),
    .B1(_12811_),
    .Y(_12813_));
 sky130_fd_sc_hd__o211ai_4 _40211_ (.A1(_12805_),
    .A2(_12808_),
    .B1(_12809_),
    .C1(_12813_),
    .Y(_12814_));
 sky130_fd_sc_hd__nand2_1 _40212_ (.A(_12811_),
    .B(_12804_),
    .Y(_12815_));
 sky130_fd_sc_hd__a21boi_2 _40213_ (.A1(_10484_),
    .A2(_11632_),
    .B1_N(_11628_),
    .Y(_12816_));
 sky130_fd_sc_hd__o211ai_4 _40214_ (.A1(_12802_),
    .A2(_12803_),
    .B1(_12810_),
    .C1(_12755_),
    .Y(_12817_));
 sky130_fd_sc_hd__nand3_2 _40215_ (.A(_12815_),
    .B(_12816_),
    .C(_12817_),
    .Y(_12818_));
 sky130_fd_sc_hd__a21bo_1 _40216_ (.A1(_11648_),
    .A2(_11661_),
    .B1_N(_11662_),
    .X(_12819_));
 sky130_fd_sc_hd__and2_1 _40217_ (.A(_25159_),
    .B(_25242_),
    .X(_12820_));
 sky130_fd_sc_hd__or3b_2 _40218_ (.A(_23718_),
    .B(_23724_),
    .C_N(_07497_),
    .X(_12821_));
 sky130_fd_sc_hd__or2_1 _40219_ (.A(_08956_),
    .B(_23725_),
    .X(_12822_));
 sky130_fd_sc_hd__o211a_2 _40220_ (.A1(_12820_),
    .A2(_11650_),
    .B1(_12821_),
    .C1(_12822_),
    .X(_12824_));
 sky130_fd_sc_hd__a221oi_4 _40221_ (.A1(_23595_),
    .A2(_07502_),
    .B1(_12822_),
    .B2(_12821_),
    .C1(_12820_),
    .Y(_12825_));
 sky130_fd_sc_hd__o2bb2a_1 _40222_ (.A1_N(_10296_),
    .A2_N(_10300_),
    .B1(_12824_),
    .B2(_12825_),
    .X(_12826_));
 sky130_fd_sc_hd__and4bb_1 _40223_ (.A_N(_12824_),
    .B_N(_12825_),
    .C(_10296_),
    .D(_10300_),
    .X(_12827_));
 sky130_fd_sc_hd__or3_4 _40224_ (.A(_11652_),
    .B(_12826_),
    .C(_12827_),
    .X(_12828_));
 sky130_fd_sc_hd__o21ai_2 _40225_ (.A1(_12826_),
    .A2(_12827_),
    .B1(_11652_),
    .Y(_12829_));
 sky130_fd_sc_hd__a211o_1 _40226_ (.A1(_12828_),
    .A2(_12829_),
    .B1(_10465_),
    .C1(_10471_),
    .X(_12830_));
 sky130_fd_sc_hd__o211ai_4 _40227_ (.A1(_10465_),
    .A2(_10471_),
    .B1(_12828_),
    .C1(_12829_),
    .Y(_12831_));
 sky130_fd_sc_hd__and3_1 _40228_ (.A(_11652_),
    .B(_11653_),
    .C(_10299_),
    .X(_12832_));
 sky130_fd_sc_hd__a221o_1 _40229_ (.A1(_10369_),
    .A2(_11654_),
    .B1(_12830_),
    .B2(_12831_),
    .C1(_12832_),
    .X(_12833_));
 sky130_fd_sc_hd__o211ai_4 _40230_ (.A1(_12832_),
    .A2(_11656_),
    .B1(_12830_),
    .C1(_12831_),
    .Y(_12835_));
 sky130_fd_sc_hd__and2_1 _40231_ (.A(_12833_),
    .B(_12835_),
    .X(_12836_));
 sky130_fd_sc_hd__or2_1 _40232_ (.A(_12819_),
    .B(_12836_),
    .X(_12837_));
 sky130_fd_sc_hd__nand2_4 _40233_ (.A(_12836_),
    .B(_12819_),
    .Y(_12838_));
 sky130_fd_sc_hd__nand2_2 _40234_ (.A(_12837_),
    .B(_12838_),
    .Y(_12839_));
 sky130_fd_sc_hd__inv_2 _40235_ (.A(_12839_),
    .Y(_12840_));
 sky130_fd_sc_hd__a21oi_1 _40236_ (.A1(_09562_),
    .A2(_10476_),
    .B1(_10474_),
    .Y(_12841_));
 sky130_fd_sc_hd__a21o_1 _40237_ (.A1(_10479_),
    .A2(_10478_),
    .B1(_12841_),
    .X(_12842_));
 sky130_fd_sc_hd__o221a_1 _40238_ (.A1(_10378_),
    .A2(_10380_),
    .B1(_12840_),
    .B2(_12842_),
    .C1(_11664_),
    .X(_12843_));
 sky130_fd_sc_hd__a21o_1 _40239_ (.A1(_10475_),
    .A2(_11635_),
    .B1(_12839_),
    .X(_12844_));
 sky130_fd_sc_hd__nand2_1 _40240_ (.A(_12843_),
    .B(_12844_),
    .Y(_12846_));
 sky130_fd_sc_hd__inv_2 _40241_ (.A(_12846_),
    .Y(_12847_));
 sky130_fd_sc_hd__a211o_1 _40242_ (.A1(_10479_),
    .A2(_10478_),
    .B1(_12840_),
    .C1(_12841_),
    .X(_12848_));
 sky130_fd_sc_hd__a22oi_2 _40243_ (.A1(_11646_),
    .A2(_11664_),
    .B1(_12844_),
    .B2(_12848_),
    .Y(_12849_));
 sky130_fd_sc_hd__o2bb2ai_1 _40244_ (.A1_N(_12814_),
    .A2_N(_12818_),
    .B1(_12847_),
    .B2(_12849_),
    .Y(_12850_));
 sky130_fd_sc_hd__a21oi_1 _40245_ (.A1(_12843_),
    .A2(_12844_),
    .B1(_12849_),
    .Y(_12851_));
 sky130_fd_sc_hd__nand3_1 _40246_ (.A(_12814_),
    .B(_12818_),
    .C(_12851_),
    .Y(_12852_));
 sky130_fd_sc_hd__nand3_2 _40247_ (.A(_11698_),
    .B(_12850_),
    .C(_12852_),
    .Y(_12853_));
 sky130_fd_sc_hd__nand2_1 _40248_ (.A(_12814_),
    .B(_12818_),
    .Y(_12854_));
 sky130_fd_sc_hd__nand2_1 _40249_ (.A(_12854_),
    .B(_12851_),
    .Y(_12855_));
 sky130_fd_sc_hd__a21boi_1 _40250_ (.A1(_11676_),
    .A2(_11644_),
    .B1_N(_11639_),
    .Y(_12857_));
 sky130_fd_sc_hd__a21o_1 _40251_ (.A1(_12843_),
    .A2(_12844_),
    .B1(_12849_),
    .X(_12858_));
 sky130_fd_sc_hd__nand3_1 _40252_ (.A(_12814_),
    .B(_12818_),
    .C(_12858_),
    .Y(_12859_));
 sky130_fd_sc_hd__nand3_2 _40253_ (.A(_12855_),
    .B(_12857_),
    .C(_12859_),
    .Y(_12860_));
 sky130_fd_sc_hd__o2111ai_4 _40254_ (.A1(_10386_),
    .A2(_11666_),
    .B1(_11697_),
    .C1(_12853_),
    .D1(_12860_),
    .Y(_12861_));
 sky130_fd_sc_hd__a31o_1 _40255_ (.A1(_10424_),
    .A2(_11671_),
    .A3(_11672_),
    .B1(_11673_),
    .X(_12862_));
 sky130_fd_sc_hd__nand2_1 _40256_ (.A(_12853_),
    .B(_12860_),
    .Y(_12863_));
 sky130_fd_sc_hd__o21a_1 _40257_ (.A1(_10386_),
    .A2(_11666_),
    .B1(_11697_),
    .X(_12864_));
 sky130_fd_sc_hd__inv_2 _40258_ (.A(_12864_),
    .Y(_12865_));
 sky130_fd_sc_hd__a22oi_4 _40259_ (.A1(_11679_),
    .A2(_12862_),
    .B1(_12863_),
    .B2(_12865_),
    .Y(_12866_));
 sky130_fd_sc_hd__nand2_1 _40260_ (.A(_12863_),
    .B(_12865_),
    .Y(_12868_));
 sky130_fd_sc_hd__a32o_1 _40261_ (.A1(_11675_),
    .A2(_11677_),
    .A3(_11678_),
    .B1(_11683_),
    .B2(_11682_),
    .X(_12869_));
 sky130_fd_sc_hd__a21oi_1 _40262_ (.A1(_12868_),
    .A2(_12861_),
    .B1(_12869_),
    .Y(_12870_));
 sky130_fd_sc_hd__a21oi_4 _40263_ (.A1(_12861_),
    .A2(_12866_),
    .B1(_12870_),
    .Y(_12871_));
 sky130_fd_sc_hd__xnor2_4 _40264_ (.A(_11696_),
    .B(_12871_),
    .Y(_00013_));
 sky130_fd_sc_hd__a21o_1 _40265_ (.A1(_12804_),
    .A2(_12755_),
    .B1(_12808_),
    .X(_12872_));
 sky130_fd_sc_hd__a31o_1 _40266_ (.A1(_12751_),
    .A2(_12748_),
    .A3(_12750_),
    .B1(_12747_),
    .X(_12873_));
 sky130_fd_sc_hd__o21ai_2 _40267_ (.A1(_12618_),
    .A2(_12738_),
    .B1(_12739_),
    .Y(_12874_));
 sky130_fd_sc_hd__buf_2 _40268_ (.A(_10935_),
    .X(_12875_));
 sky130_fd_sc_hd__clkbuf_4 _40269_ (.A(_12875_),
    .X(_12876_));
 sky130_fd_sc_hd__mux2_2 _40270_ (.A0(_02017_),
    .A1(_00397_),
    .S(_12147_),
    .X(_12878_));
 sky130_fd_sc_hd__o21a_1 _40271_ (.A1(_12151_),
    .A2(_12876_),
    .B1(_12878_),
    .X(_12879_));
 sky130_fd_sc_hd__buf_2 _40272_ (.A(_10939_),
    .X(_12880_));
 sky130_fd_sc_hd__buf_2 _40273_ (.A(_12880_),
    .X(_12881_));
 sky130_fd_sc_hd__nand2_1 _40274_ (.A(_06607_),
    .B(_12881_),
    .Y(_12882_));
 sky130_fd_sc_hd__nor2_1 _40275_ (.A(_12882_),
    .B(_12878_),
    .Y(_12883_));
 sky130_fd_sc_hd__o21ai_1 _40276_ (.A1(_12137_),
    .A2(_12135_),
    .B1(_12133_),
    .Y(_12884_));
 sky130_fd_sc_hd__clkbuf_2 _40277_ (.A(_10934_),
    .X(_12885_));
 sky130_fd_sc_hd__nor2_1 _40278_ (.A(_12885_),
    .B(_12124_),
    .Y(_12886_));
 sky130_fd_sc_hd__and2_1 _40279_ (.A(_12099_),
    .B(_12105_),
    .X(_12887_));
 sky130_fd_sc_hd__a22oi_1 _40280_ (.A1(_12116_),
    .A2(_12117_),
    .B1(_12103_),
    .B2(_12099_),
    .Y(_12889_));
 sky130_fd_sc_hd__nand3_1 _40281_ (.A(_09505_),
    .B(_10901_),
    .C(_12111_),
    .Y(_12890_));
 sky130_fd_sc_hd__a2bb2oi_1 _40282_ (.A1_N(_12106_),
    .A2_N(_12887_),
    .B1(_12889_),
    .B2(_12890_),
    .Y(_12891_));
 sky130_fd_sc_hd__a41oi_4 _40283_ (.A1(_08127_),
    .A2(_10903_),
    .A3(_10908_),
    .A4(_12109_),
    .B1(_12891_),
    .Y(_12892_));
 sky130_fd_sc_hd__o21ai_4 _40284_ (.A1(_11952_),
    .A2(_11949_),
    .B1(_12069_),
    .Y(_12893_));
 sky130_fd_sc_hd__o21ai_1 _40285_ (.A1(_11872_),
    .A2(_11868_),
    .B1(_11874_),
    .Y(_12894_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40286_ (.A(_10598_),
    .X(_12895_));
 sky130_fd_sc_hd__clkbuf_2 _40287_ (.A(_12895_),
    .X(_12896_));
 sky130_fd_sc_hd__buf_2 _40288_ (.A(_10628_),
    .X(_12897_));
 sky130_fd_sc_hd__nand2_1 _40289_ (.A(_11823_),
    .B(_11825_),
    .Y(_12898_));
 sky130_fd_sc_hd__buf_1 _40290_ (.A(net409),
    .X(_12900_));
 sky130_fd_sc_hd__and3b_1 _40291_ (.A_N(_06233_),
    .B(_12900_),
    .C(_09247_),
    .X(_12901_));
 sky130_fd_sc_hd__a22oi_1 _40292_ (.A1(_12901_),
    .A2(_11819_),
    .B1(_10584_),
    .B2(_10585_),
    .Y(_12902_));
 sky130_fd_sc_hd__o22ai_1 _40293_ (.A1(_10570_),
    .A2(_12898_),
    .B1(_11829_),
    .B2(_12902_),
    .Y(_12903_));
 sky130_fd_sc_hd__a21oi_1 _40294_ (.A1(_11824_),
    .A2(_11827_),
    .B1(_12900_),
    .Y(_12904_));
 sky130_fd_sc_hd__and3_1 _40295_ (.A(_12900_),
    .B(\delay_line[11][15] ),
    .C(_11827_),
    .X(_12905_));
 sky130_fd_sc_hd__nor2_2 _40296_ (.A(_12904_),
    .B(_12905_),
    .Y(_12906_));
 sky130_fd_sc_hd__inv_2 _40297_ (.A(_12906_),
    .Y(_12907_));
 sky130_fd_sc_hd__nand2_1 _40298_ (.A(_12903_),
    .B(_12907_),
    .Y(_12908_));
 sky130_fd_sc_hd__o211ai_2 _40299_ (.A1(_10570_),
    .A2(_12898_),
    .B1(_12906_),
    .C1(_11841_),
    .Y(_12909_));
 sky130_fd_sc_hd__nand2_1 _40300_ (.A(_12908_),
    .B(_12909_),
    .Y(_12911_));
 sky130_fd_sc_hd__nand2_1 _40301_ (.A(_11814_),
    .B(_11813_),
    .Y(_12912_));
 sky130_fd_sc_hd__a221o_2 _40302_ (.A1(_11835_),
    .A2(_10552_),
    .B1(_11807_),
    .B2(_10561_),
    .C1(_12912_),
    .X(_12913_));
 sky130_fd_sc_hd__o22a_1 _40303_ (.A1(_10557_),
    .A2(_11835_),
    .B1(_12913_),
    .B2(_11837_),
    .X(_12914_));
 sky130_fd_sc_hd__nand2_2 _40304_ (.A(_12911_),
    .B(_12914_),
    .Y(_12915_));
 sky130_fd_sc_hd__nor2_1 _40305_ (.A(_11835_),
    .B(_10557_),
    .Y(_12916_));
 sky130_fd_sc_hd__a21oi_2 _40306_ (.A1(_09245_),
    .A2(_11807_),
    .B1(_12913_),
    .Y(_12917_));
 sky130_fd_sc_hd__buf_6 _40307_ (.A(_12909_),
    .X(_12918_));
 sky130_fd_sc_hd__o211ai_4 _40308_ (.A1(_12916_),
    .A2(_12917_),
    .B1(_12908_),
    .C1(_12918_),
    .Y(_12919_));
 sky130_fd_sc_hd__o21ai_2 _40309_ (.A1(_11818_),
    .A2(_11834_),
    .B1(_11858_),
    .Y(_12920_));
 sky130_fd_sc_hd__a22oi_4 _40310_ (.A1(_12915_),
    .A2(_12919_),
    .B1(_12920_),
    .B2(_11852_),
    .Y(_12922_));
 sky130_fd_sc_hd__clkbuf_2 _40311_ (.A(_12919_),
    .X(_12923_));
 sky130_fd_sc_hd__nand3_1 _40312_ (.A(_11852_),
    .B(_12915_),
    .C(_12923_),
    .Y(_12924_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40313_ (.A(_11801_),
    .X(_12925_));
 sky130_fd_sc_hd__a31oi_1 _40314_ (.A1(_11849_),
    .A2(_11850_),
    .A3(_11832_),
    .B1(_12925_),
    .Y(_12926_));
 sky130_fd_sc_hd__a21oi_1 _40315_ (.A1(_11852_),
    .A2(_11851_),
    .B1(_11858_),
    .Y(_12927_));
 sky130_fd_sc_hd__a21oi_1 _40316_ (.A1(_11806_),
    .A2(_11846_),
    .B1(_11845_),
    .Y(_12928_));
 sky130_fd_sc_hd__o22ai_1 _40317_ (.A1(_12924_),
    .A2(_12926_),
    .B1(_12927_),
    .B2(_12928_),
    .Y(_12929_));
 sky130_fd_sc_hd__nand2_1 _40318_ (.A(_11838_),
    .B(_11839_),
    .Y(_12930_));
 sky130_fd_sc_hd__o2111a_1 _40319_ (.A1(_11849_),
    .A2(_12930_),
    .B1(_12915_),
    .C1(_12923_),
    .D1(_12920_),
    .X(_12931_));
 sky130_fd_sc_hd__o21a_1 _40320_ (.A1(_11818_),
    .A2(_11834_),
    .B1(_11852_),
    .X(_12933_));
 sky130_fd_sc_hd__nand2_1 _40321_ (.A(_11806_),
    .B(_11846_),
    .Y(_12934_));
 sky130_fd_sc_hd__a21oi_2 _40322_ (.A1(_12933_),
    .A2(_12934_),
    .B1(_12927_),
    .Y(_12935_));
 sky130_fd_sc_hd__o21ai_2 _40323_ (.A1(_12922_),
    .A2(_12931_),
    .B1(_12935_),
    .Y(_12936_));
 sky130_fd_sc_hd__o21ai_1 _40324_ (.A1(_12922_),
    .A2(_12929_),
    .B1(_12936_),
    .Y(_12937_));
 sky130_fd_sc_hd__o21ai_1 _40325_ (.A1(_12896_),
    .A2(_12897_),
    .B1(_12937_),
    .Y(_12938_));
 sky130_fd_sc_hd__a21oi_1 _40326_ (.A1(_11863_),
    .A2(_11864_),
    .B1(_11857_),
    .Y(_12939_));
 sky130_fd_sc_hd__o2111ai_1 _40327_ (.A1(_12922_),
    .A2(_12929_),
    .B1(_12936_),
    .C1(_10545_),
    .D1(_12925_),
    .Y(_12940_));
 sky130_fd_sc_hd__nand3_2 _40328_ (.A(_12938_),
    .B(_12939_),
    .C(_12940_),
    .Y(_12941_));
 sky130_fd_sc_hd__a21oi_1 _40329_ (.A1(_11850_),
    .A2(_11832_),
    .B1(_11849_),
    .Y(_12942_));
 sky130_fd_sc_hd__clkbuf_2 _40330_ (.A(_12915_),
    .X(_12944_));
 sky130_fd_sc_hd__nand2_1 _40331_ (.A(_12944_),
    .B(_12923_),
    .Y(_12945_));
 sky130_fd_sc_hd__o21ai_1 _40332_ (.A1(_12942_),
    .A2(_12926_),
    .B1(_12945_),
    .Y(_12946_));
 sky130_fd_sc_hd__o2111ai_2 _40333_ (.A1(_11849_),
    .A2(_12930_),
    .B1(_12944_),
    .C1(_12923_),
    .D1(_12920_),
    .Y(_12947_));
 sky130_fd_sc_hd__nand2_1 _40334_ (.A(_12946_),
    .B(_12947_),
    .Y(_12948_));
 sky130_fd_sc_hd__o22ai_4 _40335_ (.A1(_12896_),
    .A2(_12897_),
    .B1(_12935_),
    .B2(_12948_),
    .Y(_12949_));
 sky130_fd_sc_hd__o21a_1 _40336_ (.A1(_12922_),
    .A2(_12931_),
    .B1(_12935_),
    .X(_12950_));
 sky130_fd_sc_hd__a21o_1 _40337_ (.A1(_11863_),
    .A2(_11864_),
    .B1(_11857_),
    .X(_12951_));
 sky130_fd_sc_hd__nor2_2 _40338_ (.A(_12896_),
    .B(_10628_),
    .Y(_12952_));
 sky130_fd_sc_hd__nand2_1 _40339_ (.A(_12937_),
    .B(_12952_),
    .Y(_12953_));
 sky130_fd_sc_hd__o211ai_4 _40340_ (.A1(_12949_),
    .A2(_12950_),
    .B1(_12951_),
    .C1(_12953_),
    .Y(_12955_));
 sky130_fd_sc_hd__inv_2 _40341_ (.A(_06287_),
    .Y(_12956_));
 sky130_fd_sc_hd__nand2_1 _40342_ (.A(_12956_),
    .B(_10545_),
    .Y(_12957_));
 sky130_fd_sc_hd__nand2_1 _40343_ (.A(_10640_),
    .B(_10541_),
    .Y(_12958_));
 sky130_fd_sc_hd__o2bb2a_1 _40344_ (.A1_N(_12957_),
    .A2_N(_12958_),
    .B1(_12895_),
    .B2(_10543_),
    .X(_12959_));
 sky130_fd_sc_hd__a211oi_2 _40345_ (.A1(_12956_),
    .A2(_11802_),
    .B1(_11795_),
    .C1(_12959_),
    .Y(_12960_));
 sky130_fd_sc_hd__buf_1 _40346_ (.A(_04775_),
    .X(_12961_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40347_ (.A(_12897_),
    .X(_12962_));
 sky130_fd_sc_hd__and4_1 _40348_ (.A(_12956_),
    .B(_12925_),
    .C(_10628_),
    .D(_10607_),
    .X(_12963_));
 sky130_fd_sc_hd__o2bb2a_1 _40349_ (.A1_N(_12961_),
    .A2_N(_12962_),
    .B1(_12963_),
    .B2(_12959_),
    .X(_12964_));
 sky130_fd_sc_hd__o2bb2ai_1 _40350_ (.A1_N(_12941_),
    .A2_N(_12955_),
    .B1(_12960_),
    .B2(_12964_),
    .Y(_12966_));
 sky130_fd_sc_hd__a211oi_1 _40351_ (.A1(_12961_),
    .A2(_12962_),
    .B1(_12963_),
    .C1(_12959_),
    .Y(_12967_));
 sky130_fd_sc_hd__o211a_1 _40352_ (.A1(_12963_),
    .A2(_12959_),
    .B1(_12961_),
    .C1(_12962_),
    .X(_12968_));
 sky130_fd_sc_hd__o211ai_1 _40353_ (.A1(_12967_),
    .A2(_12968_),
    .B1(_12941_),
    .C1(_12955_),
    .Y(_12969_));
 sky130_fd_sc_hd__nand3_1 _40354_ (.A(_12894_),
    .B(_12966_),
    .C(_12969_),
    .Y(_12970_));
 sky130_fd_sc_hd__o21a_1 _40355_ (.A1(_11872_),
    .A2(_11868_),
    .B1(_11874_),
    .X(_12971_));
 sky130_fd_sc_hd__o211ai_1 _40356_ (.A1(_12960_),
    .A2(_12964_),
    .B1(_12941_),
    .C1(_12955_),
    .Y(_12972_));
 sky130_fd_sc_hd__o2bb2ai_1 _40357_ (.A1_N(_12941_),
    .A2_N(_12955_),
    .B1(_12967_),
    .B2(_12968_),
    .Y(_12973_));
 sky130_fd_sc_hd__nand3_2 _40358_ (.A(_12971_),
    .B(_12972_),
    .C(_12973_),
    .Y(_12974_));
 sky130_fd_sc_hd__o21ai_2 _40359_ (.A1(_11793_),
    .A2(_11798_),
    .B1(_11797_),
    .Y(_12975_));
 sky130_fd_sc_hd__o21a_1 _40360_ (.A1(_11797_),
    .A2(_11793_),
    .B1(_12975_),
    .X(_12977_));
 sky130_fd_sc_hd__and3_1 _40361_ (.A(_04789_),
    .B(_11883_),
    .C(_12977_),
    .X(_12978_));
 sky130_fd_sc_hd__a21oi_2 _40362_ (.A1(_04789_),
    .A2(_11883_),
    .B1(_12977_),
    .Y(_12979_));
 sky130_fd_sc_hd__nor2_1 _40363_ (.A(_12978_),
    .B(_12979_),
    .Y(_12980_));
 sky130_fd_sc_hd__a21bo_1 _40364_ (.A1(_12970_),
    .A2(_12974_),
    .B1_N(_12980_),
    .X(_12981_));
 sky130_fd_sc_hd__nor2_1 _40365_ (.A(_11893_),
    .B(_11894_),
    .Y(_12982_));
 sky130_fd_sc_hd__inv_2 _40366_ (.A(_12982_),
    .Y(_12983_));
 sky130_fd_sc_hd__a32oi_4 _40367_ (.A1(_11792_),
    .A2(_11871_),
    .A3(_11875_),
    .B1(_11882_),
    .B2(_12983_),
    .Y(_12984_));
 sky130_fd_sc_hd__clkbuf_2 _40368_ (.A(_12970_),
    .X(_12985_));
 sky130_fd_sc_hd__o211ai_2 _40369_ (.A1(_12978_),
    .A2(_12979_),
    .B1(_12985_),
    .C1(_12974_),
    .Y(_12986_));
 sky130_fd_sc_hd__nand3_4 _40370_ (.A(_12981_),
    .B(_12984_),
    .C(_12986_),
    .Y(_12988_));
 sky130_fd_sc_hd__a32o_1 _40371_ (.A1(_11792_),
    .A2(_11871_),
    .A3(_11875_),
    .B1(_11882_),
    .B2(_12983_),
    .X(_12989_));
 sky130_fd_sc_hd__nand3_2 _40372_ (.A(_12985_),
    .B(_12974_),
    .C(_12980_),
    .Y(_12990_));
 sky130_fd_sc_hd__o2bb2ai_2 _40373_ (.A1_N(_12985_),
    .A2_N(_12974_),
    .B1(_12978_),
    .B2(_12979_),
    .Y(_12991_));
 sky130_fd_sc_hd__nand3_2 _40374_ (.A(_12989_),
    .B(_12990_),
    .C(_12991_),
    .Y(_12992_));
 sky130_fd_sc_hd__clkbuf_2 _40375_ (.A(_10502_),
    .X(_12993_));
 sky130_fd_sc_hd__clkbuf_2 _40376_ (.A(_04800_),
    .X(_12994_));
 sky130_fd_sc_hd__a311oi_2 _40377_ (.A1(_10507_),
    .A2(_06200_),
    .A3(_12993_),
    .B1(_10644_),
    .C1(_12994_),
    .Y(_12995_));
 sky130_fd_sc_hd__o2111a_1 _40378_ (.A1(_10499_),
    .A2(_12994_),
    .B1(_06200_),
    .C1(_10507_),
    .D1(_12993_),
    .X(_12996_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40379_ (.A(_10502_),
    .X(_12997_));
 sky130_fd_sc_hd__a21o_1 _40380_ (.A1(_10507_),
    .A2(_12997_),
    .B1(_03125_),
    .X(_12999_));
 sky130_fd_sc_hd__o211a_1 _40381_ (.A1(_12995_),
    .A2(_12996_),
    .B1(_11908_),
    .C1(_12999_),
    .X(_13000_));
 sky130_fd_sc_hd__a211oi_2 _40382_ (.A1(_11908_),
    .A2(_12999_),
    .B1(_12995_),
    .C1(_12996_),
    .Y(_13001_));
 sky130_fd_sc_hd__or2_1 _40383_ (.A(_07867_),
    .B(_07870_),
    .X(_13002_));
 sky130_fd_sc_hd__nand2_1 _40384_ (.A(_07870_),
    .B(_07867_),
    .Y(_13003_));
 sky130_fd_sc_hd__and4_1 _40385_ (.A(_13002_),
    .B(_13003_),
    .C(_07863_),
    .D(_10526_),
    .X(_13004_));
 sky130_fd_sc_hd__inv_2 _40386_ (.A(_13004_),
    .Y(_13005_));
 sky130_fd_sc_hd__buf_1 _40387_ (.A(_07863_),
    .X(_13006_));
 sky130_fd_sc_hd__a22o_1 _40388_ (.A1(_13006_),
    .A2(_10526_),
    .B1(_13002_),
    .B2(_13003_),
    .X(_13007_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40389_ (.A(_07878_),
    .X(_13008_));
 sky130_fd_sc_hd__nor2_1 _40390_ (.A(_01702_),
    .B(_13008_),
    .Y(_13010_));
 sky130_fd_sc_hd__and3_2 _40391_ (.A(_13005_),
    .B(_13007_),
    .C(_13010_),
    .X(_13011_));
 sky130_fd_sc_hd__o2bb2a_1 _40392_ (.A1_N(_13005_),
    .A2_N(_13007_),
    .B1(_01702_),
    .B2(_13008_),
    .X(_13012_));
 sky130_fd_sc_hd__nand2_1 _40393_ (.A(_13006_),
    .B(_12993_),
    .Y(_13013_));
 sky130_fd_sc_hd__or2b_2 _40394_ (.A(_10502_),
    .B_N(_10527_),
    .X(_13014_));
 sky130_fd_sc_hd__o211a_1 _40395_ (.A1(_13011_),
    .A2(_13012_),
    .B1(_13013_),
    .C1(_13014_),
    .X(_13015_));
 sky130_fd_sc_hd__a211oi_4 _40396_ (.A1(_13013_),
    .A2(_13014_),
    .B1(_13011_),
    .C1(_13012_),
    .Y(_13016_));
 sky130_fd_sc_hd__o22ai_4 _40397_ (.A1(_13000_),
    .A2(_13001_),
    .B1(_13015_),
    .B2(_13016_),
    .Y(_13017_));
 sky130_fd_sc_hd__or4_2 _40398_ (.A(_13000_),
    .B(_13001_),
    .C(_13015_),
    .D(_13016_),
    .X(_13018_));
 sky130_fd_sc_hd__a221o_1 _40399_ (.A1(_10647_),
    .A2(_11889_),
    .B1(_13017_),
    .B2(_13018_),
    .C1(_11887_),
    .X(_13019_));
 sky130_fd_sc_hd__o211ai_4 _40400_ (.A1(_11887_),
    .A2(_11890_),
    .B1(_13017_),
    .C1(_13018_),
    .Y(_13021_));
 sky130_fd_sc_hd__and2_1 _40401_ (.A(_13019_),
    .B(_13021_),
    .X(_13022_));
 sky130_fd_sc_hd__a21o_1 _40402_ (.A1(_11912_),
    .A2(_11927_),
    .B1(_11906_),
    .X(_13023_));
 sky130_fd_sc_hd__nand2_1 _40403_ (.A(_13022_),
    .B(_13023_),
    .Y(_13024_));
 sky130_fd_sc_hd__a211o_1 _40404_ (.A1(_11912_),
    .A2(_11927_),
    .B1(_13022_),
    .C1(_11906_),
    .X(_13025_));
 sky130_fd_sc_hd__and2_2 _40405_ (.A(_13024_),
    .B(_13025_),
    .X(_13026_));
 sky130_fd_sc_hd__inv_2 _40406_ (.A(_13026_),
    .Y(_13027_));
 sky130_fd_sc_hd__a21o_1 _40407_ (.A1(_12988_),
    .A2(_12992_),
    .B1(_13027_),
    .X(_13028_));
 sky130_fd_sc_hd__a32oi_4 _40408_ (.A1(_11791_),
    .A2(_11892_),
    .A3(_11895_),
    .B1(_11902_),
    .B2(_11935_),
    .Y(_13029_));
 sky130_fd_sc_hd__nand3_1 _40409_ (.A(_13027_),
    .B(_12988_),
    .C(_12992_),
    .Y(_13030_));
 sky130_fd_sc_hd__nand3_4 _40410_ (.A(_13028_),
    .B(_13029_),
    .C(_13030_),
    .Y(_13032_));
 sky130_fd_sc_hd__a32o_1 _40411_ (.A1(_11791_),
    .A2(_11892_),
    .A3(_11895_),
    .B1(_11902_),
    .B2(_11935_),
    .X(_13033_));
 sky130_fd_sc_hd__a21o_1 _40412_ (.A1(_12988_),
    .A2(_12992_),
    .B1(_13026_),
    .X(_13034_));
 sky130_fd_sc_hd__nand3_2 _40413_ (.A(_12988_),
    .B(_12992_),
    .C(_13026_),
    .Y(_13035_));
 sky130_fd_sc_hd__nand3_4 _40414_ (.A(_13033_),
    .B(_13034_),
    .C(_13035_),
    .Y(_13036_));
 sky130_fd_sc_hd__a21boi_1 _40415_ (.A1(_11763_),
    .A2(_11782_),
    .B1_N(_11783_),
    .Y(_13037_));
 sky130_fd_sc_hd__o211ai_1 _40416_ (.A1(_01793_),
    .A2(_11757_),
    .B1(_11758_),
    .C1(_11752_),
    .Y(_13038_));
 sky130_fd_sc_hd__nand3_1 _40417_ (.A(_07703_),
    .B(_03322_),
    .C(_11749_),
    .Y(_13039_));
 sky130_fd_sc_hd__or2_1 _40418_ (.A(_11751_),
    .B(_13039_),
    .X(_13040_));
 sky130_fd_sc_hd__buf_1 _40419_ (.A(_11753_),
    .X(_13041_));
 sky130_fd_sc_hd__a31o_1 _40420_ (.A1(_07703_),
    .A2(_03322_),
    .A3(_13041_),
    .B1(_07690_),
    .X(_13043_));
 sky130_fd_sc_hd__or2_1 _40421_ (.A(_10705_),
    .B(_13039_),
    .X(_13044_));
 sky130_fd_sc_hd__clkbuf_2 _40422_ (.A(_07675_),
    .X(_13045_));
 sky130_fd_sc_hd__a21oi_1 _40423_ (.A1(_13043_),
    .A2(_13044_),
    .B1(_13045_),
    .Y(_13046_));
 sky130_fd_sc_hd__and3_1 _40424_ (.A(_13044_),
    .B(_13045_),
    .C(_13043_),
    .X(_13047_));
 sky130_fd_sc_hd__a211oi_1 _40425_ (.A1(_13038_),
    .A2(_13040_),
    .B1(_13046_),
    .C1(_13047_),
    .Y(_13048_));
 sky130_fd_sc_hd__o221a_1 _40426_ (.A1(_13039_),
    .A2(_11751_),
    .B1(_13046_),
    .B2(_13047_),
    .C1(_13038_),
    .X(_13049_));
 sky130_fd_sc_hd__buf_1 _40427_ (.A(_09148_),
    .X(_13050_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40428_ (.A(_13050_),
    .X(_13051_));
 sky130_fd_sc_hd__nand2_1 _40429_ (.A(_09125_),
    .B(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__a21oi_1 _40430_ (.A1(_09125_),
    .A2(_11738_),
    .B1(_03347_),
    .Y(_13054_));
 sky130_fd_sc_hd__and3_1 _40431_ (.A(_09124_),
    .B(_03347_),
    .C(_09148_),
    .X(_13055_));
 sky130_fd_sc_hd__or3_1 _40432_ (.A(_11748_),
    .B(_13054_),
    .C(_13055_),
    .X(_13056_));
 sky130_fd_sc_hd__o21ai_2 _40433_ (.A1(_13054_),
    .A2(_13055_),
    .B1(_11748_),
    .Y(_13057_));
 sky130_fd_sc_hd__nand2_1 _40434_ (.A(_13056_),
    .B(_13057_),
    .Y(_13058_));
 sky130_fd_sc_hd__or3_1 _40435_ (.A(_11737_),
    .B(_13052_),
    .C(_13058_),
    .X(_13059_));
 sky130_fd_sc_hd__clkbuf_2 _40436_ (.A(_13050_),
    .X(_13060_));
 sky130_fd_sc_hd__a32o_1 _40437_ (.A1(_03354_),
    .A2(_09125_),
    .A3(_13060_),
    .B1(_13056_),
    .B2(_13057_),
    .X(_13061_));
 sky130_fd_sc_hd__nand2_1 _40438_ (.A(_13059_),
    .B(_13061_),
    .Y(_13062_));
 sky130_fd_sc_hd__or2_1 _40439_ (.A(_13049_),
    .B(_13062_),
    .X(_13063_));
 sky130_fd_sc_hd__o21ai_1 _40440_ (.A1(_13048_),
    .A2(_13049_),
    .B1(_13062_),
    .Y(_13065_));
 sky130_fd_sc_hd__o21a_1 _40441_ (.A1(_13048_),
    .A2(_13063_),
    .B1(_13065_),
    .X(_13066_));
 sky130_fd_sc_hd__nand2_1 _40442_ (.A(_11776_),
    .B(_11765_),
    .Y(_13067_));
 sky130_fd_sc_hd__nor2_1 _40443_ (.A(_11919_),
    .B(_11920_),
    .Y(_13068_));
 sky130_fd_sc_hd__a31o_1 _40444_ (.A1(_10502_),
    .A2(_10520_),
    .A3(_13068_),
    .B1(_11926_),
    .X(_13069_));
 sky130_fd_sc_hd__and3_1 _40445_ (.A(_11913_),
    .B(_11914_),
    .C(_10519_),
    .X(_13070_));
 sky130_fd_sc_hd__nor2_1 _40446_ (.A(_07697_),
    .B(_07698_),
    .Y(_13071_));
 sky130_fd_sc_hd__a31o_1 _40447_ (.A1(_11915_),
    .A2(_10511_),
    .A3(_11916_),
    .B1(_13071_),
    .X(_13072_));
 sky130_fd_sc_hd__o21ai_2 _40448_ (.A1(_13070_),
    .A2(_11917_),
    .B1(_13071_),
    .Y(_13073_));
 sky130_fd_sc_hd__o21a_1 _40449_ (.A1(_13070_),
    .A2(_13072_),
    .B1(_13073_),
    .X(_13074_));
 sky130_fd_sc_hd__nand2_1 _40450_ (.A(_11770_),
    .B(_13074_),
    .Y(_13076_));
 sky130_fd_sc_hd__a21o_1 _40451_ (.A1(_11768_),
    .A2(_11772_),
    .B1(_13074_),
    .X(_13077_));
 sky130_fd_sc_hd__and3_1 _40452_ (.A(_13069_),
    .B(_13076_),
    .C(_13077_),
    .X(_13078_));
 sky130_fd_sc_hd__a21o_1 _40453_ (.A1(_13076_),
    .A2(_13077_),
    .B1(_13069_),
    .X(_13079_));
 sky130_fd_sc_hd__or2b_1 _40454_ (.A(_13078_),
    .B_N(_13079_),
    .X(_13080_));
 sky130_fd_sc_hd__a21oi_1 _40455_ (.A1(_11771_),
    .A2(_11774_),
    .B1(_13080_),
    .Y(_13081_));
 sky130_fd_sc_hd__nand2_1 _40456_ (.A(_11773_),
    .B(_11771_),
    .Y(_13082_));
 sky130_fd_sc_hd__o311a_1 _40457_ (.A1(_07690_),
    .A2(_13008_),
    .A3(_13082_),
    .B1(_13080_),
    .C1(_11771_),
    .X(_13083_));
 sky130_fd_sc_hd__or2_1 _40458_ (.A(_13081_),
    .B(_13083_),
    .X(_13084_));
 sky130_fd_sc_hd__a21oi_1 _40459_ (.A1(_13067_),
    .A2(_11780_),
    .B1(_13084_),
    .Y(_13085_));
 sky130_fd_sc_hd__and3_1 _40460_ (.A(_13067_),
    .B(_11780_),
    .C(_13084_),
    .X(_13087_));
 sky130_fd_sc_hd__nor2_1 _40461_ (.A(_13085_),
    .B(_13087_),
    .Y(_13088_));
 sky130_fd_sc_hd__xnor2_1 _40462_ (.A(_13066_),
    .B(_13088_),
    .Y(_13089_));
 sky130_fd_sc_hd__nand3_1 _40463_ (.A(_11930_),
    .B(_11944_),
    .C(_13089_),
    .Y(_13090_));
 sky130_fd_sc_hd__a21o_1 _40464_ (.A1(_11930_),
    .A2(_11944_),
    .B1(_13089_),
    .X(_13091_));
 sky130_fd_sc_hd__nand2_1 _40465_ (.A(_13090_),
    .B(_13091_),
    .Y(_13092_));
 sky130_fd_sc_hd__or2_1 _40466_ (.A(_13037_),
    .B(_13092_),
    .X(_13093_));
 sky130_fd_sc_hd__nand2_1 _40467_ (.A(_13092_),
    .B(_13037_),
    .Y(_13094_));
 sky130_fd_sc_hd__nand2_1 _40468_ (.A(_13093_),
    .B(_13094_),
    .Y(_13095_));
 sky130_fd_sc_hd__inv_2 _40469_ (.A(_13095_),
    .Y(_13096_));
 sky130_fd_sc_hd__a21o_2 _40470_ (.A1(_13032_),
    .A2(_13036_),
    .B1(_13096_),
    .X(_13098_));
 sky130_fd_sc_hd__nand3_4 _40471_ (.A(_13036_),
    .B(_13096_),
    .C(_13032_),
    .Y(_13099_));
 sky130_fd_sc_hd__nand3_2 _40472_ (.A(_12893_),
    .B(_13098_),
    .C(_13099_),
    .Y(_13100_));
 sky130_fd_sc_hd__o21ba_1 _40473_ (.A1(_12052_),
    .A2(_12000_),
    .B1_N(_11997_),
    .X(_13101_));
 sky130_fd_sc_hd__nand2_1 _40474_ (.A(_12033_),
    .B(_12011_),
    .Y(_13102_));
 sky130_fd_sc_hd__or2_1 _40475_ (.A(_12006_),
    .B(_13102_),
    .X(_13103_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40476_ (.A(_10849_),
    .X(_13104_));
 sky130_fd_sc_hd__clkbuf_2 _40477_ (.A(_12013_),
    .X(_13105_));
 sky130_fd_sc_hd__nor2_1 _40478_ (.A(_13104_),
    .B(_13105_),
    .Y(_13106_));
 sky130_fd_sc_hd__a211oi_1 _40479_ (.A1(_12036_),
    .A2(_12038_),
    .B1(_10747_),
    .C1(_13106_),
    .Y(_13107_));
 sky130_fd_sc_hd__o221a_1 _40480_ (.A1(_09391_),
    .A2(_13105_),
    .B1(_10747_),
    .B2(_13106_),
    .C1(_12038_),
    .X(_13109_));
 sky130_fd_sc_hd__a211oi_1 _40481_ (.A1(_12040_),
    .A2(_13103_),
    .B1(_13107_),
    .C1(_13109_),
    .Y(_13110_));
 sky130_fd_sc_hd__o221a_1 _40482_ (.A1(_13102_),
    .A2(_12006_),
    .B1(_13109_),
    .B2(_13107_),
    .C1(_12040_),
    .X(_13111_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40483_ (.A(_12012_),
    .X(_13112_));
 sky130_fd_sc_hd__clkbuf_2 _40484_ (.A(_12015_),
    .X(_13113_));
 sky130_fd_sc_hd__and4b_1 _40485_ (.A_N(_03457_),
    .B(_13113_),
    .C(_13104_),
    .D(_12004_),
    .X(_13114_));
 sky130_fd_sc_hd__a31oi_1 _40486_ (.A1(_13112_),
    .A2(_10749_),
    .A3(_12014_),
    .B1(_13114_),
    .Y(_13115_));
 sky130_fd_sc_hd__or3b_1 _40487_ (.A(_13110_),
    .B(_13111_),
    .C_N(_13115_),
    .X(_13116_));
 sky130_fd_sc_hd__o21bai_1 _40488_ (.A1(_13110_),
    .A2(_13111_),
    .B1_N(_13115_),
    .Y(_13117_));
 sky130_fd_sc_hd__nand2_1 _40489_ (.A(_13116_),
    .B(_13117_),
    .Y(_13118_));
 sky130_fd_sc_hd__nor3_1 _40490_ (.A(_12032_),
    .B(_12043_),
    .C(_12045_),
    .Y(_13120_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40491_ (.A(_08010_),
    .X(_13121_));
 sky130_fd_sc_hd__and3b_1 _40492_ (.A_N(_12033_),
    .B(_13121_),
    .C(_12012_),
    .X(_13122_));
 sky130_fd_sc_hd__mux2_1 _40493_ (.A0(_13102_),
    .A1(_12003_),
    .S(_13121_),
    .X(_13123_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40494_ (.A(_06157_),
    .X(_13124_));
 sky130_fd_sc_hd__nor2_2 _40495_ (.A(_13124_),
    .B(_12015_),
    .Y(_13125_));
 sky130_fd_sc_hd__and2_1 _40496_ (.A(_13124_),
    .B(_12015_),
    .X(_13126_));
 sky130_fd_sc_hd__or3_1 _40497_ (.A(_12003_),
    .B(_13125_),
    .C(_13126_),
    .X(_13127_));
 sky130_fd_sc_hd__o21ai_2 _40498_ (.A1(_13125_),
    .A2(_13126_),
    .B1(_12012_),
    .Y(_13128_));
 sky130_fd_sc_hd__nand3_1 _40499_ (.A(_13123_),
    .B(_13127_),
    .C(_13128_),
    .Y(_13129_));
 sky130_fd_sc_hd__nand3b_1 _40500_ (.A_N(_12033_),
    .B(_13121_),
    .C(_12012_),
    .Y(_13131_));
 sky130_fd_sc_hd__a22o_1 _40501_ (.A1(_13131_),
    .A2(_13123_),
    .B1(_13127_),
    .B2(_13128_),
    .X(_13132_));
 sky130_fd_sc_hd__o21a_1 _40502_ (.A1(_13122_),
    .A2(_13129_),
    .B1(_13132_),
    .X(_13133_));
 sky130_fd_sc_hd__buf_1 _40503_ (.A(_12029_),
    .X(_13134_));
 sky130_fd_sc_hd__buf_1 _40504_ (.A(_13134_),
    .X(_13135_));
 sky130_fd_sc_hd__o21ai_2 _40505_ (.A1(_11977_),
    .A2(net246),
    .B1(_13134_),
    .Y(_13136_));
 sky130_fd_sc_hd__o21ai_1 _40506_ (.A1(_13135_),
    .A2(_11977_),
    .B1(_13136_),
    .Y(_13137_));
 sky130_fd_sc_hd__and2_1 _40507_ (.A(_12030_),
    .B(_13137_),
    .X(_13138_));
 sky130_fd_sc_hd__buf_1 _40508_ (.A(_12025_),
    .X(_13139_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40509_ (.A(_13134_),
    .X(_13140_));
 sky130_fd_sc_hd__o2111a_1 _40510_ (.A1(_10796_),
    .A2(net223),
    .B1(_13139_),
    .C1(_13140_),
    .D1(_13136_),
    .X(_13142_));
 sky130_fd_sc_hd__nor2_1 _40511_ (.A(_13138_),
    .B(_13142_),
    .Y(_13143_));
 sky130_fd_sc_hd__nand2_1 _40512_ (.A(_13133_),
    .B(_13143_),
    .Y(_13144_));
 sky130_fd_sc_hd__or2_1 _40513_ (.A(_13133_),
    .B(_13143_),
    .X(_13145_));
 sky130_fd_sc_hd__o211a_1 _40514_ (.A1(_12032_),
    .A2(_13120_),
    .B1(_13144_),
    .C1(_13145_),
    .X(_13146_));
 sky130_fd_sc_hd__a211o_1 _40515_ (.A1(_13144_),
    .A2(_13145_),
    .B1(_12032_),
    .C1(_13120_),
    .X(_13147_));
 sky130_fd_sc_hd__and2b_1 _40516_ (.A_N(_13146_),
    .B(_13147_),
    .X(_13148_));
 sky130_fd_sc_hd__xnor2_2 _40517_ (.A(_13118_),
    .B(_13148_),
    .Y(_13149_));
 sky130_fd_sc_hd__o31ai_2 _40518_ (.A1(_11744_),
    .A2(net189),
    .A3(_11762_),
    .B1(_11760_),
    .Y(_13150_));
 sky130_fd_sc_hd__nor2_1 _40519_ (.A(_01745_),
    .B(_09355_),
    .Y(_13151_));
 sky130_fd_sc_hd__and2_1 _40520_ (.A(_06091_),
    .B(_01745_),
    .X(_13153_));
 sky130_fd_sc_hd__or2_1 _40521_ (.A(_13151_),
    .B(_13153_),
    .X(_13154_));
 sky130_fd_sc_hd__a21oi_2 _40522_ (.A1(_06432_),
    .A2(_09139_),
    .B1(_11972_),
    .Y(_13155_));
 sky130_fd_sc_hd__nor2_2 _40523_ (.A(_13154_),
    .B(_13155_),
    .Y(_13156_));
 sky130_fd_sc_hd__o21a_1 _40524_ (.A1(_13151_),
    .A2(_13153_),
    .B1(_13155_),
    .X(_13157_));
 sky130_fd_sc_hd__nor4_1 _40525_ (.A(_01747_),
    .B(_12026_),
    .C(_13156_),
    .D(_13157_),
    .Y(_13158_));
 sky130_fd_sc_hd__inv_2 _40526_ (.A(_13158_),
    .Y(_13159_));
 sky130_fd_sc_hd__o22ai_1 _40527_ (.A1(_01747_),
    .A2(_12026_),
    .B1(_13156_),
    .B2(_13157_),
    .Y(_13160_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40528_ (.A(_06432_),
    .X(_13161_));
 sky130_fd_sc_hd__nand3_1 _40529_ (.A(_13159_),
    .B(_13160_),
    .C(_13161_),
    .Y(_13162_));
 sky130_fd_sc_hd__a21o_1 _40530_ (.A1(_13159_),
    .A2(_13160_),
    .B1(_13161_),
    .X(_13164_));
 sky130_fd_sc_hd__or2_1 _40531_ (.A(_11743_),
    .B(net190),
    .X(_13165_));
 sky130_fd_sc_hd__a21oi_1 _40532_ (.A1(_13162_),
    .A2(_13164_),
    .B1(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__and3_1 _40533_ (.A(_13165_),
    .B(_13162_),
    .C(_13164_),
    .X(_13167_));
 sky130_fd_sc_hd__nor2_1 _40534_ (.A(_13166_),
    .B(_13167_),
    .Y(_13168_));
 sky130_fd_sc_hd__xor2_1 _40535_ (.A(_11981_),
    .B(_13168_),
    .X(_13169_));
 sky130_fd_sc_hd__nor2_1 _40536_ (.A(_13150_),
    .B(_13169_),
    .Y(_13170_));
 sky130_fd_sc_hd__nand2_1 _40537_ (.A(_13169_),
    .B(_13150_),
    .Y(_13171_));
 sky130_fd_sc_hd__and2b_1 _40538_ (.A_N(_13170_),
    .B(_13171_),
    .X(_13172_));
 sky130_fd_sc_hd__a211o_1 _40539_ (.A1(_10694_),
    .A2(_10695_),
    .B1(_11981_),
    .C1(_11982_),
    .X(_13173_));
 sky130_fd_sc_hd__o21ai_1 _40540_ (.A1(_10810_),
    .A2(_11984_),
    .B1(_13173_),
    .Y(_13175_));
 sky130_fd_sc_hd__nand2_1 _40541_ (.A(_13172_),
    .B(_13175_),
    .Y(_13176_));
 sky130_fd_sc_hd__or2_1 _40542_ (.A(_13175_),
    .B(_13172_),
    .X(_13177_));
 sky130_fd_sc_hd__nand2_1 _40543_ (.A(_13176_),
    .B(_13177_),
    .Y(_13178_));
 sky130_fd_sc_hd__o211ai_2 _40544_ (.A1(_11992_),
    .A2(_11993_),
    .B1(_11990_),
    .C1(_13178_),
    .Y(_13179_));
 sky130_fd_sc_hd__a21o_1 _40545_ (.A1(_11990_),
    .A2(_11995_),
    .B1(_13178_),
    .X(_13180_));
 sky130_fd_sc_hd__nand2_1 _40546_ (.A(_13179_),
    .B(_13180_),
    .Y(_13181_));
 sky130_fd_sc_hd__xor2_1 _40547_ (.A(_13149_),
    .B(_13181_),
    .X(_13182_));
 sky130_fd_sc_hd__a21o_1 _40548_ (.A1(_11736_),
    .A2(_11785_),
    .B1(_11961_),
    .X(_13183_));
 sky130_fd_sc_hd__nor2_1 _40549_ (.A(_13182_),
    .B(_13183_),
    .Y(_13184_));
 sky130_fd_sc_hd__nand2_1 _40550_ (.A(_13183_),
    .B(_13182_),
    .Y(_13186_));
 sky130_fd_sc_hd__or2b_1 _40551_ (.A(_13184_),
    .B_N(_13186_),
    .X(_13187_));
 sky130_fd_sc_hd__xor2_1 _40552_ (.A(_13101_),
    .B(_13187_),
    .X(_13188_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40553_ (.A(_13188_),
    .X(_13189_));
 sky130_fd_sc_hd__nand2_1 _40554_ (.A(_13100_),
    .B(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__nand3_1 _40555_ (.A(_13095_),
    .B(_13032_),
    .C(_13036_),
    .Y(_13191_));
 sky130_fd_sc_hd__a21o_1 _40556_ (.A1(_13032_),
    .A2(_13036_),
    .B1(_13095_),
    .X(_13192_));
 sky130_fd_sc_hd__nand3b_2 _40557_ (.A_N(_12893_),
    .B(_13191_),
    .C(_13192_),
    .Y(_13193_));
 sky130_fd_sc_hd__inv_2 _40558_ (.A(_13193_),
    .Y(_13194_));
 sky130_fd_sc_hd__a2bb2o_1 _40559_ (.A1_N(_12070_),
    .A2_N(_12068_),
    .B1(_12061_),
    .B2(_11958_),
    .X(_13195_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40560_ (.A(_13193_),
    .X(_13197_));
 sky130_fd_sc_hd__a21o_1 _40561_ (.A1(_13197_),
    .A2(_13100_),
    .B1(_13189_),
    .X(_13198_));
 sky130_fd_sc_hd__o211a_1 _40562_ (.A1(_13190_),
    .A2(_13194_),
    .B1(_13195_),
    .C1(_13198_),
    .X(_13199_));
 sky130_fd_sc_hd__a21bo_1 _40563_ (.A1(_13197_),
    .A2(_13100_),
    .B1_N(_13188_),
    .X(_13200_));
 sky130_fd_sc_hd__o2bb2a_1 _40564_ (.A1_N(_12061_),
    .A2_N(_11958_),
    .B1(_12070_),
    .B2(_12068_),
    .X(_13201_));
 sky130_fd_sc_hd__nand3b_1 _40565_ (.A_N(_13189_),
    .B(_13197_),
    .C(_13100_),
    .Y(_13202_));
 sky130_fd_sc_hd__o21ai_2 _40566_ (.A1(_11966_),
    .A2(_12059_),
    .B1(_12058_),
    .Y(_13203_));
 sky130_fd_sc_hd__o21a_1 _40567_ (.A1(_10853_),
    .A2(_11707_),
    .B1(_11708_),
    .X(_13204_));
 sky130_fd_sc_hd__clkbuf_2 _40568_ (.A(_13104_),
    .X(_13205_));
 sky130_fd_sc_hd__nor2_1 _40569_ (.A(_13205_),
    .B(net445),
    .Y(_13206_));
 sky130_fd_sc_hd__and3_1 _40570_ (.A(_12008_),
    .B(_12021_),
    .C(_13206_),
    .X(_13208_));
 sky130_fd_sc_hd__clkbuf_2 _40571_ (.A(_13206_),
    .X(_13209_));
 sky130_fd_sc_hd__a21oi_2 _40572_ (.A1(_12008_),
    .A2(_12021_),
    .B1(_13209_),
    .Y(_13210_));
 sky130_fd_sc_hd__o221a_1 _40573_ (.A1(_13208_),
    .A2(_13210_),
    .B1(_12022_),
    .B2(_12051_),
    .C1(_12050_),
    .X(_13211_));
 sky130_fd_sc_hd__or3b_1 _40574_ (.A(_12019_),
    .B(_12051_),
    .C_N(_12021_),
    .X(_13212_));
 sky130_fd_sc_hd__a211oi_4 _40575_ (.A1(_12050_),
    .A2(_13212_),
    .B1(_13208_),
    .C1(_13210_),
    .Y(_13213_));
 sky130_fd_sc_hd__nor3_2 _40576_ (.A(_13204_),
    .B(_13211_),
    .C(_13213_),
    .Y(_13214_));
 sky130_fd_sc_hd__o221ai_1 _40577_ (.A1(_10853_),
    .A2(_11709_),
    .B1(_13211_),
    .B2(_13213_),
    .C1(_11708_),
    .Y(_13215_));
 sky130_fd_sc_hd__or2b_1 _40578_ (.A(_13214_),
    .B_N(_13215_),
    .X(_13216_));
 sky130_fd_sc_hd__o211a_1 _40579_ (.A1(_11710_),
    .A2(_11711_),
    .B1(_11718_),
    .C1(_13216_),
    .X(_13217_));
 sky130_fd_sc_hd__o21a_1 _40580_ (.A1(_11710_),
    .A2(_11711_),
    .B1(_11718_),
    .X(_13219_));
 sky130_fd_sc_hd__or3b_2 _40581_ (.A(_13219_),
    .B(_13214_),
    .C_N(_13215_),
    .X(_13220_));
 sky130_fd_sc_hd__and2b_1 _40582_ (.A_N(_13217_),
    .B(_13220_),
    .X(_13221_));
 sky130_fd_sc_hd__xnor2_2 _40583_ (.A(_13203_),
    .B(_13221_),
    .Y(_13222_));
 sky130_fd_sc_hd__xnor2_1 _40584_ (.A(_11725_),
    .B(_13222_),
    .Y(_13223_));
 sky130_fd_sc_hd__a31o_1 _40585_ (.A1(_13200_),
    .A2(_13201_),
    .A3(_13202_),
    .B1(_13223_),
    .X(_13224_));
 sky130_fd_sc_hd__o21ai_2 _40586_ (.A1(_12073_),
    .A2(_12093_),
    .B1(_12085_),
    .Y(_13225_));
 sky130_fd_sc_hd__o211ai_2 _40587_ (.A1(_13190_),
    .A2(_13194_),
    .B1(_13195_),
    .C1(_13198_),
    .Y(_13226_));
 sky130_fd_sc_hd__nand3_2 _40588_ (.A(_13200_),
    .B(_13201_),
    .C(_13202_),
    .Y(_13227_));
 sky130_fd_sc_hd__and4_1 _40589_ (.A(_11721_),
    .B(_11717_),
    .C(_11718_),
    .D(_13222_),
    .X(_13228_));
 sky130_fd_sc_hd__nor2_1 _40590_ (.A(_11725_),
    .B(_13222_),
    .Y(_13230_));
 sky130_fd_sc_hd__o2bb2ai_1 _40591_ (.A1_N(_13226_),
    .A2_N(_13227_),
    .B1(_13228_),
    .B2(_13230_),
    .Y(_13231_));
 sky130_fd_sc_hd__o211ai_4 _40592_ (.A1(_13199_),
    .A2(_13224_),
    .B1(_13225_),
    .C1(_13231_),
    .Y(_13232_));
 sky130_fd_sc_hd__nor2_1 _40593_ (.A(_12092_),
    .B(_12079_),
    .Y(_13233_));
 sky130_fd_sc_hd__o211ai_2 _40594_ (.A1(_13228_),
    .A2(_13230_),
    .B1(_13226_),
    .C1(_13227_),
    .Y(_13234_));
 sky130_fd_sc_hd__inv_2 _40595_ (.A(_13222_),
    .Y(_13235_));
 sky130_fd_sc_hd__nand2_1 _40596_ (.A(_11725_),
    .B(_13235_),
    .Y(_13236_));
 sky130_fd_sc_hd__inv_2 _40597_ (.A(_13236_),
    .Y(_13237_));
 sky130_fd_sc_hd__nor2_1 _40598_ (.A(_11725_),
    .B(_13235_),
    .Y(_13238_));
 sky130_fd_sc_hd__o2bb2ai_1 _40599_ (.A1_N(_13226_),
    .A2_N(_13227_),
    .B1(_13237_),
    .B2(_13238_),
    .Y(_13239_));
 sky130_fd_sc_hd__o211ai_4 _40600_ (.A1(_12073_),
    .A2(_13233_),
    .B1(_13234_),
    .C1(_13239_),
    .Y(_13241_));
 sky130_fd_sc_hd__a21oi_1 _40601_ (.A1(_10865_),
    .A2(_11733_),
    .B1(_11728_),
    .Y(_13242_));
 sky130_fd_sc_hd__a21boi_1 _40602_ (.A1(_13232_),
    .A2(_13241_),
    .B1_N(_13242_),
    .Y(_13243_));
 sky130_fd_sc_hd__o211a_2 _40603_ (.A1(_11728_),
    .A2(_12091_),
    .B1(_13232_),
    .C1(_13241_),
    .X(_13244_));
 sky130_fd_sc_hd__a32o_1 _40604_ (.A1(_12089_),
    .A2(_12090_),
    .A3(_12094_),
    .B1(_12088_),
    .B2(_12096_),
    .X(_13245_));
 sky130_fd_sc_hd__o21bai_2 _40605_ (.A1(_13243_),
    .A2(_13244_),
    .B1_N(_13245_),
    .Y(_13246_));
 sky130_fd_sc_hd__a21bo_1 _40606_ (.A1(_13232_),
    .A2(_13241_),
    .B1_N(_13242_),
    .X(_13247_));
 sky130_fd_sc_hd__o211ai_1 _40607_ (.A1(_11728_),
    .A2(_12091_),
    .B1(_13232_),
    .C1(_13241_),
    .Y(_13248_));
 sky130_fd_sc_hd__nand3_2 _40608_ (.A(_13245_),
    .B(_13247_),
    .C(_13248_),
    .Y(_13249_));
 sky130_fd_sc_hd__nand2_1 _40609_ (.A(_13246_),
    .B(_13249_),
    .Y(_13250_));
 sky130_fd_sc_hd__clkbuf_2 _40610_ (.A(_13250_),
    .X(_13252_));
 sky130_fd_sc_hd__nand2_1 _40611_ (.A(_12892_),
    .B(_13252_),
    .Y(_13253_));
 sky130_fd_sc_hd__nand2_2 _40612_ (.A(_13245_),
    .B(_13247_),
    .Y(_13254_));
 sky130_fd_sc_hd__nand3_1 _40613_ (.A(_12106_),
    .B(_12099_),
    .C(_12105_),
    .Y(_13255_));
 sky130_fd_sc_hd__o21ai_1 _40614_ (.A1(_10905_),
    .A2(_10898_),
    .B1(_13255_),
    .Y(_13256_));
 sky130_fd_sc_hd__a21oi_1 _40615_ (.A1(_10490_),
    .A2(_10902_),
    .B1(_13256_),
    .Y(_13257_));
 sky130_fd_sc_hd__nand2_1 _40616_ (.A(_12099_),
    .B(_12105_),
    .Y(_13258_));
 sky130_fd_sc_hd__and2_1 _40617_ (.A(_10896_),
    .B(_12100_),
    .X(_13259_));
 sky130_fd_sc_hd__a22oi_2 _40618_ (.A1(_12116_),
    .A2(_12117_),
    .B1(_13258_),
    .B2(_13259_),
    .Y(_13260_));
 sky130_fd_sc_hd__nand4b_2 _40619_ (.A_N(_10491_),
    .B(_13260_),
    .C(_13255_),
    .D(_10902_),
    .Y(_13261_));
 sky130_fd_sc_hd__o22a_1 _40620_ (.A1(_08124_),
    .A2(_08125_),
    .B1(_06582_),
    .B2(_05094_),
    .X(_13263_));
 sky130_fd_sc_hd__o22ai_4 _40621_ (.A1(_12107_),
    .A2(_13257_),
    .B1(_13261_),
    .B2(_13263_),
    .Y(_13264_));
 sky130_fd_sc_hd__o211ai_4 _40622_ (.A1(_13254_),
    .A2(_13244_),
    .B1(_13246_),
    .C1(_13264_),
    .Y(_13265_));
 sky130_fd_sc_hd__o211a_1 _40623_ (.A1(_12723_),
    .A2(_12726_),
    .B1(_13253_),
    .C1(_13265_),
    .X(_13266_));
 sky130_fd_sc_hd__a21o_1 _40624_ (.A1(_12721_),
    .A2(_12727_),
    .B1(_12723_),
    .X(_13267_));
 sky130_fd_sc_hd__a21oi_1 _40625_ (.A1(_13253_),
    .A2(_13265_),
    .B1(_13267_),
    .Y(_13268_));
 sky130_fd_sc_hd__o21ai_1 _40626_ (.A1(_13266_),
    .A2(_13268_),
    .B1(_12127_),
    .Y(_13269_));
 sky130_fd_sc_hd__buf_2 _40627_ (.A(_12723_),
    .X(_13270_));
 sky130_fd_sc_hd__o211ai_1 _40628_ (.A1(_13270_),
    .A2(_12726_),
    .B1(_13253_),
    .C1(_13265_),
    .Y(_13271_));
 sky130_fd_sc_hd__a21o_1 _40629_ (.A1(_13253_),
    .A2(_13265_),
    .B1(_13267_),
    .X(_13272_));
 sky130_fd_sc_hd__nand3_1 _40630_ (.A(_10934_),
    .B(_13271_),
    .C(_13272_),
    .Y(_13274_));
 sky130_fd_sc_hd__and2b_1 _40631_ (.A_N(_12729_),
    .B(_12719_),
    .X(_13275_));
 sky130_fd_sc_hd__nor2_1 _40632_ (.A(_12718_),
    .B(_13275_),
    .Y(_13276_));
 sky130_fd_sc_hd__nand3_2 _40633_ (.A(_13269_),
    .B(_13274_),
    .C(_13276_),
    .Y(_13277_));
 sky130_fd_sc_hd__nand3_1 _40634_ (.A(_13272_),
    .B(_10939_),
    .C(_13271_),
    .Y(_13278_));
 sky130_fd_sc_hd__o21ai_1 _40635_ (.A1(_13266_),
    .A2(_13268_),
    .B1(_10934_),
    .Y(_13279_));
 sky130_fd_sc_hd__o211ai_2 _40636_ (.A1(_12718_),
    .A2(_13275_),
    .B1(_13278_),
    .C1(_13279_),
    .Y(_13280_));
 sky130_fd_sc_hd__buf_4 _40637_ (.A(_13280_),
    .X(_13281_));
 sky130_fd_sc_hd__o211ai_4 _40638_ (.A1(_12122_),
    .A2(_12886_),
    .B1(_13277_),
    .C1(_13281_),
    .Y(_13282_));
 sky130_fd_sc_hd__o21ai_1 _40639_ (.A1(_10935_),
    .A2(_12124_),
    .B1(_12128_),
    .Y(_13283_));
 sky130_fd_sc_hd__a21o_1 _40640_ (.A1(_13277_),
    .A2(_13281_),
    .B1(_13283_),
    .X(_13285_));
 sky130_fd_sc_hd__nand3_1 _40641_ (.A(_12884_),
    .B(_13282_),
    .C(_13285_),
    .Y(_13286_));
 sky130_fd_sc_hd__clkbuf_2 _40642_ (.A(_13286_),
    .X(_13287_));
 sky130_fd_sc_hd__o211a_1 _40643_ (.A1(_12122_),
    .A2(_12886_),
    .B1(_13277_),
    .C1(_13281_),
    .X(_13288_));
 sky130_fd_sc_hd__a21oi_1 _40644_ (.A1(_13277_),
    .A2(_13281_),
    .B1(_13283_),
    .Y(_13289_));
 sky130_fd_sc_hd__o221ai_4 _40645_ (.A1(_12137_),
    .A2(_12135_),
    .B1(_13288_),
    .B2(_13289_),
    .C1(_12133_),
    .Y(_13290_));
 sky130_fd_sc_hd__o211ai_1 _40646_ (.A1(_12879_),
    .A2(_12883_),
    .B1(_13287_),
    .C1(_13290_),
    .Y(_13291_));
 sky130_fd_sc_hd__and3_1 _40647_ (.A(_06607_),
    .B(_12880_),
    .C(_12878_),
    .X(_13292_));
 sky130_fd_sc_hd__buf_2 _40648_ (.A(_06607_),
    .X(_13293_));
 sky130_fd_sc_hd__buf_2 _40649_ (.A(_12880_),
    .X(_13294_));
 sky130_fd_sc_hd__clkbuf_2 _40650_ (.A(_13294_),
    .X(_13296_));
 sky130_fd_sc_hd__a21oi_1 _40651_ (.A1(_13293_),
    .A2(_13296_),
    .B1(_12878_),
    .Y(_13297_));
 sky130_fd_sc_hd__o2bb2ai_1 _40652_ (.A1_N(_13286_),
    .A2_N(_13290_),
    .B1(_13292_),
    .B2(_13297_),
    .Y(_13298_));
 sky130_fd_sc_hd__nand3_1 _40653_ (.A(_12874_),
    .B(_13291_),
    .C(_13298_),
    .Y(_13299_));
 sky130_fd_sc_hd__o2bb2ai_1 _40654_ (.A1_N(_13287_),
    .A2_N(_13290_),
    .B1(_12879_),
    .B2(_12883_),
    .Y(_13300_));
 sky130_fd_sc_hd__inv_2 _40655_ (.A(_12874_),
    .Y(_13301_));
 sky130_fd_sc_hd__o211ai_1 _40656_ (.A1(_13292_),
    .A2(_13297_),
    .B1(_13287_),
    .C1(_13290_),
    .Y(_13302_));
 sky130_fd_sc_hd__nand3_1 _40657_ (.A(_13300_),
    .B(_13301_),
    .C(_13302_),
    .Y(_13303_));
 sky130_fd_sc_hd__a21o_1 _40658_ (.A1(_12144_),
    .A2(_12158_),
    .B1(_12166_),
    .X(_13304_));
 sky130_fd_sc_hd__a21o_1 _40659_ (.A1(_13299_),
    .A2(_13303_),
    .B1(_13304_),
    .X(_13305_));
 sky130_fd_sc_hd__clkbuf_2 _40660_ (.A(_13299_),
    .X(_13307_));
 sky130_fd_sc_hd__nand3_1 _40661_ (.A(_13304_),
    .B(_13307_),
    .C(_13303_),
    .Y(_13308_));
 sky130_fd_sc_hd__a31oi_4 _40662_ (.A1(_12606_),
    .A2(_12565_),
    .A3(_12564_),
    .B1(_12604_),
    .Y(_13309_));
 sky130_fd_sc_hd__clkbuf_2 _40663_ (.A(_10168_),
    .X(_13310_));
 sky130_fd_sc_hd__and4b_1 _40664_ (.A_N(_08784_),
    .B(_13310_),
    .C(_04266_),
    .D(_12558_),
    .X(_13311_));
 sky130_fd_sc_hd__o21a_1 _40665_ (.A1(_12558_),
    .A2(_10168_),
    .B1(_06990_),
    .X(_13312_));
 sky130_fd_sc_hd__a211oi_1 _40666_ (.A1(_12558_),
    .A2(_13310_),
    .B1(_06994_),
    .C1(_13312_),
    .Y(_13313_));
 sky130_fd_sc_hd__o221a_1 _40667_ (.A1(_11329_),
    .A2(_12561_),
    .B1(_13311_),
    .B2(_13313_),
    .C1(_12564_),
    .X(_13314_));
 sky130_fd_sc_hd__a211oi_1 _40668_ (.A1(_12563_),
    .A2(_12564_),
    .B1(_13311_),
    .C1(_13313_),
    .Y(_13315_));
 sky130_fd_sc_hd__or4_1 _40669_ (.A(_11363_),
    .B(_12573_),
    .C(net191),
    .D(_11362_),
    .X(_13316_));
 sky130_fd_sc_hd__buf_1 _40670_ (.A(net329),
    .X(_13318_));
 sky130_fd_sc_hd__and4_1 _40671_ (.A(_05509_),
    .B(_02221_),
    .C(_12568_),
    .D(_13318_),
    .X(_13319_));
 sky130_fd_sc_hd__a21oi_1 _40672_ (.A1(_13318_),
    .A2(_12568_),
    .B1(_05500_),
    .Y(_13320_));
 sky130_fd_sc_hd__and3_1 _40673_ (.A(_05500_),
    .B(_13318_),
    .C(_12568_),
    .X(_13321_));
 sky130_fd_sc_hd__o2111ai_2 _40674_ (.A1(_13320_),
    .A2(_13321_),
    .B1(_02220_),
    .C1(_04319_),
    .D1(_04317_),
    .Y(_13322_));
 sky130_fd_sc_hd__a311o_1 _40675_ (.A1(_02220_),
    .A2(_04319_),
    .A3(_04317_),
    .B1(_13320_),
    .C1(_13321_),
    .X(_13323_));
 sky130_fd_sc_hd__o211ai_1 _40676_ (.A1(_12572_),
    .A2(_13319_),
    .B1(_13322_),
    .C1(_13323_),
    .Y(_13324_));
 sky130_fd_sc_hd__inv_2 _40677_ (.A(_13324_),
    .Y(_13325_));
 sky130_fd_sc_hd__a211oi_1 _40678_ (.A1(_13322_),
    .A2(_13323_),
    .B1(_12572_),
    .C1(_13319_),
    .Y(_13326_));
 sky130_fd_sc_hd__nor4_1 _40679_ (.A(_12574_),
    .B(_12573_),
    .C(_13325_),
    .D(_13326_),
    .Y(_13327_));
 sky130_fd_sc_hd__o22a_1 _40680_ (.A1(_12574_),
    .A2(_12573_),
    .B1(_13325_),
    .B2(_13326_),
    .X(_13329_));
 sky130_fd_sc_hd__a211oi_2 _40681_ (.A1(_12578_),
    .A2(_13316_),
    .B1(net145),
    .C1(_13329_),
    .Y(_13330_));
 sky130_fd_sc_hd__buf_1 _40682_ (.A(_13327_),
    .X(_13331_));
 sky130_fd_sc_hd__o211ai_1 _40683_ (.A1(_13331_),
    .A2(_13329_),
    .B1(_12578_),
    .C1(_13316_),
    .Y(_13332_));
 sky130_fd_sc_hd__nand2b_1 _40684_ (.A_N(_13330_),
    .B(_13332_),
    .Y(_13333_));
 sky130_fd_sc_hd__nor2_1 _40685_ (.A(_12590_),
    .B(_12591_),
    .Y(_13334_));
 sky130_fd_sc_hd__and3_1 _40686_ (.A(_10154_),
    .B(_11345_),
    .C(_13334_),
    .X(_13335_));
 sky130_fd_sc_hd__buf_1 _40687_ (.A(_11349_),
    .X(_13336_));
 sky130_fd_sc_hd__xor2_1 _40688_ (.A(net334),
    .B(\delay_line[26][15] ),
    .X(_13337_));
 sky130_fd_sc_hd__or2_1 _40689_ (.A(_10146_),
    .B(_13337_),
    .X(_13338_));
 sky130_fd_sc_hd__nand2_1 _40690_ (.A(_10146_),
    .B(_13337_),
    .Y(_13340_));
 sky130_fd_sc_hd__a21bo_1 _40691_ (.A1(_05531_),
    .A2(_12584_),
    .B1_N(_12585_),
    .X(_13341_));
 sky130_fd_sc_hd__a21oi_1 _40692_ (.A1(_13338_),
    .A2(_13340_),
    .B1(_13341_),
    .Y(_13342_));
 sky130_fd_sc_hd__and3_1 _40693_ (.A(_13341_),
    .B(_13338_),
    .C(_13340_),
    .X(_13343_));
 sky130_fd_sc_hd__nor2_1 _40694_ (.A(_13342_),
    .B(_13343_),
    .Y(_13344_));
 sky130_fd_sc_hd__a21oi_1 _40695_ (.A1(_12579_),
    .A2(_13334_),
    .B1(_12590_),
    .Y(_13345_));
 sky130_fd_sc_hd__xnor2_1 _40696_ (.A(_13344_),
    .B(_13345_),
    .Y(_13346_));
 sky130_fd_sc_hd__nand2_1 _40697_ (.A(_13336_),
    .B(_13346_),
    .Y(_13347_));
 sky130_fd_sc_hd__or2_1 _40698_ (.A(_13336_),
    .B(_13346_),
    .X(_13348_));
 sky130_fd_sc_hd__o211ai_2 _40699_ (.A1(_12597_),
    .A2(_13335_),
    .B1(_13347_),
    .C1(_13348_),
    .Y(_13349_));
 sky130_fd_sc_hd__a221o_1 _40700_ (.A1(_13334_),
    .A2(net244),
    .B1(_13347_),
    .B2(_13348_),
    .C1(_12597_),
    .X(_13351_));
 sky130_fd_sc_hd__o211ai_1 _40701_ (.A1(_11351_),
    .A2(_11348_),
    .B1(_12599_),
    .C1(_12600_),
    .Y(_13352_));
 sky130_fd_sc_hd__o31ai_2 _40702_ (.A1(_12582_),
    .A2(_12596_),
    .A3(_12597_),
    .B1(_13352_),
    .Y(_13353_));
 sky130_fd_sc_hd__and3_1 _40703_ (.A(_13349_),
    .B(_13351_),
    .C(_13353_),
    .X(_13354_));
 sky130_fd_sc_hd__a21oi_1 _40704_ (.A1(_13349_),
    .A2(_13351_),
    .B1(_13353_),
    .Y(_13355_));
 sky130_fd_sc_hd__or2_1 _40705_ (.A(_13354_),
    .B(_13355_),
    .X(_13356_));
 sky130_fd_sc_hd__xnor2_1 _40706_ (.A(_13333_),
    .B(_13356_),
    .Y(_13357_));
 sky130_fd_sc_hd__o21ai_1 _40707_ (.A1(_13314_),
    .A2(_13315_),
    .B1(_13357_),
    .Y(_13358_));
 sky130_fd_sc_hd__or3_2 _40708_ (.A(_13314_),
    .B(_13315_),
    .C(_13357_),
    .X(_13359_));
 sky130_fd_sc_hd__nand2_1 _40709_ (.A(_13358_),
    .B(_13359_),
    .Y(_13360_));
 sky130_fd_sc_hd__xnor2_1 _40710_ (.A(_13309_),
    .B(_13360_),
    .Y(_13362_));
 sky130_fd_sc_hd__o21ai_1 _40711_ (.A1(_11400_),
    .A2(_11403_),
    .B1(_12551_),
    .Y(_13363_));
 sky130_fd_sc_hd__nand2_1 _40712_ (.A(_11398_),
    .B(_12546_),
    .Y(_13364_));
 sky130_fd_sc_hd__or2b_1 _40713_ (.A(_12544_),
    .B_N(_11382_),
    .X(_13365_));
 sky130_fd_sc_hd__buf_1 _40714_ (.A(_08857_),
    .X(_13366_));
 sky130_fd_sc_hd__or4b_1 _40715_ (.A(_10237_),
    .B(_08859_),
    .C(_06962_),
    .D_N(_13366_),
    .X(_13367_));
 sky130_fd_sc_hd__a22o_1 _40716_ (.A1(_04353_),
    .A2(_13366_),
    .B1(_05410_),
    .B2(_05413_),
    .X(_13368_));
 sky130_fd_sc_hd__and2_1 _40717_ (.A(_13367_),
    .B(_13368_),
    .X(_13369_));
 sky130_fd_sc_hd__nand2_1 _40718_ (.A(_13365_),
    .B(_13369_),
    .Y(_13370_));
 sky130_fd_sc_hd__a21o_1 _40719_ (.A1(_13367_),
    .A2(_13368_),
    .B1(_13365_),
    .X(_13371_));
 sky130_fd_sc_hd__nand3b_1 _40720_ (.A_N(_08864_),
    .B(_10244_),
    .C(_12543_),
    .Y(_13373_));
 sky130_fd_sc_hd__a21oi_1 _40721_ (.A1(_13370_),
    .A2(_13371_),
    .B1(_13373_),
    .Y(_13374_));
 sky130_fd_sc_hd__and3_1 _40722_ (.A(_13373_),
    .B(_13370_),
    .C(_13371_),
    .X(_13375_));
 sky130_fd_sc_hd__a2bb2o_1 _40723_ (.A1_N(_11390_),
    .A2_N(_13365_),
    .B1(_11387_),
    .B2(_12545_),
    .X(_13376_));
 sky130_fd_sc_hd__or3b_2 _40724_ (.A(_13374_),
    .B(_13375_),
    .C_N(_13376_),
    .X(_13377_));
 sky130_fd_sc_hd__o21bai_1 _40725_ (.A1(_13374_),
    .A2(_13375_),
    .B1_N(_13376_),
    .Y(_13378_));
 sky130_fd_sc_hd__and2_1 _40726_ (.A(_13377_),
    .B(_13378_),
    .X(_13379_));
 sky130_fd_sc_hd__and3_1 _40727_ (.A(_11393_),
    .B(_12546_),
    .C(_13379_),
    .X(_13380_));
 sky130_fd_sc_hd__a21oi_1 _40728_ (.A1(_11393_),
    .A2(_12546_),
    .B1(_13379_),
    .Y(_13381_));
 sky130_fd_sc_hd__or2_1 _40729_ (.A(_13380_),
    .B(_13381_),
    .X(_13382_));
 sky130_fd_sc_hd__a21oi_2 _40730_ (.A1(_13363_),
    .A2(_13364_),
    .B1(_13382_),
    .Y(_13384_));
 sky130_fd_sc_hd__and3_1 _40731_ (.A(_13363_),
    .B(_13364_),
    .C(_13382_),
    .X(_13385_));
 sky130_fd_sc_hd__nor2_4 _40732_ (.A(_13384_),
    .B(_13385_),
    .Y(_13386_));
 sky130_fd_sc_hd__o21ai_1 _40733_ (.A1(_10188_),
    .A2(_10190_),
    .B1(_11450_),
    .Y(_13387_));
 sky130_fd_sc_hd__nor2_1 _40734_ (.A(_11447_),
    .B(_11448_),
    .Y(_13388_));
 sky130_fd_sc_hd__a21o_1 _40735_ (.A1(_13387_),
    .A2(_13388_),
    .B1(_12508_),
    .X(_13389_));
 sky130_fd_sc_hd__a32o_1 _40736_ (.A1(_11442_),
    .A2(_06941_),
    .A3(_10183_),
    .B1(_12507_),
    .B2(_13389_),
    .X(_13390_));
 sky130_fd_sc_hd__xnor2_2 _40737_ (.A(\delay_line[29][14] ),
    .B(_12506_),
    .Y(_13391_));
 sky130_fd_sc_hd__xnor2_2 _40738_ (.A(_13390_),
    .B(_13391_),
    .Y(_13392_));
 sky130_fd_sc_hd__o211a_1 _40739_ (.A1(_10220_),
    .A2(_10223_),
    .B1(_11432_),
    .C1(_12533_),
    .X(_13393_));
 sky130_fd_sc_hd__inv_2 _40740_ (.A(_13393_),
    .Y(_13395_));
 sky130_fd_sc_hd__or3_1 _40741_ (.A(_02110_),
    .B(_12513_),
    .C(_10210_),
    .X(_13396_));
 sky130_fd_sc_hd__a211o_1 _40742_ (.A1(_08895_),
    .A2(_11410_),
    .B1(_10205_),
    .C1(_10208_),
    .X(_13397_));
 sky130_fd_sc_hd__a211oi_1 _40743_ (.A1(_13396_),
    .A2(_13397_),
    .B1(_12514_),
    .C1(net176),
    .Y(_13398_));
 sky130_fd_sc_hd__o211a_1 _40744_ (.A1(_12514_),
    .A2(net176),
    .B1(_13396_),
    .C1(_13397_),
    .X(_13399_));
 sky130_fd_sc_hd__or2_1 _40745_ (.A(_13398_),
    .B(_13399_),
    .X(_13400_));
 sky130_fd_sc_hd__o21ba_1 _40746_ (.A1(_12519_),
    .A2(net187),
    .B1_N(_13400_),
    .X(_13401_));
 sky130_fd_sc_hd__nor3b_1 _40747_ (.A(_12519_),
    .B(net187),
    .C_N(_13400_),
    .Y(_13402_));
 sky130_fd_sc_hd__nor2_1 _40748_ (.A(_13401_),
    .B(_13402_),
    .Y(_13403_));
 sky130_fd_sc_hd__nor2_1 _40749_ (.A(net164),
    .B(_12528_),
    .Y(_13404_));
 sky130_fd_sc_hd__xnor2_1 _40750_ (.A(_13403_),
    .B(_13404_),
    .Y(_13406_));
 sky130_fd_sc_hd__or4b_2 _40751_ (.A(_12528_),
    .B(_12529_),
    .C(_12530_),
    .D_N(_13406_),
    .X(_13407_));
 sky130_fd_sc_hd__or2_1 _40752_ (.A(_12531_),
    .B(_13406_),
    .X(_13408_));
 sky130_fd_sc_hd__nand2_1 _40753_ (.A(_13407_),
    .B(_13408_),
    .Y(_13409_));
 sky130_fd_sc_hd__a21oi_1 _40754_ (.A1(_13395_),
    .A2(_12539_),
    .B1(_13409_),
    .Y(_13410_));
 sky130_fd_sc_hd__and3_1 _40755_ (.A(_13395_),
    .B(_12539_),
    .C(_13409_),
    .X(_13411_));
 sky130_fd_sc_hd__or2_1 _40756_ (.A(_13410_),
    .B(_13411_),
    .X(_13412_));
 sky130_fd_sc_hd__xnor2_2 _40757_ (.A(_13392_),
    .B(_13412_),
    .Y(_13413_));
 sky130_fd_sc_hd__xor2_4 _40758_ (.A(_13386_),
    .B(_13413_),
    .X(_13414_));
 sky130_fd_sc_hd__nand2_1 _40759_ (.A(_13362_),
    .B(_13414_),
    .Y(_13415_));
 sky130_fd_sc_hd__or2_1 _40760_ (.A(_13362_),
    .B(_13414_),
    .X(_13417_));
 sky130_fd_sc_hd__nand2_2 _40761_ (.A(_13415_),
    .B(_13417_),
    .Y(_13418_));
 sky130_fd_sc_hd__o211ai_2 _40762_ (.A1(_12388_),
    .A2(_12489_),
    .B1(_12490_),
    .C1(_13418_),
    .Y(_13419_));
 sky130_fd_sc_hd__or2_1 _40763_ (.A(_12388_),
    .B(_12489_),
    .X(_13420_));
 sky130_fd_sc_hd__a21o_1 _40764_ (.A1(_12490_),
    .A2(_13420_),
    .B1(_13418_),
    .X(_13421_));
 sky130_fd_sc_hd__a21bo_1 _40765_ (.A1(_12556_),
    .A2(_12607_),
    .B1_N(_12610_),
    .X(_13422_));
 sky130_fd_sc_hd__a21oi_2 _40766_ (.A1(_13419_),
    .A2(_13421_),
    .B1(_13422_),
    .Y(_13423_));
 sky130_fd_sc_hd__and3_1 _40767_ (.A(_13422_),
    .B(_13419_),
    .C(_13421_),
    .X(_13424_));
 sky130_fd_sc_hd__o21ai_1 _40768_ (.A1(_12444_),
    .A2(_12448_),
    .B1(_12445_),
    .Y(_13425_));
 sky130_fd_sc_hd__buf_1 _40769_ (.A(_07164_),
    .X(_13426_));
 sky130_fd_sc_hd__buf_1 _40770_ (.A(_07159_),
    .X(_13428_));
 sky130_fd_sc_hd__or4b_1 _40771_ (.A(_13426_),
    .B(_13428_),
    .C(_12432_),
    .D_N(_12420_),
    .X(_13429_));
 sky130_fd_sc_hd__or2_1 _40772_ (.A(_13426_),
    .B(_13428_),
    .X(_13430_));
 sky130_fd_sc_hd__o21ai_1 _40773_ (.A1(_12432_),
    .A2(_11277_),
    .B1(_13430_),
    .Y(_13431_));
 sky130_fd_sc_hd__a21oi_1 _40774_ (.A1(_13430_),
    .A2(_12420_),
    .B1(_11269_),
    .Y(_13432_));
 sky130_fd_sc_hd__and3_1 _40775_ (.A(_13430_),
    .B(_12420_),
    .C(_11269_),
    .X(_13433_));
 sky130_fd_sc_hd__a211o_1 _40776_ (.A1(_13429_),
    .A2(_13431_),
    .B1(_13432_),
    .C1(_13433_),
    .X(_13434_));
 sky130_fd_sc_hd__o211ai_1 _40777_ (.A1(_13433_),
    .A2(_13432_),
    .B1(_13431_),
    .C1(_13429_),
    .Y(_13435_));
 sky130_fd_sc_hd__nor2_1 _40778_ (.A(_12431_),
    .B(_12433_),
    .Y(_13436_));
 sky130_fd_sc_hd__a221o_1 _40779_ (.A1(_13434_),
    .A2(_13435_),
    .B1(_12424_),
    .B2(_12434_),
    .C1(_13436_),
    .X(_13437_));
 sky130_fd_sc_hd__and2_1 _40780_ (.A(_12424_),
    .B(_12434_),
    .X(_13439_));
 sky130_fd_sc_hd__o211ai_1 _40781_ (.A1(_13436_),
    .A2(_13439_),
    .B1(_13434_),
    .C1(_13435_),
    .Y(_13440_));
 sky130_fd_sc_hd__nand2_1 _40782_ (.A(_13437_),
    .B(_13440_),
    .Y(_13441_));
 sky130_fd_sc_hd__xnor2_1 _40783_ (.A(_12423_),
    .B(_13441_),
    .Y(_13442_));
 sky130_fd_sc_hd__o21a_1 _40784_ (.A1(_12437_),
    .A2(_12441_),
    .B1(_13442_),
    .X(_13443_));
 sky130_fd_sc_hd__inv_2 _40785_ (.A(_13443_),
    .Y(_13444_));
 sky130_fd_sc_hd__a211o_1 _40786_ (.A1(_11270_),
    .A2(_12440_),
    .B1(_13442_),
    .C1(_12437_),
    .X(_13445_));
 sky130_fd_sc_hd__nand2_1 _40787_ (.A(_13444_),
    .B(_13445_),
    .Y(_13446_));
 sky130_fd_sc_hd__inv_2 _40788_ (.A(_13446_),
    .Y(_13447_));
 sky130_fd_sc_hd__nand2_1 _40789_ (.A(_13425_),
    .B(_13447_),
    .Y(_13448_));
 sky130_fd_sc_hd__or2_1 _40790_ (.A(_13447_),
    .B(_13425_),
    .X(_13450_));
 sky130_fd_sc_hd__inv_2 _40791_ (.A(_12480_),
    .Y(_13451_));
 sky130_fd_sc_hd__a21o_1 _40792_ (.A1(_12452_),
    .A2(_13451_),
    .B1(_12478_),
    .X(_13452_));
 sky130_fd_sc_hd__and3_1 _40793_ (.A(_12469_),
    .B(_12453_),
    .C(_10057_),
    .X(_13453_));
 sky130_fd_sc_hd__and2b_1 _40794_ (.A_N(_10036_),
    .B(_10039_),
    .X(_13454_));
 sky130_fd_sc_hd__buf_1 _40795_ (.A(_10039_),
    .X(_13455_));
 sky130_fd_sc_hd__and2b_1 _40796_ (.A_N(_13455_),
    .B(_10036_),
    .X(_13456_));
 sky130_fd_sc_hd__or2_1 _40797_ (.A(_13455_),
    .B(_12454_),
    .X(_13457_));
 sky130_fd_sc_hd__o31a_1 _40798_ (.A1(_11237_),
    .A2(_13454_),
    .A3(_13456_),
    .B1(_13457_),
    .X(_13458_));
 sky130_fd_sc_hd__a21oi_1 _40799_ (.A1(_08456_),
    .A2(_10038_),
    .B1(_13458_),
    .Y(_13459_));
 sky130_fd_sc_hd__o311a_1 _40800_ (.A1(_11237_),
    .A2(_13454_),
    .A3(_13456_),
    .B1(_12459_),
    .C1(_13457_),
    .X(_13461_));
 sky130_fd_sc_hd__a211o_1 _40801_ (.A1(_12457_),
    .A2(_12462_),
    .B1(_13459_),
    .C1(_13461_),
    .X(_13462_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40802_ (.A(_11237_),
    .X(_13463_));
 sky130_fd_sc_hd__o211ai_2 _40803_ (.A1(_13459_),
    .A2(_13461_),
    .B1(_12457_),
    .C1(_12462_),
    .Y(_13464_));
 sky130_fd_sc_hd__buf_1 _40804_ (.A(_10036_),
    .X(_13465_));
 sky130_fd_sc_hd__or3_1 _40805_ (.A(_13465_),
    .B(_12469_),
    .C(_11233_),
    .X(_13466_));
 sky130_fd_sc_hd__and4_1 _40806_ (.A(_13462_),
    .B(_13463_),
    .C(_13464_),
    .D(_13466_),
    .X(_13467_));
 sky130_fd_sc_hd__and3b_1 _40807_ (.A_N(_13465_),
    .B(_13463_),
    .C(_12453_),
    .X(_13468_));
 sky130_fd_sc_hd__o2bb2a_1 _40808_ (.A1_N(_13464_),
    .A2_N(_13462_),
    .B1(_13468_),
    .B2(_12469_),
    .X(_13469_));
 sky130_fd_sc_hd__a21o_1 _40809_ (.A1(_11245_),
    .A2(_11244_),
    .B1(_12464_),
    .X(_13470_));
 sky130_fd_sc_hd__o221a_1 _40810_ (.A1(_12466_),
    .A2(_12467_),
    .B1(_13467_),
    .B2(_13469_),
    .C1(_13470_),
    .X(_13472_));
 sky130_fd_sc_hd__a211o_1 _40811_ (.A1(_13470_),
    .A2(_12468_),
    .B1(_13467_),
    .C1(_13469_),
    .X(_13473_));
 sky130_fd_sc_hd__and2b_1 _40812_ (.A_N(_13472_),
    .B(_13473_),
    .X(_13474_));
 sky130_fd_sc_hd__xnor2_1 _40813_ (.A(_13453_),
    .B(_13474_),
    .Y(_13475_));
 sky130_fd_sc_hd__o21a_1 _40814_ (.A1(_11234_),
    .A2(_12474_),
    .B1(_12475_),
    .X(_13476_));
 sky130_fd_sc_hd__or2_1 _40815_ (.A(_13475_),
    .B(_13476_),
    .X(_13477_));
 sky130_fd_sc_hd__nand2_1 _40816_ (.A(_13475_),
    .B(_13476_),
    .Y(_13478_));
 sky130_fd_sc_hd__nand2_1 _40817_ (.A(_13477_),
    .B(_13478_),
    .Y(_13479_));
 sky130_fd_sc_hd__xnor2_2 _40818_ (.A(_13452_),
    .B(_13479_),
    .Y(_13480_));
 sky130_fd_sc_hd__a21oi_1 _40819_ (.A1(_13448_),
    .A2(_13450_),
    .B1(_13480_),
    .Y(_13481_));
 sky130_fd_sc_hd__and3_1 _40820_ (.A(_13448_),
    .B(_13450_),
    .C(_13480_),
    .X(_13483_));
 sky130_fd_sc_hd__a21oi_1 _40821_ (.A1(_12415_),
    .A2(_12413_),
    .B1(_12411_),
    .Y(_13484_));
 sky130_fd_sc_hd__and4b_1 _40822_ (.A_N(_11219_),
    .B(_12403_),
    .C(_08408_),
    .D(_10005_),
    .X(_13485_));
 sky130_fd_sc_hd__nor2_1 _40823_ (.A(_12406_),
    .B(_13485_),
    .Y(_13486_));
 sky130_fd_sc_hd__or3b_1 _40824_ (.A(_11202_),
    .B(_12391_),
    .C_N(_11219_),
    .X(_13487_));
 sky130_fd_sc_hd__buf_1 _40825_ (.A(_10008_),
    .X(_13488_));
 sky130_fd_sc_hd__and3_1 _40826_ (.A(_07084_),
    .B(_13488_),
    .C(_11209_),
    .X(_13489_));
 sky130_fd_sc_hd__buf_1 _40827_ (.A(_11205_),
    .X(_13490_));
 sky130_fd_sc_hd__nor2_1 _40828_ (.A(_11205_),
    .B(_11209_),
    .Y(_13491_));
 sky130_fd_sc_hd__a221o_1 _40829_ (.A1(_11206_),
    .A2(_10008_),
    .B1(_04144_),
    .B2(_13490_),
    .C1(_13491_),
    .X(_13492_));
 sky130_fd_sc_hd__a21o_1 _40830_ (.A1(_13490_),
    .A2(_04144_),
    .B1(_13491_),
    .X(_13494_));
 sky130_fd_sc_hd__nand3_1 _40831_ (.A(_13494_),
    .B(_13488_),
    .C(_11206_),
    .Y(_13495_));
 sky130_fd_sc_hd__or4bb_1 _40832_ (.A(_13489_),
    .B(_12397_),
    .C_N(_13492_),
    .D_N(_13495_),
    .X(_13496_));
 sky130_fd_sc_hd__a2bb2o_1 _40833_ (.A1_N(_13489_),
    .A2_N(_12397_),
    .B1(_13492_),
    .B2(_13495_),
    .X(_13497_));
 sky130_fd_sc_hd__nand4_2 _40834_ (.A(_13496_),
    .B(_12391_),
    .C(_12393_),
    .D(_13497_),
    .Y(_13498_));
 sky130_fd_sc_hd__a22o_1 _40835_ (.A1(_12391_),
    .A2(_12393_),
    .B1(_13496_),
    .B2(_13497_),
    .X(_13499_));
 sky130_fd_sc_hd__a21oi_1 _40836_ (.A1(_12392_),
    .A2(_12400_),
    .B1(_12399_),
    .Y(_13500_));
 sky130_fd_sc_hd__a21oi_1 _40837_ (.A1(_13498_),
    .A2(_13499_),
    .B1(_13500_),
    .Y(_13501_));
 sky130_fd_sc_hd__nor2_1 _40838_ (.A(_13487_),
    .B(_13501_),
    .Y(_13502_));
 sky130_fd_sc_hd__a31o_1 _40839_ (.A1(_13500_),
    .A2(_13498_),
    .A3(_13499_),
    .B1(_13502_),
    .X(_13503_));
 sky130_fd_sc_hd__a21o_1 _40840_ (.A1(_13487_),
    .A2(_13501_),
    .B1(_13503_),
    .X(_13505_));
 sky130_fd_sc_hd__and2_1 _40841_ (.A(_13486_),
    .B(_13505_),
    .X(_13506_));
 sky130_fd_sc_hd__nor2_1 _40842_ (.A(_13505_),
    .B(_13486_),
    .Y(_13507_));
 sky130_fd_sc_hd__or2_1 _40843_ (.A(_13506_),
    .B(_13507_),
    .X(_13508_));
 sky130_fd_sc_hd__xnor2_1 _40844_ (.A(_13484_),
    .B(_13508_),
    .Y(_13509_));
 sky130_fd_sc_hd__o21a_1 _40845_ (.A1(_13481_),
    .A2(_13483_),
    .B1(_13509_),
    .X(_13510_));
 sky130_fd_sc_hd__nor3_2 _40846_ (.A(_13509_),
    .B(_13481_),
    .C(_13483_),
    .Y(_13511_));
 sky130_fd_sc_hd__o211a_1 _40847_ (.A1(_13510_),
    .A2(_13511_),
    .B1(_12297_),
    .C1(net87),
    .X(_13512_));
 sky130_fd_sc_hd__a211oi_4 _40848_ (.A1(_12297_),
    .A2(net87),
    .B1(_13510_),
    .C1(_13511_),
    .Y(_13513_));
 sky130_fd_sc_hd__a211oi_4 _40849_ (.A1(_12484_),
    .A2(_12487_),
    .B1(_13512_),
    .C1(_13513_),
    .Y(_13514_));
 sky130_fd_sc_hd__o221a_1 _40850_ (.A1(_12417_),
    .A2(_12485_),
    .B1(_13512_),
    .B2(_13513_),
    .C1(_12484_),
    .X(_13516_));
 sky130_fd_sc_hd__nand3_1 _40851_ (.A(_11151_),
    .B(_11156_),
    .C(_12343_),
    .Y(_13517_));
 sky130_fd_sc_hd__and3_1 _40852_ (.A(_02434_),
    .B(_11131_),
    .C(_08611_),
    .X(_13518_));
 sky130_fd_sc_hd__buf_1 _40853_ (.A(_09925_),
    .X(_13519_));
 sky130_fd_sc_hd__nor2_1 _40854_ (.A(_03955_),
    .B(_03956_),
    .Y(_13520_));
 sky130_fd_sc_hd__buf_1 _40855_ (.A(_09926_),
    .X(_13521_));
 sky130_fd_sc_hd__nor2_1 _40856_ (.A(_09926_),
    .B(_08598_),
    .Y(_13522_));
 sky130_fd_sc_hd__a221o_1 _40857_ (.A1(_09924_),
    .A2(_13519_),
    .B1(_13520_),
    .B2(_13521_),
    .C1(_13522_),
    .X(_13523_));
 sky130_fd_sc_hd__a21o_1 _40858_ (.A1(_09926_),
    .A2(_13520_),
    .B1(_13522_),
    .X(_13524_));
 sky130_fd_sc_hd__nand3_1 _40859_ (.A(_13524_),
    .B(_13519_),
    .C(_09924_),
    .Y(_13525_));
 sky130_fd_sc_hd__a22oi_2 _40860_ (.A1(_08600_),
    .A2(_12330_),
    .B1(_13523_),
    .B2(_13525_),
    .Y(_13527_));
 sky130_fd_sc_hd__and4_1 _40861_ (.A(_08600_),
    .B(_12330_),
    .C(_13523_),
    .D(_13525_),
    .X(_13528_));
 sky130_fd_sc_hd__a2111oi_1 _40862_ (.A1(_11131_),
    .A2(_12327_),
    .B1(_02434_),
    .C1(_13527_),
    .D1(_13528_),
    .Y(_13529_));
 sky130_fd_sc_hd__and3_1 _40863_ (.A(_12327_),
    .B(_12324_),
    .C(_11131_),
    .X(_13530_));
 sky130_fd_sc_hd__o22a_1 _40864_ (.A1(_13530_),
    .A2(_02434_),
    .B1(_13527_),
    .B2(_13528_),
    .X(_13531_));
 sky130_fd_sc_hd__a21oi_1 _40865_ (.A1(_12325_),
    .A2(_12334_),
    .B1(_12333_),
    .Y(_13532_));
 sky130_fd_sc_hd__o21bai_1 _40866_ (.A1(net175),
    .A2(_13531_),
    .B1_N(_13532_),
    .Y(_13533_));
 sky130_fd_sc_hd__a2111o_1 _40867_ (.A1(_12325_),
    .A2(_12334_),
    .B1(net175),
    .C1(_13531_),
    .D1(_12333_),
    .X(_13534_));
 sky130_fd_sc_hd__a21boi_2 _40868_ (.A1(_13518_),
    .A2(_13533_),
    .B1_N(_13534_),
    .Y(_13535_));
 sky130_fd_sc_hd__o21ai_1 _40869_ (.A1(_13518_),
    .A2(_13533_),
    .B1(_13535_),
    .Y(_13536_));
 sky130_fd_sc_hd__o21ai_1 _40870_ (.A1(_11144_),
    .A2(_12336_),
    .B1(_11132_),
    .Y(_13538_));
 sky130_fd_sc_hd__nand2_1 _40871_ (.A(_12337_),
    .B(_13538_),
    .Y(_13539_));
 sky130_fd_sc_hd__xnor2_1 _40872_ (.A(_13536_),
    .B(_13539_),
    .Y(_13540_));
 sky130_fd_sc_hd__a21o_1 _40873_ (.A1(_12342_),
    .A2(_13517_),
    .B1(_13540_),
    .X(_13541_));
 sky130_fd_sc_hd__and3_1 _40874_ (.A(_11160_),
    .B(_11165_),
    .C(_12351_),
    .X(_13542_));
 sky130_fd_sc_hd__buf_1 _40875_ (.A(net389),
    .X(_13543_));
 sky130_fd_sc_hd__mux2_1 _40876_ (.A0(_13543_),
    .A1(_11164_),
    .S(net388),
    .X(_13544_));
 sky130_fd_sc_hd__buf_1 _40877_ (.A(_11164_),
    .X(_13545_));
 sky130_fd_sc_hd__and3_1 _40878_ (.A(_11157_),
    .B(_13545_),
    .C(_13543_),
    .X(_13546_));
 sky130_fd_sc_hd__a21o_1 _40879_ (.A1(_13545_),
    .A2(_13543_),
    .B1(_11157_),
    .X(_13547_));
 sky130_fd_sc_hd__and3b_1 _40880_ (.A_N(_13546_),
    .B(_13547_),
    .C(_13544_),
    .X(_13549_));
 sky130_fd_sc_hd__o21ba_1 _40881_ (.A1(_11157_),
    .A2(_13544_),
    .B1_N(_13549_),
    .X(_13550_));
 sky130_fd_sc_hd__o21a_1 _40882_ (.A1(_12356_),
    .A2(_13542_),
    .B1(_13550_),
    .X(_13551_));
 sky130_fd_sc_hd__buf_2 _40883_ (.A(_11160_),
    .X(_13552_));
 sky130_fd_sc_hd__a311o_1 _40884_ (.A1(_13552_),
    .A2(_11165_),
    .A3(_12351_),
    .B1(_12356_),
    .C1(_13550_),
    .X(_13553_));
 sky130_fd_sc_hd__or2b_1 _40885_ (.A(_13551_),
    .B_N(_13553_),
    .X(_13554_));
 sky130_fd_sc_hd__xnor2_1 _40886_ (.A(_12355_),
    .B(_13554_),
    .Y(_13555_));
 sky130_fd_sc_hd__a21oi_1 _40887_ (.A1(_12362_),
    .A2(_12365_),
    .B1(_13555_),
    .Y(_13556_));
 sky130_fd_sc_hd__and3_1 _40888_ (.A(_12362_),
    .B(_12365_),
    .C(_13555_),
    .X(_13557_));
 sky130_fd_sc_hd__nor2_1 _40889_ (.A(_13556_),
    .B(_13557_),
    .Y(_13558_));
 sky130_fd_sc_hd__o21a_1 _40890_ (.A1(_12367_),
    .A2(_12370_),
    .B1(_13558_),
    .X(_13560_));
 sky130_fd_sc_hd__nor3_1 _40891_ (.A(_12367_),
    .B(_12370_),
    .C(_13558_),
    .Y(_13561_));
 sky130_fd_sc_hd__nor2_1 _40892_ (.A(_13560_),
    .B(_13561_),
    .Y(_13562_));
 sky130_fd_sc_hd__nand3_2 _40893_ (.A(_12342_),
    .B(_13517_),
    .C(_13540_),
    .Y(_13563_));
 sky130_fd_sc_hd__nand3_1 _40894_ (.A(_13541_),
    .B(_13562_),
    .C(_13563_),
    .Y(_13564_));
 sky130_fd_sc_hd__a21o_1 _40895_ (.A1(_13563_),
    .A2(_13541_),
    .B1(_13562_),
    .X(_13565_));
 sky130_fd_sc_hd__a21o_1 _40896_ (.A1(_11094_),
    .A2(_12319_),
    .B1(_12316_),
    .X(_13566_));
 sky130_fd_sc_hd__buf_1 _40897_ (.A(_11096_),
    .X(_13567_));
 sky130_fd_sc_hd__buf_1 _40898_ (.A(_07214_),
    .X(_13568_));
 sky130_fd_sc_hd__or4b_1 _40899_ (.A(_13567_),
    .B(_13568_),
    .C(_12311_),
    .D_N(_11093_),
    .X(_13569_));
 sky130_fd_sc_hd__or2_1 _40900_ (.A(_11096_),
    .B(_07214_),
    .X(_13571_));
 sky130_fd_sc_hd__o21ai_1 _40901_ (.A1(_12311_),
    .A2(_11102_),
    .B1(_13571_),
    .Y(_13572_));
 sky130_fd_sc_hd__buf_1 _40902_ (.A(_11093_),
    .X(_13573_));
 sky130_fd_sc_hd__a21oi_1 _40903_ (.A1(_13571_),
    .A2(_13573_),
    .B1(_09971_),
    .Y(_13574_));
 sky130_fd_sc_hd__and3_1 _40904_ (.A(_13571_),
    .B(_11093_),
    .C(_09971_),
    .X(_13575_));
 sky130_fd_sc_hd__a211o_1 _40905_ (.A1(_13569_),
    .A2(_13572_),
    .B1(_13574_),
    .C1(_13575_),
    .X(_13576_));
 sky130_fd_sc_hd__o211ai_1 _40906_ (.A1(_13575_),
    .A2(_13574_),
    .B1(_13572_),
    .C1(_13569_),
    .Y(_13577_));
 sky130_fd_sc_hd__nor2_1 _40907_ (.A(_12310_),
    .B(_12312_),
    .Y(_13578_));
 sky130_fd_sc_hd__a221o_1 _40908_ (.A1(_13576_),
    .A2(_13577_),
    .B1(_12304_),
    .B2(_12313_),
    .C1(_13578_),
    .X(_13579_));
 sky130_fd_sc_hd__and2_1 _40909_ (.A(_12304_),
    .B(_12313_),
    .X(_13580_));
 sky130_fd_sc_hd__and2_1 _40910_ (.A(_13576_),
    .B(_13577_),
    .X(_13582_));
 sky130_fd_sc_hd__o21ai_1 _40911_ (.A1(_13578_),
    .A2(_13580_),
    .B1(_13582_),
    .Y(_13583_));
 sky130_fd_sc_hd__nand2_1 _40912_ (.A(_13579_),
    .B(_13583_),
    .Y(_13584_));
 sky130_fd_sc_hd__xnor2_1 _40913_ (.A(_12303_),
    .B(_13584_),
    .Y(_13585_));
 sky130_fd_sc_hd__and2_1 _40914_ (.A(_13566_),
    .B(_13585_),
    .X(_13586_));
 sky130_fd_sc_hd__nor2_1 _40915_ (.A(_13585_),
    .B(_13566_),
    .Y(_13587_));
 sky130_fd_sc_hd__or2_1 _40916_ (.A(_13586_),
    .B(_13587_),
    .X(_13588_));
 sky130_fd_sc_hd__inv_2 _40917_ (.A(_13588_),
    .Y(_13589_));
 sky130_fd_sc_hd__and2_1 _40918_ (.A(_12320_),
    .B(_12301_),
    .X(_13590_));
 sky130_fd_sc_hd__o21bai_2 _40919_ (.A1(_12321_),
    .A2(_12322_),
    .B1_N(_13590_),
    .Y(_13591_));
 sky130_fd_sc_hd__xor2_1 _40920_ (.A(_13589_),
    .B(_13591_),
    .X(_13593_));
 sky130_fd_sc_hd__a21o_1 _40921_ (.A1(_13564_),
    .A2(_13565_),
    .B1(_13593_),
    .X(_13594_));
 sky130_fd_sc_hd__nand3_2 _40922_ (.A(_13565_),
    .B(_13593_),
    .C(_13564_),
    .Y(_13595_));
 sky130_fd_sc_hd__o21ai_4 _40923_ (.A1(_12373_),
    .A2(_12377_),
    .B1(_12378_),
    .Y(_13596_));
 sky130_fd_sc_hd__a21oi_4 _40924_ (.A1(_13594_),
    .A2(_13595_),
    .B1(_13596_),
    .Y(_13597_));
 sky130_fd_sc_hd__nand3_4 _40925_ (.A(_13596_),
    .B(_13594_),
    .C(_13595_),
    .Y(_13598_));
 sky130_fd_sc_hd__or2b_1 _40926_ (.A(_13597_),
    .B_N(_13598_),
    .X(_13599_));
 sky130_fd_sc_hd__clkbuf_2 _40927_ (.A(_12222_),
    .X(_13600_));
 sky130_fd_sc_hd__nor2_1 _40928_ (.A(_12228_),
    .B(_11024_),
    .Y(_13601_));
 sky130_fd_sc_hd__and2_1 _40929_ (.A(_11024_),
    .B(_12228_),
    .X(_13602_));
 sky130_fd_sc_hd__nand2_1 _40930_ (.A(_11024_),
    .B(_08695_),
    .Y(_13604_));
 sky130_fd_sc_hd__o31a_1 _40931_ (.A1(_08695_),
    .A2(_13601_),
    .A3(_13602_),
    .B1(_13604_),
    .X(_13605_));
 sky130_fd_sc_hd__a21oi_1 _40932_ (.A1(_12232_),
    .A2(_12234_),
    .B1(_13605_),
    .Y(_13606_));
 sky130_fd_sc_hd__o311a_1 _40933_ (.A1(_08695_),
    .A2(_13601_),
    .A3(_13602_),
    .B1(_12237_),
    .C1(_13604_),
    .X(_13607_));
 sky130_fd_sc_hd__a211o_1 _40934_ (.A1(_12233_),
    .A2(_12239_),
    .B1(_13606_),
    .C1(_13607_),
    .X(_13608_));
 sky130_fd_sc_hd__o211ai_2 _40935_ (.A1(_13606_),
    .A2(_13607_),
    .B1(_12233_),
    .C1(_12239_),
    .Y(_13609_));
 sky130_fd_sc_hd__buf_1 _40936_ (.A(_12228_),
    .X(_13610_));
 sky130_fd_sc_hd__or3_1 _40937_ (.A(_13610_),
    .B(_12227_),
    .C(_11012_),
    .X(_13611_));
 sky130_fd_sc_hd__and4_1 _40938_ (.A(_13608_),
    .B(_12222_),
    .C(_13609_),
    .D(_13611_),
    .X(_13612_));
 sky130_fd_sc_hd__and3b_1 _40939_ (.A_N(_13610_),
    .B(_12222_),
    .C(_11011_),
    .X(_13613_));
 sky130_fd_sc_hd__o2bb2a_1 _40940_ (.A1_N(_13609_),
    .A2_N(_13608_),
    .B1(_13613_),
    .B2(_12227_),
    .X(_13615_));
 sky130_fd_sc_hd__o221ai_2 _40941_ (.A1(_12223_),
    .A2(_12243_),
    .B1(_13612_),
    .B2(_13615_),
    .C1(_12244_),
    .Y(_13616_));
 sky130_fd_sc_hd__or3b_1 _40942_ (.A(_12223_),
    .B(_12243_),
    .C_N(_12244_),
    .X(_13617_));
 sky130_fd_sc_hd__a211o_1 _40943_ (.A1(_12244_),
    .A2(_13617_),
    .B1(_13612_),
    .C1(_13615_),
    .X(_13618_));
 sky130_fd_sc_hd__o311a_1 _40944_ (.A1(_11013_),
    .A2(_12219_),
    .A3(_13600_),
    .B1(_13616_),
    .C1(_13618_),
    .X(_13619_));
 sky130_fd_sc_hd__a2111oi_1 _40945_ (.A1(_13616_),
    .A2(_13618_),
    .B1(_11013_),
    .C1(_12219_),
    .D1(_13600_),
    .Y(_13620_));
 sky130_fd_sc_hd__nor2_1 _40946_ (.A(_13619_),
    .B(_13620_),
    .Y(_13621_));
 sky130_fd_sc_hd__nand3_1 _40947_ (.A(_13621_),
    .B(_12250_),
    .C(_12248_),
    .Y(_13622_));
 sky130_fd_sc_hd__a21o_1 _40948_ (.A1(_12248_),
    .A2(_12250_),
    .B1(_13621_),
    .X(_13623_));
 sky130_fd_sc_hd__nand2_1 _40949_ (.A(_13622_),
    .B(_13623_),
    .Y(_13624_));
 sky130_fd_sc_hd__or3b_1 _40950_ (.A(_12252_),
    .B(_12255_),
    .C_N(_13624_),
    .X(_13626_));
 sky130_fd_sc_hd__o21bai_1 _40951_ (.A1(_12252_),
    .A2(_12255_),
    .B1_N(_13624_),
    .Y(_13627_));
 sky130_fd_sc_hd__and2_2 _40952_ (.A(_13626_),
    .B(_13627_),
    .X(_13628_));
 sky130_fd_sc_hd__a31oi_4 _40953_ (.A1(_11002_),
    .A2(_12177_),
    .A3(_12213_),
    .B1(_12211_),
    .Y(_13629_));
 sky130_fd_sc_hd__o221a_1 _40954_ (.A1(_07427_),
    .A2(_12199_),
    .B1(_10979_),
    .B2(_02589_),
    .C1(_07423_),
    .X(_13630_));
 sky130_fd_sc_hd__o21a_1 _40955_ (.A1(_12202_),
    .A2(_12195_),
    .B1(_12197_),
    .X(_13631_));
 sky130_fd_sc_hd__clkbuf_2 _40956_ (.A(_07416_),
    .X(_13632_));
 sky130_fd_sc_hd__or3b_1 _40957_ (.A(_07425_),
    .B(_13632_),
    .C_N(_12179_),
    .X(_13633_));
 sky130_fd_sc_hd__buf_1 _40958_ (.A(_05687_),
    .X(_13634_));
 sky130_fd_sc_hd__nor2_1 _40959_ (.A(_13634_),
    .B(_05688_),
    .Y(_13635_));
 sky130_fd_sc_hd__or2_1 _40960_ (.A(_09799_),
    .B(_13635_),
    .X(_13637_));
 sky130_fd_sc_hd__a21oi_2 _40961_ (.A1(_09803_),
    .A2(_12188_),
    .B1(_05691_),
    .Y(_13638_));
 sky130_fd_sc_hd__or3b_1 _40962_ (.A(_13634_),
    .B(_05688_),
    .C_N(_09799_),
    .X(_13639_));
 sky130_fd_sc_hd__and3_1 _40963_ (.A(_13637_),
    .B(_13638_),
    .C(_13639_),
    .X(_13640_));
 sky130_fd_sc_hd__a21oi_2 _40964_ (.A1(_13639_),
    .A2(_13637_),
    .B1(_13638_),
    .Y(_13641_));
 sky130_fd_sc_hd__a211o_1 _40965_ (.A1(_08736_),
    .A2(_13633_),
    .B1(_13640_),
    .C1(_13641_),
    .X(_13642_));
 sky130_fd_sc_hd__o221ai_4 _40966_ (.A1(_12183_),
    .A2(_13632_),
    .B1(_13641_),
    .B2(_13640_),
    .C1(_08736_),
    .Y(_13643_));
 sky130_fd_sc_hd__a211oi_2 _40967_ (.A1(_13642_),
    .A2(_13643_),
    .B1(_12180_),
    .C1(net220),
    .Y(_13644_));
 sky130_fd_sc_hd__o21a_1 _40968_ (.A1(_10980_),
    .A2(_10979_),
    .B1(_05697_),
    .X(_13645_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _40969_ (.A(_09799_),
    .X(_13646_));
 sky130_fd_sc_hd__a21o_1 _40970_ (.A1(_07423_),
    .A2(_13646_),
    .B1(_12199_),
    .X(_13648_));
 sky130_fd_sc_hd__o21ai_2 _40971_ (.A1(_12188_),
    .A2(_13645_),
    .B1(_13648_),
    .Y(_13649_));
 sky130_fd_sc_hd__o211ai_2 _40972_ (.A1(_12180_),
    .A2(net220),
    .B1(_13642_),
    .C1(_13643_),
    .Y(_13650_));
 sky130_fd_sc_hd__nand2_1 _40973_ (.A(_13649_),
    .B(_13650_),
    .Y(_13651_));
 sky130_fd_sc_hd__and2b_1 _40974_ (.A_N(_13644_),
    .B(_13650_),
    .X(_13652_));
 sky130_fd_sc_hd__o22a_1 _40975_ (.A1(_13644_),
    .A2(_13651_),
    .B1(_13649_),
    .B2(_13652_),
    .X(_13653_));
 sky130_fd_sc_hd__xor2_1 _40976_ (.A(_13631_),
    .B(_13653_),
    .X(_13654_));
 sky130_fd_sc_hd__xnor2_1 _40977_ (.A(_13630_),
    .B(_13654_),
    .Y(_13655_));
 sky130_fd_sc_hd__o311a_1 _40978_ (.A1(_10973_),
    .A2(_10994_),
    .A3(_12205_),
    .B1(_12206_),
    .C1(_13655_),
    .X(_13656_));
 sky130_fd_sc_hd__or3_1 _40979_ (.A(_10973_),
    .B(_10994_),
    .C(_12208_),
    .X(_13657_));
 sky130_fd_sc_hd__a21o_1 _40980_ (.A1(_12206_),
    .A2(_13657_),
    .B1(_13655_),
    .X(_13659_));
 sky130_fd_sc_hd__or2b_2 _40981_ (.A(_13656_),
    .B_N(_13659_),
    .X(_13660_));
 sky130_fd_sc_hd__xor2_4 _40982_ (.A(_13629_),
    .B(_13660_),
    .X(_13661_));
 sky130_fd_sc_hd__xnor2_4 _40983_ (.A(_13628_),
    .B(_13661_),
    .Y(_13662_));
 sky130_fd_sc_hd__nand3b_1 _40984_ (.A_N(_12279_),
    .B(_12280_),
    .C(_12282_),
    .Y(_13663_));
 sky130_fd_sc_hd__buf_1 _40985_ (.A(_09846_),
    .X(_13664_));
 sky130_fd_sc_hd__a21o_1 _40986_ (.A1(_11059_),
    .A2(_13664_),
    .B1(_09849_),
    .X(_13665_));
 sky130_fd_sc_hd__o21ai_1 _40987_ (.A1(_12260_),
    .A2(_12264_),
    .B1(_13665_),
    .Y(_13666_));
 sky130_fd_sc_hd__buf_1 _40988_ (.A(_07336_),
    .X(_13667_));
 sky130_fd_sc_hd__nand3b_1 _40989_ (.A_N(_08652_),
    .B(_11050_),
    .C(_07336_),
    .Y(_13668_));
 sky130_fd_sc_hd__or3b_1 _40990_ (.A(_05602_),
    .B(_05603_),
    .C_N(_04106_),
    .X(_13670_));
 sky130_fd_sc_hd__or2_1 _40991_ (.A(_09846_),
    .B(_07351_),
    .X(_13671_));
 sky130_fd_sc_hd__and4_1 _40992_ (.A(_05606_),
    .B(_12259_),
    .C(_13670_),
    .D(_13671_),
    .X(_13672_));
 sky130_fd_sc_hd__a22oi_1 _40993_ (.A1(_05606_),
    .A2(_12259_),
    .B1(_13670_),
    .B2(_13671_),
    .Y(_13673_));
 sky130_fd_sc_hd__a211oi_1 _40994_ (.A1(_08658_),
    .A2(_13668_),
    .B1(_13672_),
    .C1(_13673_),
    .Y(_13674_));
 sky130_fd_sc_hd__o211a_1 _40995_ (.A1(_13672_),
    .A2(_13673_),
    .B1(_08658_),
    .C1(_13668_),
    .X(_13675_));
 sky130_fd_sc_hd__o221a_1 _40996_ (.A1(_13667_),
    .A2(_11052_),
    .B1(_13674_),
    .B2(_13675_),
    .C1(_12269_),
    .X(_13676_));
 sky130_fd_sc_hd__o2bb2a_1 _40997_ (.A1_N(_12265_),
    .A2_N(_12267_),
    .B1(_13667_),
    .B2(_11052_),
    .X(_13677_));
 sky130_fd_sc_hd__or3_1 _40998_ (.A(_13674_),
    .B(_13675_),
    .C(_13677_),
    .X(_13678_));
 sky130_fd_sc_hd__and2b_1 _40999_ (.A_N(_13676_),
    .B(_13678_),
    .X(_13679_));
 sky130_fd_sc_hd__and2_1 _41000_ (.A(_13666_),
    .B(_13678_),
    .X(_13681_));
 sky130_fd_sc_hd__inv_2 _41001_ (.A(_13681_),
    .Y(_13682_));
 sky130_fd_sc_hd__o22a_1 _41002_ (.A1(_13666_),
    .A2(_13679_),
    .B1(_13676_),
    .B2(_13682_),
    .X(_13683_));
 sky130_fd_sc_hd__a21oi_1 _41003_ (.A1(_12271_),
    .A2(_12278_),
    .B1(_13683_),
    .Y(_13684_));
 sky130_fd_sc_hd__and3_1 _41004_ (.A(_13683_),
    .B(_12278_),
    .C(_12271_),
    .X(_13685_));
 sky130_fd_sc_hd__nor2_1 _41005_ (.A(_13684_),
    .B(_13685_),
    .Y(_13686_));
 sky130_fd_sc_hd__o221a_1 _41006_ (.A1(_08644_),
    .A2(_09853_),
    .B1(_11057_),
    .B2(_11058_),
    .C1(_13686_),
    .X(_13687_));
 sky130_fd_sc_hd__buf_1 _41007_ (.A(_09849_),
    .X(_13688_));
 sky130_fd_sc_hd__o221a_1 _41008_ (.A1(_09865_),
    .A2(_13688_),
    .B1(_11057_),
    .B2(_11058_),
    .C1(_11069_),
    .X(_13689_));
 sky130_fd_sc_hd__nor2_1 _41009_ (.A(_13689_),
    .B(_13686_),
    .Y(_13690_));
 sky130_fd_sc_hd__or2_1 _41010_ (.A(_13687_),
    .B(_13690_),
    .X(_13692_));
 sky130_fd_sc_hd__and3_1 _41011_ (.A(_12280_),
    .B(_13663_),
    .C(_13692_),
    .X(_13693_));
 sky130_fd_sc_hd__a21o_1 _41012_ (.A1(_12280_),
    .A2(_13663_),
    .B1(_13692_),
    .X(_13694_));
 sky130_fd_sc_hd__and2b_1 _41013_ (.A_N(_13693_),
    .B(_13694_),
    .X(_13695_));
 sky130_fd_sc_hd__a31oi_4 _41014_ (.A1(_11083_),
    .A2(_12290_),
    .A3(_12287_),
    .B1(_12285_),
    .Y(_13696_));
 sky130_fd_sc_hd__xor2_4 _41015_ (.A(_13695_),
    .B(_13696_),
    .X(_13697_));
 sky130_fd_sc_hd__xnor2_4 _41016_ (.A(_13662_),
    .B(_13697_),
    .Y(_13698_));
 sky130_fd_sc_hd__xnor2_2 _41017_ (.A(_13599_),
    .B(_13698_),
    .Y(_13699_));
 sky130_fd_sc_hd__a21oi_4 _41018_ (.A1(_12380_),
    .A2(_12382_),
    .B1(_13699_),
    .Y(_13700_));
 sky130_fd_sc_hd__and3_4 _41019_ (.A(_13699_),
    .B(_12382_),
    .C(_12380_),
    .X(_13701_));
 sky130_fd_sc_hd__o22a_1 _41020_ (.A1(_13514_),
    .A2(_13516_),
    .B1(_13700_),
    .B2(_13701_),
    .X(_13703_));
 sky130_fd_sc_hd__nor4_1 _41021_ (.A(_13514_),
    .B(_13516_),
    .C(_13700_),
    .D(_13701_),
    .Y(_13704_));
 sky130_fd_sc_hd__a211oi_1 _41022_ (.A1(_12495_),
    .A2(_12385_),
    .B1(_13703_),
    .C1(net73),
    .Y(_13705_));
 sky130_fd_sc_hd__o221a_1 _41023_ (.A1(_12492_),
    .A2(_12494_),
    .B1(_13703_),
    .B2(net73),
    .C1(_12385_),
    .X(_13706_));
 sky130_fd_sc_hd__o22a_1 _41024_ (.A1(_13423_),
    .A2(_13424_),
    .B1(_13705_),
    .B2(_13706_),
    .X(_13707_));
 sky130_fd_sc_hd__nor4_1 _41025_ (.A(_13423_),
    .B(_13424_),
    .C(_13705_),
    .D(_13706_),
    .Y(_13708_));
 sky130_fd_sc_hd__a21o_1 _41026_ (.A1(_12615_),
    .A2(_12499_),
    .B1(_12498_),
    .X(_13709_));
 sky130_fd_sc_hd__o21bai_1 _41027_ (.A1(_13707_),
    .A2(_13708_),
    .B1_N(_13709_),
    .Y(_13710_));
 sky130_fd_sc_hd__or3b_2 _41028_ (.A(_13707_),
    .B(_13708_),
    .C_N(_13709_),
    .X(_13711_));
 sky130_fd_sc_hd__nand2_2 _41029_ (.A(_13710_),
    .B(_13711_),
    .Y(_13712_));
 sky130_fd_sc_hd__or2b_1 _41030_ (.A(_12733_),
    .B_N(_12731_),
    .X(_13714_));
 sky130_fd_sc_hd__and3_1 _41031_ (.A(_12503_),
    .B(_12609_),
    .C(_12610_),
    .X(_13715_));
 sky130_fd_sc_hd__a221o_1 _41032_ (.A1(_11308_),
    .A2(_11310_),
    .B1(_12609_),
    .B2(_12610_),
    .C1(_11307_),
    .X(_13716_));
 sky130_fd_sc_hd__and2b_1 _41033_ (.A_N(_12502_),
    .B(_13716_),
    .X(_13717_));
 sky130_fd_sc_hd__or2b_1 _41034_ (.A(_11524_),
    .B_N(_09582_),
    .X(_13718_));
 sky130_fd_sc_hd__or2b_1 _41035_ (.A(_09582_),
    .B_N(_11524_),
    .X(_13719_));
 sky130_fd_sc_hd__a22o_1 _41036_ (.A1(_09586_),
    .A2(_12633_),
    .B1(_13718_),
    .B2(_13719_),
    .X(_13720_));
 sky130_fd_sc_hd__nand4_2 _41037_ (.A(_09586_),
    .B(_13718_),
    .C(_13719_),
    .D(_12633_),
    .Y(_13721_));
 sky130_fd_sc_hd__and3_1 _41038_ (.A(_13720_),
    .B(_12640_),
    .C(_13721_),
    .X(_13722_));
 sky130_fd_sc_hd__a21oi_1 _41039_ (.A1(_13721_),
    .A2(_13720_),
    .B1(_12640_),
    .Y(_13723_));
 sky130_fd_sc_hd__and4bb_1 _41040_ (.A_N(_13722_),
    .B_N(_13723_),
    .C(_12634_),
    .D(_12635_),
    .X(_13725_));
 sky130_fd_sc_hd__o2bb2a_1 _41041_ (.A1_N(_12634_),
    .A2_N(_12635_),
    .B1(_13722_),
    .B2(_13723_),
    .X(_13726_));
 sky130_fd_sc_hd__a211oi_2 _41042_ (.A1(_12641_),
    .A2(_12642_),
    .B1(_13725_),
    .C1(_13726_),
    .Y(_13727_));
 sky130_fd_sc_hd__o211a_1 _41043_ (.A1(_13725_),
    .A2(_13726_),
    .B1(_12641_),
    .C1(_12642_),
    .X(_13728_));
 sky130_fd_sc_hd__nor4_1 _41044_ (.A(_13727_),
    .B(_12644_),
    .C(_12645_),
    .D(_13728_),
    .Y(_13729_));
 sky130_fd_sc_hd__o22a_1 _41045_ (.A1(_13727_),
    .A2(_13728_),
    .B1(_12644_),
    .B2(_12645_),
    .X(_13730_));
 sky130_fd_sc_hd__o221ai_4 _41046_ (.A1(_12650_),
    .A2(_12652_),
    .B1(net150),
    .B2(_13730_),
    .C1(_12655_),
    .Y(_13731_));
 sky130_fd_sc_hd__or2_1 _41047_ (.A(net151),
    .B(_13730_),
    .X(_13732_));
 sky130_fd_sc_hd__a21o_1 _41048_ (.A1(_12653_),
    .A2(_12655_),
    .B1(_13732_),
    .X(_13733_));
 sky130_fd_sc_hd__o21ai_1 _41049_ (.A1(_11518_),
    .A2(_11521_),
    .B1(_12678_),
    .Y(_13734_));
 sky130_fd_sc_hd__nor3_1 _41050_ (.A(_12666_),
    .B(_12667_),
    .C(_12670_),
    .Y(_13736_));
 sky130_fd_sc_hd__and2_1 _41051_ (.A(_12671_),
    .B(_12656_),
    .X(_13737_));
 sky130_fd_sc_hd__clkbuf_2 _41052_ (.A(_09619_),
    .X(_13738_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41053_ (.A(_12660_),
    .X(_13739_));
 sky130_fd_sc_hd__buf_1 _41054_ (.A(_12659_),
    .X(_13740_));
 sky130_fd_sc_hd__and3_1 _41055_ (.A(_09633_),
    .B(_13739_),
    .C(_13740_),
    .X(_13741_));
 sky130_fd_sc_hd__a41o_1 _41056_ (.A1(_06812_),
    .A2(_12657_),
    .A3(_12661_),
    .A4(_13738_),
    .B1(_13741_),
    .X(_13742_));
 sky130_fd_sc_hd__and3b_1 _41057_ (.A_N(_12660_),
    .B(_12659_),
    .C(_12664_),
    .X(_13743_));
 sky130_fd_sc_hd__and2_1 _41058_ (.A(_11496_),
    .B(_12660_),
    .X(_13744_));
 sky130_fd_sc_hd__xnor2_1 _41059_ (.A(_09619_),
    .B(_12659_),
    .Y(_13745_));
 sky130_fd_sc_hd__xor2_1 _41060_ (.A(_13744_),
    .B(_13745_),
    .X(_13747_));
 sky130_fd_sc_hd__o21a_1 _41061_ (.A1(_12666_),
    .A2(_13743_),
    .B1(_13747_),
    .X(_13748_));
 sky130_fd_sc_hd__a311oi_1 _41062_ (.A1(_12662_),
    .A2(_12663_),
    .A3(_12665_),
    .B1(_13747_),
    .C1(_13743_),
    .Y(_13749_));
 sky130_fd_sc_hd__nor2_1 _41063_ (.A(_13748_),
    .B(_13749_),
    .Y(_13750_));
 sky130_fd_sc_hd__xor2_1 _41064_ (.A(_13742_),
    .B(_13750_),
    .X(_13751_));
 sky130_fd_sc_hd__o21ai_1 _41065_ (.A1(_13736_),
    .A2(_13737_),
    .B1(_13751_),
    .Y(_13752_));
 sky130_fd_sc_hd__or3_1 _41066_ (.A(_13736_),
    .B(_13737_),
    .C(_13751_),
    .X(_13753_));
 sky130_fd_sc_hd__and2_1 _41067_ (.A(_13752_),
    .B(_13753_),
    .X(_13754_));
 sky130_fd_sc_hd__xor2_1 _41068_ (.A(_12673_),
    .B(_13754_),
    .X(_13755_));
 sky130_fd_sc_hd__a21oi_1 _41069_ (.A1(_11516_),
    .A2(_12676_),
    .B1(_13755_),
    .Y(_13756_));
 sky130_fd_sc_hd__o21a_1 _41070_ (.A1(net125),
    .A2(_12679_),
    .B1(_13755_),
    .X(_13758_));
 sky130_fd_sc_hd__a21oi_1 _41071_ (.A1(_13734_),
    .A2(_13756_),
    .B1(_13758_),
    .Y(_13759_));
 sky130_fd_sc_hd__nand3_1 _41072_ (.A(_13731_),
    .B(_13733_),
    .C(_13759_),
    .Y(_13760_));
 sky130_fd_sc_hd__a21o_1 _41073_ (.A1(_13731_),
    .A2(_13733_),
    .B1(_13759_),
    .X(_13761_));
 sky130_fd_sc_hd__nand2_1 _41074_ (.A(_13760_),
    .B(_13761_),
    .Y(_13762_));
 sky130_fd_sc_hd__or2_1 _41075_ (.A(_11480_),
    .B(net177),
    .X(_13763_));
 sky130_fd_sc_hd__o211ai_1 _41076_ (.A1(_11477_),
    .A2(_06780_),
    .B1(_06785_),
    .C1(_12623_),
    .Y(_13764_));
 sky130_fd_sc_hd__o31a_1 _41077_ (.A1(_06785_),
    .A2(_11477_),
    .A3(_06780_),
    .B1(_13764_),
    .X(_13765_));
 sky130_fd_sc_hd__a31oi_1 _41078_ (.A1(_12624_),
    .A2(_12626_),
    .A3(_13763_),
    .B1(_13765_),
    .Y(_13766_));
 sky130_fd_sc_hd__a21boi_4 _41079_ (.A1(_12628_),
    .A2(_12630_),
    .B1_N(_13765_),
    .Y(_13767_));
 sky130_fd_sc_hd__a21oi_1 _41080_ (.A1(_12630_),
    .A2(_13766_),
    .B1(_13767_),
    .Y(_13769_));
 sky130_fd_sc_hd__inv_2 _41081_ (.A(_13769_),
    .Y(_13770_));
 sky130_fd_sc_hd__and3_1 _41082_ (.A(_13760_),
    .B(_13770_),
    .C(_13761_),
    .X(_13771_));
 sky130_fd_sc_hd__a2111o_1 _41083_ (.A1(_13762_),
    .A2(_13769_),
    .B1(_12555_),
    .C1(_12542_),
    .D1(_13771_),
    .X(_13772_));
 sky130_fd_sc_hd__inv_2 _41084_ (.A(_13760_),
    .Y(_13773_));
 sky130_fd_sc_hd__nor2_1 _41085_ (.A(_13773_),
    .B(_13770_),
    .Y(_13774_));
 sky130_fd_sc_hd__o21a_1 _41086_ (.A1(_12540_),
    .A2(_12553_),
    .B1(_12541_),
    .X(_13775_));
 sky130_fd_sc_hd__a221o_1 _41087_ (.A1(_13770_),
    .A2(_13762_),
    .B1(_13774_),
    .B2(_13761_),
    .C1(_13775_),
    .X(_13776_));
 sky130_fd_sc_hd__o21ai_1 _41088_ (.A1(_12632_),
    .A2(_12685_),
    .B1(_12683_),
    .Y(_13777_));
 sky130_fd_sc_hd__a21o_1 _41089_ (.A1(_13772_),
    .A2(_13776_),
    .B1(_13777_),
    .X(_13778_));
 sky130_fd_sc_hd__nand3_2 _41090_ (.A(_13777_),
    .B(_13772_),
    .C(_13776_),
    .Y(_13780_));
 sky130_fd_sc_hd__o21ai_1 _41091_ (.A1(_12687_),
    .A2(_12690_),
    .B1(_12693_),
    .Y(_13781_));
 sky130_fd_sc_hd__a21o_1 _41092_ (.A1(_13778_),
    .A2(_13780_),
    .B1(_13781_),
    .X(_13782_));
 sky130_fd_sc_hd__nand3_2 _41093_ (.A(_13781_),
    .B(_13778_),
    .C(_13780_),
    .Y(_13783_));
 sky130_fd_sc_hd__nand2_1 _41094_ (.A(_13782_),
    .B(_13783_),
    .Y(_13784_));
 sky130_fd_sc_hd__o21ai_1 _41095_ (.A1(_12699_),
    .A2(_12704_),
    .B1(_12700_),
    .Y(_13785_));
 sky130_fd_sc_hd__or4_1 _41096_ (.A(_11569_),
    .B(_11571_),
    .C(_12707_),
    .D(_09698_),
    .X(_13786_));
 sky130_fd_sc_hd__mux2_1 _41097_ (.A0(_08251_),
    .A1(_06682_),
    .S(_03704_),
    .X(_13787_));
 sky130_fd_sc_hd__o2111a_1 _41098_ (.A1(_12706_),
    .A2(_12709_),
    .B1(_12710_),
    .C1(_13786_),
    .D1(_13787_),
    .X(_13788_));
 sky130_fd_sc_hd__o211a_1 _41099_ (.A1(_12706_),
    .A2(_12709_),
    .B1(_12710_),
    .C1(_13786_),
    .X(_13789_));
 sky130_fd_sc_hd__nor2_1 _41100_ (.A(_13789_),
    .B(_13787_),
    .Y(_13791_));
 sky130_fd_sc_hd__or3_2 _41101_ (.A(_13785_),
    .B(_13788_),
    .C(_13791_),
    .X(_13792_));
 sky130_fd_sc_hd__o21ai_1 _41102_ (.A1(_13788_),
    .A2(_13791_),
    .B1(_13785_),
    .Y(_13793_));
 sky130_fd_sc_hd__and3_1 _41103_ (.A(_12696_),
    .B(_13792_),
    .C(_13793_),
    .X(_13794_));
 sky130_fd_sc_hd__a21oi_1 _41104_ (.A1(_13792_),
    .A2(_13793_),
    .B1(_12696_),
    .Y(_13795_));
 sky130_fd_sc_hd__nand2_1 _41105_ (.A(_11580_),
    .B(_12715_),
    .Y(_13796_));
 sky130_fd_sc_hd__o211a_1 _41106_ (.A1(_13794_),
    .A2(_13795_),
    .B1(_12714_),
    .C1(_13796_),
    .X(_13797_));
 sky130_fd_sc_hd__a211oi_2 _41107_ (.A1(_12714_),
    .A2(_13796_),
    .B1(_13794_),
    .C1(_13795_),
    .Y(_13798_));
 sky130_fd_sc_hd__or2_1 _41108_ (.A(_13797_),
    .B(_13798_),
    .X(_13799_));
 sky130_fd_sc_hd__and2_1 _41109_ (.A(_11588_),
    .B(_12725_),
    .X(_13800_));
 sky130_fd_sc_hd__nor2_1 _41110_ (.A(_11588_),
    .B(_12727_),
    .Y(_13802_));
 sky130_fd_sc_hd__or2_2 _41111_ (.A(_13800_),
    .B(_13802_),
    .X(_13803_));
 sky130_fd_sc_hd__nor2_1 _41112_ (.A(_13799_),
    .B(_13803_),
    .Y(_13804_));
 sky130_fd_sc_hd__o21a_1 _41113_ (.A1(_13800_),
    .A2(_13802_),
    .B1(_13799_),
    .X(_13805_));
 sky130_fd_sc_hd__nor2_2 _41114_ (.A(_13804_),
    .B(_13805_),
    .Y(_13806_));
 sky130_fd_sc_hd__xnor2_1 _41115_ (.A(_13784_),
    .B(_13806_),
    .Y(_13807_));
 sky130_fd_sc_hd__o21a_1 _41116_ (.A1(_13715_),
    .A2(_13717_),
    .B1(_13807_),
    .X(_13808_));
 sky130_fd_sc_hd__nor3_1 _41117_ (.A(_13715_),
    .B(_13717_),
    .C(_13807_),
    .Y(_13809_));
 sky130_fd_sc_hd__nor2_1 _41118_ (.A(_13808_),
    .B(_13809_),
    .Y(_13810_));
 sky130_fd_sc_hd__nor2_1 _41119_ (.A(_13714_),
    .B(_13810_),
    .Y(_13811_));
 sky130_fd_sc_hd__and2_1 _41120_ (.A(_13810_),
    .B(_13714_),
    .X(_13813_));
 sky130_fd_sc_hd__nor2_1 _41121_ (.A(_13811_),
    .B(_13813_),
    .Y(_13814_));
 sky130_fd_sc_hd__xor2_2 _41122_ (.A(_13712_),
    .B(_13814_),
    .X(_13815_));
 sky130_fd_sc_hd__a21boi_2 _41123_ (.A1(_12173_),
    .A2(_12616_),
    .B1_N(_12743_),
    .Y(_13816_));
 sky130_fd_sc_hd__xor2_2 _41124_ (.A(_13815_),
    .B(_13816_),
    .X(_13817_));
 sky130_fd_sc_hd__a21o_1 _41125_ (.A1(_13305_),
    .A2(_13308_),
    .B1(_13817_),
    .X(_13818_));
 sky130_fd_sc_hd__nand3_1 _41126_ (.A(_13305_),
    .B(_13308_),
    .C(_13817_),
    .Y(_13819_));
 sky130_fd_sc_hd__nand3_1 _41127_ (.A(_12873_),
    .B(_13818_),
    .C(_13819_),
    .Y(_13820_));
 sky130_fd_sc_hd__buf_1 _41128_ (.A(_13820_),
    .X(_13821_));
 sky130_fd_sc_hd__a21oi_1 _41129_ (.A1(_13305_),
    .A2(_13308_),
    .B1(_13817_),
    .Y(_13822_));
 sky130_fd_sc_hd__and3_1 _41130_ (.A(_13305_),
    .B(_13817_),
    .C(_13308_),
    .X(_13824_));
 sky130_fd_sc_hd__a31oi_1 _41131_ (.A1(_12751_),
    .A2(_12748_),
    .A3(_12750_),
    .B1(_12747_),
    .Y(_13825_));
 sky130_fd_sc_hd__o21ai_1 _41132_ (.A1(_13822_),
    .A2(_13824_),
    .B1(_13825_),
    .Y(_13826_));
 sky130_fd_sc_hd__clkbuf_2 _41133_ (.A(_13826_),
    .X(_13827_));
 sky130_fd_sc_hd__a21oi_1 _41134_ (.A1(_12159_),
    .A2(_12161_),
    .B1(_12162_),
    .Y(_13828_));
 sky130_fd_sc_hd__a31oi_2 _41135_ (.A1(_12159_),
    .A2(_12161_),
    .A3(_12162_),
    .B1(_12171_),
    .Y(_13829_));
 sky130_fd_sc_hd__or3b_2 _41136_ (.A(_08982_),
    .B(_08975_),
    .C_N(_10467_),
    .X(_13830_));
 sky130_fd_sc_hd__or2_1 _41137_ (.A(_08967_),
    .B(_12762_),
    .X(_13831_));
 sky130_fd_sc_hd__and2_1 _41138_ (.A(_04533_),
    .B(_10302_),
    .X(_13832_));
 sky130_fd_sc_hd__nor2_2 _41139_ (.A(_10302_),
    .B(_04533_),
    .Y(_13833_));
 sky130_fd_sc_hd__o211ai_1 _41140_ (.A1(_03033_),
    .A2(_08974_),
    .B1(_12765_),
    .C1(_12766_),
    .Y(_13835_));
 sky130_fd_sc_hd__o2111ai_1 _41141_ (.A1(_08973_),
    .A2(_09000_),
    .B1(_12765_),
    .C1(_13835_),
    .D1(_10304_),
    .Y(_13836_));
 sky130_fd_sc_hd__or2_1 _41142_ (.A(_08973_),
    .B(_09000_),
    .X(_13837_));
 sky130_fd_sc_hd__a22o_1 _41143_ (.A1(_12765_),
    .A2(_13835_),
    .B1(_13837_),
    .B2(_10304_),
    .X(_13838_));
 sky130_fd_sc_hd__or4bb_2 _41144_ (.A(_13832_),
    .B(_13833_),
    .C_N(_13836_),
    .D_N(_13838_),
    .X(_13839_));
 sky130_fd_sc_hd__a2bb2o_1 _41145_ (.A1_N(_13832_),
    .A2_N(_13833_),
    .B1(_13836_),
    .B2(_13838_),
    .X(_13840_));
 sky130_fd_sc_hd__a211o_1 _41146_ (.A1(_13839_),
    .A2(_13840_),
    .B1(_12771_),
    .C1(net163),
    .X(_13841_));
 sky130_fd_sc_hd__o211ai_4 _41147_ (.A1(_12771_),
    .A2(net163),
    .B1(_13839_),
    .C1(_13840_),
    .Y(_13842_));
 sky130_fd_sc_hd__a22o_2 _41148_ (.A1(_13830_),
    .A2(_13831_),
    .B1(_13841_),
    .B2(_13842_),
    .X(_13843_));
 sky130_fd_sc_hd__clkbuf_2 _41149_ (.A(_24238_),
    .X(_13844_));
 sky130_fd_sc_hd__a21boi_2 _41150_ (.A1(_24256_),
    .A2(_13844_),
    .B1_N(_10436_),
    .Y(_13846_));
 sky130_fd_sc_hd__and4b_1 _41151_ (.A_N(_10436_),
    .B(_00437_),
    .C(_24238_),
    .D(_06644_),
    .X(_13847_));
 sky130_fd_sc_hd__and3_1 _41152_ (.A(_12150_),
    .B(_12155_),
    .C(_12156_),
    .X(_13848_));
 sky130_fd_sc_hd__or4_1 _41153_ (.A(_12154_),
    .B(_13846_),
    .C(_13847_),
    .D(_13848_),
    .X(_13849_));
 sky130_fd_sc_hd__o22ai_2 _41154_ (.A1(_13846_),
    .A2(_13847_),
    .B1(_13848_),
    .B2(_12154_),
    .Y(_13850_));
 sky130_fd_sc_hd__and3_1 _41155_ (.A(_13849_),
    .B(_12785_),
    .C(_13850_),
    .X(_13851_));
 sky130_fd_sc_hd__a21oi_1 _41156_ (.A1(_13850_),
    .A2(_13849_),
    .B1(_12785_),
    .Y(_13852_));
 sky130_fd_sc_hd__or2_2 _41157_ (.A(_13851_),
    .B(_13852_),
    .X(_13853_));
 sky130_fd_sc_hd__a21boi_2 _41158_ (.A1(_12788_),
    .A2(_12787_),
    .B1_N(_12786_),
    .Y(_13854_));
 sky130_fd_sc_hd__xor2_1 _41159_ (.A(_13853_),
    .B(_13854_),
    .X(_13855_));
 sky130_fd_sc_hd__nand4_4 _41160_ (.A(_13830_),
    .B(_13831_),
    .C(_13841_),
    .D(_13842_),
    .Y(_13857_));
 sky130_fd_sc_hd__nand3_1 _41161_ (.A(_13843_),
    .B(_13855_),
    .C(_13857_),
    .Y(_13858_));
 sky130_fd_sc_hd__a21o_1 _41162_ (.A1(_13857_),
    .A2(_13843_),
    .B1(_13855_),
    .X(_13859_));
 sky130_fd_sc_hd__nand2_1 _41163_ (.A(_13858_),
    .B(_13859_),
    .Y(_13860_));
 sky130_fd_sc_hd__o21bai_4 _41164_ (.A1(_13828_),
    .A2(_13829_),
    .B1_N(_13860_),
    .Y(_13861_));
 sky130_fd_sc_hd__o21ai_1 _41165_ (.A1(_11699_),
    .A2(_11700_),
    .B1(_12164_),
    .Y(_13862_));
 sky130_fd_sc_hd__nand3_1 _41166_ (.A(_12169_),
    .B(_13862_),
    .C(_13860_),
    .Y(_13863_));
 sky130_fd_sc_hd__a21bo_1 _41167_ (.A1(_12780_),
    .A2(_12792_),
    .B1_N(_12793_),
    .X(_13864_));
 sky130_fd_sc_hd__a21o_1 _41168_ (.A1(_13861_),
    .A2(_13863_),
    .B1(_13864_),
    .X(_13865_));
 sky130_fd_sc_hd__nand3_1 _41169_ (.A(_13864_),
    .B(_13861_),
    .C(_13863_),
    .Y(_13866_));
 sky130_fd_sc_hd__nand4_1 _41170_ (.A(_13821_),
    .B(_13827_),
    .C(_13865_),
    .D(_13866_),
    .Y(_13868_));
 sky130_fd_sc_hd__and2_1 _41171_ (.A(_13865_),
    .B(_13866_),
    .X(_13869_));
 sky130_fd_sc_hd__a21o_1 _41172_ (.A1(_13821_),
    .A2(_13827_),
    .B1(_13869_),
    .X(_13870_));
 sky130_fd_sc_hd__nand3_1 _41173_ (.A(_12872_),
    .B(_13868_),
    .C(_13870_),
    .Y(_13871_));
 sky130_fd_sc_hd__nand2_1 _41174_ (.A(_13865_),
    .B(_13866_),
    .Y(_13872_));
 sky130_fd_sc_hd__a21o_1 _41175_ (.A1(_13820_),
    .A2(_13826_),
    .B1(_13872_),
    .X(_13873_));
 sky130_fd_sc_hd__nand3_1 _41176_ (.A(_13821_),
    .B(_13827_),
    .C(_13872_),
    .Y(_13874_));
 sky130_fd_sc_hd__nand3b_2 _41177_ (.A_N(_12872_),
    .B(_13873_),
    .C(_13874_),
    .Y(_13875_));
 sky130_fd_sc_hd__o31ai_4 _41178_ (.A1(_10468_),
    .A2(_12824_),
    .A3(_12825_),
    .B1(_12828_),
    .Y(_13876_));
 sky130_fd_sc_hd__o21a_1 _41179_ (.A1(_25242_),
    .A2(_25240_),
    .B1(_08956_),
    .X(_13877_));
 sky130_fd_sc_hd__a21boi_2 _41180_ (.A1(_25247_),
    .A2(_25251_),
    .B1_N(_07507_),
    .Y(_13879_));
 sky130_fd_sc_hd__and3b_1 _41181_ (.A_N(_08959_),
    .B(_25247_),
    .C(_25251_),
    .X(_13880_));
 sky130_fd_sc_hd__o22a_1 _41182_ (.A1(_23724_),
    .A2(_13877_),
    .B1(_13879_),
    .B2(_13880_),
    .X(_13881_));
 sky130_fd_sc_hd__a2111oi_1 _41183_ (.A1(_25242_),
    .A2(_07597_),
    .B1(_13877_),
    .C1(_13879_),
    .D1(_13880_),
    .Y(_13882_));
 sky130_fd_sc_hd__and4bb_1 _41184_ (.A_N(_13881_),
    .B_N(net243),
    .C(_08966_),
    .D(_10461_),
    .X(_13883_));
 sky130_fd_sc_hd__inv_2 _41185_ (.A(_13883_),
    .Y(_13884_));
 sky130_fd_sc_hd__a2bb2o_1 _41186_ (.A1_N(_13881_),
    .A2_N(net243),
    .B1(_10297_),
    .B2(_10461_),
    .X(_13885_));
 sky130_fd_sc_hd__nand3_1 _41187_ (.A(_13884_),
    .B(_13885_),
    .C(_12824_),
    .Y(_13886_));
 sky130_fd_sc_hd__a21o_1 _41188_ (.A1(_13884_),
    .A2(_13885_),
    .B1(_12824_),
    .X(_13887_));
 sky130_fd_sc_hd__a211oi_1 _41189_ (.A1(_10458_),
    .A2(_12774_),
    .B1(_12772_),
    .C1(_12773_),
    .Y(_13888_));
 sky130_fd_sc_hd__a211oi_1 _41190_ (.A1(_13886_),
    .A2(_13887_),
    .B1(_13888_),
    .C1(_12777_),
    .Y(_13890_));
 sky130_fd_sc_hd__o211a_1 _41191_ (.A1(_13888_),
    .A2(_12777_),
    .B1(_13886_),
    .C1(_13887_),
    .X(_13891_));
 sky130_fd_sc_hd__nor2_2 _41192_ (.A(_13890_),
    .B(_13891_),
    .Y(_13892_));
 sky130_fd_sc_hd__xnor2_2 _41193_ (.A(_13876_),
    .B(_13892_),
    .Y(_13893_));
 sky130_fd_sc_hd__and3_1 _41194_ (.A(_12831_),
    .B(_12835_),
    .C(_13893_),
    .X(_13894_));
 sky130_fd_sc_hd__a21oi_4 _41195_ (.A1(_12831_),
    .A2(_12835_),
    .B1(_13893_),
    .Y(_13895_));
 sky130_fd_sc_hd__nor2_2 _41196_ (.A(_13894_),
    .B(_13895_),
    .Y(_13896_));
 sky130_fd_sc_hd__a21oi_1 _41197_ (.A1(_10967_),
    .A2(_11624_),
    .B1(_12796_),
    .Y(_13897_));
 sky130_fd_sc_hd__a211oi_1 _41198_ (.A1(_12800_),
    .A2(_12799_),
    .B1(_13896_),
    .C1(_13897_),
    .Y(_13898_));
 sky130_fd_sc_hd__o21a_1 _41199_ (.A1(_12797_),
    .A2(_12759_),
    .B1(_12800_),
    .X(_13899_));
 sky130_fd_sc_hd__o21ai_1 _41200_ (.A1(_13897_),
    .A2(_13899_),
    .B1(_13896_),
    .Y(_13901_));
 sky130_fd_sc_hd__and2b_1 _41201_ (.A_N(_13898_),
    .B(_13901_),
    .X(_13902_));
 sky130_fd_sc_hd__xnor2_2 _41202_ (.A(_12838_),
    .B(_13902_),
    .Y(_13903_));
 sky130_fd_sc_hd__a21o_1 _41203_ (.A1(_13871_),
    .A2(_13875_),
    .B1(_13903_),
    .X(_13904_));
 sky130_fd_sc_hd__a32oi_4 _41204_ (.A1(_12816_),
    .A2(_12817_),
    .A3(_12815_),
    .B1(_12814_),
    .B2(_12858_),
    .Y(_13905_));
 sky130_fd_sc_hd__nand3_1 _41205_ (.A(_13871_),
    .B(_13875_),
    .C(_13903_),
    .Y(_13906_));
 sky130_fd_sc_hd__nand3_1 _41206_ (.A(_13904_),
    .B(_13905_),
    .C(_13906_),
    .Y(_13907_));
 sky130_fd_sc_hd__nand3b_1 _41207_ (.A_N(_13903_),
    .B(_13871_),
    .C(_13875_),
    .Y(_13908_));
 sky130_fd_sc_hd__nand2_1 _41208_ (.A(_13871_),
    .B(_13875_),
    .Y(_13909_));
 sky130_fd_sc_hd__nand2_1 _41209_ (.A(_13909_),
    .B(_13903_),
    .Y(_13910_));
 sky130_fd_sc_hd__nand3b_2 _41210_ (.A_N(_13905_),
    .B(_13908_),
    .C(_13910_),
    .Y(_13912_));
 sky130_fd_sc_hd__a21o_1 _41211_ (.A1(_12840_),
    .A2(_12842_),
    .B1(_12843_),
    .X(_13913_));
 sky130_fd_sc_hd__a21o_1 _41212_ (.A1(_13907_),
    .A2(_13912_),
    .B1(_13913_),
    .X(_13914_));
 sky130_fd_sc_hd__nand3_1 _41213_ (.A(_13913_),
    .B(_13907_),
    .C(_13912_),
    .Y(_13915_));
 sky130_fd_sc_hd__a32o_1 _41214_ (.A1(_11698_),
    .A2(_12850_),
    .A3(_12852_),
    .B1(_12860_),
    .B2(_12864_),
    .X(_13916_));
 sky130_fd_sc_hd__a21o_1 _41215_ (.A1(_13914_),
    .A2(_13915_),
    .B1(_13916_),
    .X(_13917_));
 sky130_fd_sc_hd__nand3_1 _41216_ (.A(_13916_),
    .B(_13914_),
    .C(_13915_),
    .Y(_13918_));
 sky130_fd_sc_hd__nand2_2 _41217_ (.A(_13917_),
    .B(_13918_),
    .Y(_13919_));
 sky130_fd_sc_hd__nand3_1 _41218_ (.A(_11690_),
    .B(_11694_),
    .C(_12871_),
    .Y(_13920_));
 sky130_fd_sc_hd__a21o_1 _41219_ (.A1(_12868_),
    .A2(_12861_),
    .B1(_12869_),
    .X(_13921_));
 sky130_fd_sc_hd__a22oi_1 _41220_ (.A1(_12861_),
    .A2(_12866_),
    .B1(_13921_),
    .B2(_11685_),
    .Y(_13923_));
 sky130_fd_sc_hd__nand2_2 _41221_ (.A(_13920_),
    .B(_13923_),
    .Y(_13924_));
 sky130_fd_sc_hd__a41o_2 _41222_ (.A1(_10422_),
    .A2(_11690_),
    .A3(_11692_),
    .A4(_12871_),
    .B1(_13924_),
    .X(_13925_));
 sky130_fd_sc_hd__xnor2_4 _41223_ (.A(_13919_),
    .B(_13925_),
    .Y(_00014_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41224_ (.A(_02017_),
    .X(_13926_));
 sky130_fd_sc_hd__and3_1 _41225_ (.A(_13844_),
    .B(_09543_),
    .C(_13926_),
    .X(_13927_));
 sky130_fd_sc_hd__a21oi_2 _41226_ (.A1(_13844_),
    .A2(_13926_),
    .B1(_09543_),
    .Y(_13928_));
 sky130_fd_sc_hd__a32o_1 _41227_ (.A1(_12893_),
    .A2(_13098_),
    .A3(_13099_),
    .B1(_13197_),
    .B2(_13189_),
    .X(_13929_));
 sky130_fd_sc_hd__a32oi_4 _41228_ (.A1(_12989_),
    .A2(_12990_),
    .A3(_12991_),
    .B1(_12988_),
    .B2(_13026_),
    .Y(_13930_));
 sky130_fd_sc_hd__nand2_1 _41229_ (.A(_12985_),
    .B(_12990_),
    .Y(_13931_));
 sky130_fd_sc_hd__nand2_2 _41230_ (.A(_12936_),
    .B(_12949_),
    .Y(_13933_));
 sky130_fd_sc_hd__and3_1 _41231_ (.A(_11823_),
    .B(_11825_),
    .C(_12900_),
    .X(_13934_));
 sky130_fd_sc_hd__a31o_1 _41232_ (.A1(_10567_),
    .A2(_11824_),
    .A3(_11827_),
    .B1(_11826_),
    .X(_13935_));
 sky130_fd_sc_hd__a21oi_1 _41233_ (.A1(_07763_),
    .A2(net178),
    .B1(_10583_),
    .Y(_13936_));
 sky130_fd_sc_hd__o22ai_1 _41234_ (.A1(_10571_),
    .A2(_10572_),
    .B1(_10575_),
    .B2(_13936_),
    .Y(_13937_));
 sky130_fd_sc_hd__a2bb2oi_2 _41235_ (.A1_N(_10570_),
    .A2_N(_12898_),
    .B1(_13935_),
    .B2(_13937_),
    .Y(_13938_));
 sky130_fd_sc_hd__o22ai_2 _41236_ (.A1(_10568_),
    .A2(_13934_),
    .B1(_12906_),
    .B2(_13938_),
    .Y(_13939_));
 sky130_fd_sc_hd__nand2_1 _41237_ (.A(_13939_),
    .B(_12914_),
    .Y(_13940_));
 sky130_fd_sc_hd__clkbuf_2 _41238_ (.A(_13940_),
    .X(_13941_));
 sky130_fd_sc_hd__o22ai_4 _41239_ (.A1(_10557_),
    .A2(_11835_),
    .B1(_12913_),
    .B2(_11837_),
    .Y(_13942_));
 sky130_fd_sc_hd__o221ai_4 _41240_ (.A1(_10568_),
    .A2(_13934_),
    .B1(_12906_),
    .B2(_13938_),
    .C1(_13942_),
    .Y(_13944_));
 sky130_fd_sc_hd__clkbuf_2 _41241_ (.A(_13944_),
    .X(_13945_));
 sky130_fd_sc_hd__buf_2 _41242_ (.A(_12908_),
    .X(_13946_));
 sky130_fd_sc_hd__a31oi_4 _41243_ (.A1(_13942_),
    .A2(_13946_),
    .A3(_12918_),
    .B1(_11858_),
    .Y(_13947_));
 sky130_fd_sc_hd__a221oi_1 _41244_ (.A1(_12911_),
    .A2(_12914_),
    .B1(_13941_),
    .B2(_13945_),
    .C1(_13947_),
    .Y(_13948_));
 sky130_fd_sc_hd__a31o_1 _41245_ (.A1(_13942_),
    .A2(_13946_),
    .A3(_12918_),
    .B1(_12895_),
    .X(_13949_));
 sky130_fd_sc_hd__nand2_1 _41246_ (.A(_13944_),
    .B(_13940_),
    .Y(_13950_));
 sky130_fd_sc_hd__a21oi_2 _41247_ (.A1(_12944_),
    .A2(_13949_),
    .B1(_13950_),
    .Y(_13951_));
 sky130_fd_sc_hd__a21oi_4 _41248_ (.A1(_13946_),
    .A2(_12918_),
    .B1(_13942_),
    .Y(_13952_));
 sky130_fd_sc_hd__o211a_1 _41249_ (.A1(_12916_),
    .A2(_12917_),
    .B1(_13946_),
    .C1(_12918_),
    .X(_13953_));
 sky130_fd_sc_hd__nor2_1 _41250_ (.A(_13952_),
    .B(_13953_),
    .Y(_13955_));
 sky130_fd_sc_hd__a21oi_1 _41251_ (.A1(_11851_),
    .A2(_12895_),
    .B1(_12942_),
    .Y(_13956_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41252_ (.A(_11858_),
    .X(_13957_));
 sky130_fd_sc_hd__a21oi_1 _41253_ (.A1(_12944_),
    .A2(_12923_),
    .B1(_13957_),
    .Y(_13958_));
 sky130_fd_sc_hd__a21oi_1 _41254_ (.A1(_13955_),
    .A2(_13956_),
    .B1(_13958_),
    .Y(_13959_));
 sky130_fd_sc_hd__o21ai_1 _41255_ (.A1(_13948_),
    .A2(_13951_),
    .B1(_13959_),
    .Y(_13960_));
 sky130_fd_sc_hd__o21ai_1 _41256_ (.A1(_13957_),
    .A2(_13953_),
    .B1(_13950_),
    .Y(_13961_));
 sky130_fd_sc_hd__o211ai_4 _41257_ (.A1(_13952_),
    .A2(_13947_),
    .B1(_13941_),
    .C1(_13944_),
    .Y(_13962_));
 sky130_fd_sc_hd__o21ai_1 _41258_ (.A1(_13952_),
    .A2(_13953_),
    .B1(_12925_),
    .Y(_13963_));
 sky130_fd_sc_hd__nand2_1 _41259_ (.A(_12947_),
    .B(_13963_),
    .Y(_13964_));
 sky130_fd_sc_hd__o211ai_2 _41260_ (.A1(_13952_),
    .A2(_13961_),
    .B1(_13962_),
    .C1(_13964_),
    .Y(_13966_));
 sky130_fd_sc_hd__a21o_1 _41261_ (.A1(_13960_),
    .A2(_13966_),
    .B1(_11803_),
    .X(_13967_));
 sky130_fd_sc_hd__clkbuf_2 _41262_ (.A(_12896_),
    .X(_13968_));
 sky130_fd_sc_hd__clkbuf_2 _41263_ (.A(_12897_),
    .X(_13969_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41264_ (.A(_13960_),
    .X(_13970_));
 sky130_fd_sc_hd__clkbuf_2 _41265_ (.A(_13966_),
    .X(_13971_));
 sky130_fd_sc_hd__o211ai_2 _41266_ (.A1(_13968_),
    .A2(_13969_),
    .B1(_13970_),
    .C1(_13971_),
    .Y(_13972_));
 sky130_fd_sc_hd__nand3_2 _41267_ (.A(_13933_),
    .B(_13967_),
    .C(_13972_),
    .Y(_13973_));
 sky130_fd_sc_hd__clkbuf_2 _41268_ (.A(_11803_),
    .X(_13974_));
 sky130_fd_sc_hd__a21oi_1 _41269_ (.A1(_13970_),
    .A2(_13971_),
    .B1(_13974_),
    .Y(_13975_));
 sky130_fd_sc_hd__o211a_1 _41270_ (.A1(_13968_),
    .A2(_12962_),
    .B1(_13970_),
    .C1(_13971_),
    .X(_13977_));
 sky130_fd_sc_hd__and2b_1 _41271_ (.A_N(_12950_),
    .B(_12949_),
    .X(_13978_));
 sky130_fd_sc_hd__o21ai_2 _41272_ (.A1(_13975_),
    .A2(_13977_),
    .B1(_13978_),
    .Y(_13979_));
 sky130_fd_sc_hd__clkbuf_2 _41273_ (.A(_10545_),
    .X(_13980_));
 sky130_fd_sc_hd__o2bb2ai_4 _41274_ (.A1_N(_13973_),
    .A2_N(_13979_),
    .B1(_12956_),
    .B2(_13980_),
    .Y(_13981_));
 sky130_fd_sc_hd__buf_2 _41275_ (.A(_13969_),
    .X(_13982_));
 sky130_fd_sc_hd__nand4_1 _41276_ (.A(_13979_),
    .B(_10640_),
    .C(_13973_),
    .D(_13982_),
    .Y(_13983_));
 sky130_fd_sc_hd__o21ai_1 _41277_ (.A1(_12967_),
    .A2(_12968_),
    .B1(_12941_),
    .Y(_13984_));
 sky130_fd_sc_hd__nand2_2 _41278_ (.A(_12955_),
    .B(_13984_),
    .Y(_13985_));
 sky130_fd_sc_hd__a21oi_2 _41279_ (.A1(_13981_),
    .A2(_13983_),
    .B1(_13985_),
    .Y(_13986_));
 sky130_fd_sc_hd__nand2_1 _41280_ (.A(_13970_),
    .B(_13971_),
    .Y(_13988_));
 sky130_fd_sc_hd__o211ai_4 _41281_ (.A1(_13933_),
    .A2(_13988_),
    .B1(_10640_),
    .C1(_13969_),
    .Y(_13989_));
 sky130_fd_sc_hd__and3_1 _41282_ (.A(_13933_),
    .B(_13967_),
    .C(_13972_),
    .X(_13990_));
 sky130_fd_sc_hd__o211a_1 _41283_ (.A1(_13989_),
    .A2(_13990_),
    .B1(_13985_),
    .C1(_13981_),
    .X(_13991_));
 sky130_fd_sc_hd__o21ai_1 _41284_ (.A1(_12963_),
    .A2(_12960_),
    .B1(_12961_),
    .Y(_13992_));
 sky130_fd_sc_hd__o21ai_1 _41285_ (.A1(_12961_),
    .A2(_12963_),
    .B1(_13992_),
    .Y(_13993_));
 sky130_fd_sc_hd__buf_1 _41286_ (.A(_13993_),
    .X(_13994_));
 sky130_fd_sc_hd__o21ai_2 _41287_ (.A1(_13986_),
    .A2(_13991_),
    .B1(_13994_),
    .Y(_13995_));
 sky130_fd_sc_hd__a21o_1 _41288_ (.A1(_13981_),
    .A2(_13983_),
    .B1(_13985_),
    .X(_13996_));
 sky130_fd_sc_hd__o211ai_4 _41289_ (.A1(_13989_),
    .A2(_13990_),
    .B1(_13985_),
    .C1(_13981_),
    .Y(_13997_));
 sky130_fd_sc_hd__nand3b_2 _41290_ (.A_N(_13994_),
    .B(_13996_),
    .C(_13997_),
    .Y(_13999_));
 sky130_fd_sc_hd__nand3_2 _41291_ (.A(_13931_),
    .B(_13995_),
    .C(_13999_),
    .Y(_14000_));
 sky130_fd_sc_hd__o21bai_1 _41292_ (.A1(_13986_),
    .A2(_13991_),
    .B1_N(_13993_),
    .Y(_14001_));
 sky130_fd_sc_hd__a21boi_1 _41293_ (.A1(_12974_),
    .A2(_12980_),
    .B1_N(_12985_),
    .Y(_14002_));
 sky130_fd_sc_hd__nand3_1 _41294_ (.A(_13994_),
    .B(_13996_),
    .C(_13997_),
    .Y(_14003_));
 sky130_fd_sc_hd__nand3_1 _41295_ (.A(_14001_),
    .B(_14002_),
    .C(_14003_),
    .Y(_14004_));
 sky130_fd_sc_hd__clkbuf_2 _41296_ (.A(_14004_),
    .X(_14005_));
 sky130_fd_sc_hd__o2111ai_2 _41297_ (.A1(_11797_),
    .A2(_11793_),
    .B1(_11883_),
    .C1(_04789_),
    .D1(_12975_),
    .Y(_14006_));
 sky130_fd_sc_hd__clkbuf_2 _41298_ (.A(_12997_),
    .X(_14007_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41299_ (.A(_12997_),
    .X(_14008_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41300_ (.A(_10644_),
    .X(_14010_));
 sky130_fd_sc_hd__a32oi_1 _41301_ (.A1(_11905_),
    .A2(_10643_),
    .A3(_14008_),
    .B1(_14010_),
    .B2(_10500_),
    .Y(_14011_));
 sky130_fd_sc_hd__a41o_1 _41302_ (.A1(_11905_),
    .A2(_10643_),
    .A3(_10500_),
    .A4(_14007_),
    .B1(_14011_),
    .X(_14012_));
 sky130_fd_sc_hd__buf_1 _41303_ (.A(_10527_),
    .X(_14013_));
 sky130_fd_sc_hd__nor2_1 _41304_ (.A(_07863_),
    .B(_09153_),
    .Y(_14014_));
 sky130_fd_sc_hd__and2_1 _41305_ (.A(_06363_),
    .B(_07695_),
    .X(_14015_));
 sky130_fd_sc_hd__a211oi_1 _41306_ (.A1(_10526_),
    .A2(_09203_),
    .B1(_14014_),
    .C1(_14015_),
    .Y(_14016_));
 sky130_fd_sc_hd__o211a_1 _41307_ (.A1(_14014_),
    .A2(_14015_),
    .B1(_10526_),
    .C1(_09203_),
    .X(_14017_));
 sky130_fd_sc_hd__or4_1 _41308_ (.A(_07867_),
    .B(_14016_),
    .C(_07878_),
    .D(_14017_),
    .X(_14018_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41309_ (.A(_14018_),
    .X(_14019_));
 sky130_fd_sc_hd__o21ai_1 _41310_ (.A1(_14017_),
    .A2(_14016_),
    .B1(_13002_),
    .Y(_14021_));
 sky130_fd_sc_hd__a22oi_1 _41311_ (.A1(_14013_),
    .A2(_14008_),
    .B1(_14019_),
    .B2(_14021_),
    .Y(_14022_));
 sky130_fd_sc_hd__and4_1 _41312_ (.A(_14019_),
    .B(_14021_),
    .C(_14013_),
    .D(_12997_),
    .X(_14023_));
 sky130_fd_sc_hd__or2_1 _41313_ (.A(_14022_),
    .B(_14023_),
    .X(_14024_));
 sky130_fd_sc_hd__xnor2_1 _41314_ (.A(_14012_),
    .B(_14024_),
    .Y(_14025_));
 sky130_fd_sc_hd__nand3_1 _41315_ (.A(_12975_),
    .B(_14006_),
    .C(_14025_),
    .Y(_14026_));
 sky130_fd_sc_hd__a21o_1 _41316_ (.A1(_12975_),
    .A2(_14006_),
    .B1(_14025_),
    .X(_14027_));
 sky130_fd_sc_hd__nand2_1 _41317_ (.A(_14026_),
    .B(_14027_),
    .Y(_14028_));
 sky130_fd_sc_hd__or2b_1 _41318_ (.A(_13000_),
    .B_N(_13018_),
    .X(_14029_));
 sky130_fd_sc_hd__or2b_1 _41319_ (.A(_14028_),
    .B_N(_14029_),
    .X(_14030_));
 sky130_fd_sc_hd__inv_2 _41320_ (.A(_14030_),
    .Y(_14032_));
 sky130_fd_sc_hd__and3b_1 _41321_ (.A_N(_13000_),
    .B(_13018_),
    .C(_14028_),
    .X(_14033_));
 sky130_fd_sc_hd__o2bb2ai_1 _41322_ (.A1_N(_14000_),
    .A2_N(_14005_),
    .B1(_14032_),
    .B2(_14033_),
    .Y(_14034_));
 sky130_fd_sc_hd__nor2_1 _41323_ (.A(_14029_),
    .B(_14028_),
    .Y(_14035_));
 sky130_fd_sc_hd__and2_1 _41324_ (.A(_14029_),
    .B(_14028_),
    .X(_14036_));
 sky130_fd_sc_hd__o211ai_2 _41325_ (.A1(_14035_),
    .A2(_14036_),
    .B1(_14000_),
    .C1(_14005_),
    .Y(_14037_));
 sky130_fd_sc_hd__nand3b_4 _41326_ (.A_N(_13930_),
    .B(_14034_),
    .C(_14037_),
    .Y(_14038_));
 sky130_fd_sc_hd__o2bb2ai_1 _41327_ (.A1_N(_14000_),
    .A2_N(_14005_),
    .B1(_14035_),
    .B2(_14036_),
    .Y(_14039_));
 sky130_fd_sc_hd__o211ai_2 _41328_ (.A1(_14032_),
    .A2(_14033_),
    .B1(_14000_),
    .C1(_14005_),
    .Y(_14040_));
 sky130_fd_sc_hd__nand3_4 _41329_ (.A(_14039_),
    .B(_13930_),
    .C(_14040_),
    .Y(_14041_));
 sky130_fd_sc_hd__clkbuf_2 _41330_ (.A(_11919_),
    .X(_14043_));
 sky130_fd_sc_hd__a221o_1 _41331_ (.A1(_07691_),
    .A2(_11772_),
    .B1(_13007_),
    .B2(_13010_),
    .C1(_13004_),
    .X(_14044_));
 sky130_fd_sc_hd__o21ai_2 _41332_ (.A1(_13004_),
    .A2(_13011_),
    .B1(_07698_),
    .Y(_14045_));
 sky130_fd_sc_hd__a221oi_1 _41333_ (.A1(_14007_),
    .A2(_14043_),
    .B1(_14044_),
    .B2(_14045_),
    .C1(_13016_),
    .Y(_14046_));
 sky130_fd_sc_hd__and3b_1 _41334_ (.A_N(_13006_),
    .B(_14013_),
    .C(_12993_),
    .X(_14047_));
 sky130_fd_sc_hd__o211a_1 _41335_ (.A1(_13016_),
    .A2(_14047_),
    .B1(_14044_),
    .C1(_14045_),
    .X(_14048_));
 sky130_fd_sc_hd__or2_1 _41336_ (.A(_14046_),
    .B(_14048_),
    .X(_14049_));
 sky130_fd_sc_hd__a21oi_1 _41337_ (.A1(_13073_),
    .A2(_13076_),
    .B1(_14049_),
    .Y(_14050_));
 sky130_fd_sc_hd__and3_1 _41338_ (.A(_13073_),
    .B(_13076_),
    .C(_14049_),
    .X(_14051_));
 sky130_fd_sc_hd__or2_1 _41339_ (.A(_14050_),
    .B(_14051_),
    .X(_14052_));
 sky130_fd_sc_hd__nor3b_1 _41340_ (.A(_13078_),
    .B(_13081_),
    .C_N(_14052_),
    .Y(_14054_));
 sky130_fd_sc_hd__nor2_1 _41341_ (.A(_04646_),
    .B(_09148_),
    .Y(_14055_));
 sky130_fd_sc_hd__a31o_1 _41342_ (.A1(_04635_),
    .A2(_04636_),
    .A3(_11738_),
    .B1(_14055_),
    .X(_14056_));
 sky130_fd_sc_hd__xor2_1 _41343_ (.A(_11748_),
    .B(_14056_),
    .X(_14057_));
 sky130_fd_sc_hd__and3b_1 _41344_ (.A_N(_09125_),
    .B(_03349_),
    .C(_13050_),
    .X(_14058_));
 sky130_fd_sc_hd__xnor2_1 _41345_ (.A(_14057_),
    .B(_14058_),
    .Y(_14059_));
 sky130_fd_sc_hd__buf_1 _41346_ (.A(_11768_),
    .X(_14060_));
 sky130_fd_sc_hd__and2b_1 _41347_ (.A_N(_13041_),
    .B(_14060_),
    .X(_14061_));
 sky130_fd_sc_hd__o21ai_1 _41348_ (.A1(_14060_),
    .A2(_03314_),
    .B1(_11749_),
    .Y(_14062_));
 sky130_fd_sc_hd__a21oi_1 _41349_ (.A1(_14060_),
    .A2(_03314_),
    .B1(_14062_),
    .Y(_14063_));
 sky130_fd_sc_hd__or3b_1 _41350_ (.A(_03314_),
    .B(_07703_),
    .C_N(_13041_),
    .X(_14065_));
 sky130_fd_sc_hd__nand3_1 _41351_ (.A(_13044_),
    .B(_13045_),
    .C(_13043_),
    .Y(_14066_));
 sky130_fd_sc_hd__o211a_1 _41352_ (.A1(_14061_),
    .A2(_14063_),
    .B1(_14065_),
    .C1(_14066_),
    .X(_14067_));
 sky130_fd_sc_hd__a211o_1 _41353_ (.A1(_14066_),
    .A2(_14065_),
    .B1(_14063_),
    .C1(_14061_),
    .X(_14068_));
 sky130_fd_sc_hd__or2b_1 _41354_ (.A(_14067_),
    .B_N(_14068_),
    .X(_14069_));
 sky130_fd_sc_hd__xnor2_1 _41355_ (.A(_14059_),
    .B(_14069_),
    .Y(_14070_));
 sky130_fd_sc_hd__o21ba_1 _41356_ (.A1(_13078_),
    .A2(_13081_),
    .B1_N(_14052_),
    .X(_14071_));
 sky130_fd_sc_hd__nor3_2 _41357_ (.A(_14054_),
    .B(_14070_),
    .C(_14071_),
    .Y(_14072_));
 sky130_fd_sc_hd__o21a_1 _41358_ (.A1(_14071_),
    .A2(_14054_),
    .B1(_14070_),
    .X(_14073_));
 sky130_fd_sc_hd__o211ai_2 _41359_ (.A1(_14072_),
    .A2(_14073_),
    .B1(_13021_),
    .C1(_13024_),
    .Y(_14074_));
 sky130_fd_sc_hd__a211o_1 _41360_ (.A1(_13021_),
    .A2(_13024_),
    .B1(_14072_),
    .C1(_14073_),
    .X(_14076_));
 sky130_fd_sc_hd__a21o_1 _41361_ (.A1(_13066_),
    .A2(_13088_),
    .B1(_13085_),
    .X(_14077_));
 sky130_fd_sc_hd__and3_1 _41362_ (.A(_14074_),
    .B(_14076_),
    .C(_14077_),
    .X(_14078_));
 sky130_fd_sc_hd__a21oi_1 _41363_ (.A1(_14074_),
    .A2(_14076_),
    .B1(_14077_),
    .Y(_14079_));
 sky130_fd_sc_hd__nor2_2 _41364_ (.A(_14078_),
    .B(_14079_),
    .Y(_14080_));
 sky130_fd_sc_hd__a21o_1 _41365_ (.A1(_14038_),
    .A2(_14041_),
    .B1(_14080_),
    .X(_14081_));
 sky130_fd_sc_hd__nand3_4 _41366_ (.A(_14038_),
    .B(_14041_),
    .C(_14080_),
    .Y(_14082_));
 sky130_fd_sc_hd__a32o_2 _41367_ (.A1(_13033_),
    .A2(_13034_),
    .A3(_13035_),
    .B1(_13032_),
    .B2(_13096_),
    .X(_14083_));
 sky130_fd_sc_hd__a21oi_2 _41368_ (.A1(_14081_),
    .A2(_14082_),
    .B1(_14083_),
    .Y(_14084_));
 sky130_fd_sc_hd__a21oi_4 _41369_ (.A1(_14038_),
    .A2(_14041_),
    .B1(_14080_),
    .Y(_14085_));
 sky130_fd_sc_hd__nand2_2 _41370_ (.A(_14083_),
    .B(_14082_),
    .Y(_14087_));
 sky130_fd_sc_hd__nor2_1 _41371_ (.A(_14085_),
    .B(_14087_),
    .Y(_14088_));
 sky130_fd_sc_hd__o21a_1 _41372_ (.A1(_13149_),
    .A2(_13181_),
    .B1(_13180_),
    .X(_14089_));
 sky130_fd_sc_hd__and4_1 _41373_ (.A(_12014_),
    .B(_12037_),
    .C(_12036_),
    .D(_13112_),
    .X(_14090_));
 sky130_fd_sc_hd__a41oi_2 _41374_ (.A1(_13205_),
    .A2(_10747_),
    .A3(_12036_),
    .A4(_12038_),
    .B1(_14090_),
    .Y(_14091_));
 sky130_fd_sc_hd__and3_1 _41375_ (.A(_13123_),
    .B(_13127_),
    .C(_13128_),
    .X(_14092_));
 sky130_fd_sc_hd__a221oi_2 _41376_ (.A1(_09391_),
    .A2(_13104_),
    .B1(_13128_),
    .B2(_13124_),
    .C1(_13105_),
    .Y(_14093_));
 sky130_fd_sc_hd__a21o_1 _41377_ (.A1(_09391_),
    .A2(_13104_),
    .B1(_12013_),
    .X(_14094_));
 sky130_fd_sc_hd__o211a_1 _41378_ (.A1(_13105_),
    .A2(_13124_),
    .B1(_14094_),
    .C1(_13128_),
    .X(_14095_));
 sky130_fd_sc_hd__or4_1 _41379_ (.A(_13122_),
    .B(_14092_),
    .C(_14093_),
    .D(_14095_),
    .X(_14096_));
 sky130_fd_sc_hd__o22ai_2 _41380_ (.A1(_13122_),
    .A2(_14092_),
    .B1(_14093_),
    .B2(_14095_),
    .Y(_14098_));
 sky130_fd_sc_hd__and2_1 _41381_ (.A(_14096_),
    .B(_14098_),
    .X(_14099_));
 sky130_fd_sc_hd__xnor2_1 _41382_ (.A(_14091_),
    .B(_14099_),
    .Y(_14100_));
 sky130_fd_sc_hd__o211a_1 _41383_ (.A1(_13122_),
    .A2(_13129_),
    .B1(_13132_),
    .C1(_13143_),
    .X(_14101_));
 sky130_fd_sc_hd__or3_1 _41384_ (.A(_13136_),
    .B(_13156_),
    .C(net186),
    .X(_14102_));
 sky130_fd_sc_hd__o21ai_1 _41385_ (.A1(_13140_),
    .A2(_13156_),
    .B1(_14102_),
    .Y(_14103_));
 sky130_fd_sc_hd__o21ai_1 _41386_ (.A1(_13154_),
    .A2(_13155_),
    .B1(_13159_),
    .Y(_14104_));
 sky130_fd_sc_hd__and4bb_1 _41387_ (.A_N(_11977_),
    .B_N(net246),
    .C(_13135_),
    .D(_14104_),
    .X(_14105_));
 sky130_fd_sc_hd__a21oi_1 _41388_ (.A1(_13121_),
    .A2(_12011_),
    .B1(_13139_),
    .Y(_14106_));
 sky130_fd_sc_hd__and3_1 _41389_ (.A(_08010_),
    .B(_13139_),
    .C(_12011_),
    .X(_14107_));
 sky130_fd_sc_hd__nor2_1 _41390_ (.A(_14106_),
    .B(_14107_),
    .Y(_14109_));
 sky130_fd_sc_hd__xor2_1 _41391_ (.A(_12013_),
    .B(_14109_),
    .X(_14110_));
 sky130_fd_sc_hd__o21ai_1 _41392_ (.A1(_14103_),
    .A2(_14105_),
    .B1(_14110_),
    .Y(_14111_));
 sky130_fd_sc_hd__or3_1 _41393_ (.A(_14110_),
    .B(_14103_),
    .C(_14105_),
    .X(_14112_));
 sky130_fd_sc_hd__and2_1 _41394_ (.A(_14111_),
    .B(_14112_),
    .X(_14113_));
 sky130_fd_sc_hd__o21a_1 _41395_ (.A1(_13142_),
    .A2(_14101_),
    .B1(_14113_),
    .X(_14114_));
 sky130_fd_sc_hd__a211oi_1 _41396_ (.A1(_13133_),
    .A2(_13143_),
    .B1(_14113_),
    .C1(_13142_),
    .Y(_14115_));
 sky130_fd_sc_hd__nor2_1 _41397_ (.A(_14114_),
    .B(_14115_),
    .Y(_14116_));
 sky130_fd_sc_hd__nor2_1 _41398_ (.A(_14100_),
    .B(_14116_),
    .Y(_14117_));
 sky130_fd_sc_hd__and2_1 _41399_ (.A(_14100_),
    .B(_14116_),
    .X(_14118_));
 sky130_fd_sc_hd__nor2_1 _41400_ (.A(_14117_),
    .B(_14118_),
    .Y(_14120_));
 sky130_fd_sc_hd__and2_1 _41401_ (.A(_03338_),
    .B(_07946_),
    .X(_14121_));
 sky130_fd_sc_hd__nor2_1 _41402_ (.A(_10802_),
    .B(_07946_),
    .Y(_14122_));
 sky130_fd_sc_hd__o21a_1 _41403_ (.A1(_14121_),
    .A2(_14122_),
    .B1(_10687_),
    .X(_14123_));
 sky130_fd_sc_hd__or3_1 _41404_ (.A(_09139_),
    .B(_14121_),
    .C(_14122_),
    .X(_14124_));
 sky130_fd_sc_hd__or4b_1 _41405_ (.A(_03341_),
    .B(_14123_),
    .C(_10797_),
    .D_N(_14124_),
    .X(_14125_));
 sky130_fd_sc_hd__o21ai_1 _41406_ (.A1(_14121_),
    .A2(_14122_),
    .B1(_11738_),
    .Y(_14126_));
 sky130_fd_sc_hd__a2bb2o_1 _41407_ (.A1_N(_12026_),
    .A2_N(_03341_),
    .B1(_14126_),
    .B2(_14124_),
    .X(_14127_));
 sky130_fd_sc_hd__and3_1 _41408_ (.A(_14125_),
    .B(_14127_),
    .C(_13051_),
    .X(_14128_));
 sky130_fd_sc_hd__a21oi_1 _41409_ (.A1(_14125_),
    .A2(_14127_),
    .B1(_13060_),
    .Y(_14129_));
 sky130_fd_sc_hd__or2_1 _41410_ (.A(_14128_),
    .B(_14129_),
    .X(_14131_));
 sky130_fd_sc_hd__o311a_1 _41411_ (.A1(_11737_),
    .A2(_13052_),
    .A3(_13058_),
    .B1(_14131_),
    .C1(_13057_),
    .X(_14132_));
 sky130_fd_sc_hd__a21o_1 _41412_ (.A1(_13057_),
    .A2(_13059_),
    .B1(_14131_),
    .X(_14133_));
 sky130_fd_sc_hd__inv_2 _41413_ (.A(_14133_),
    .Y(_14134_));
 sky130_fd_sc_hd__or3_1 _41414_ (.A(_14132_),
    .B(_14134_),
    .C(_13162_),
    .X(_14135_));
 sky130_fd_sc_hd__o21ai_1 _41415_ (.A1(_14132_),
    .A2(_14134_),
    .B1(_13162_),
    .Y(_14136_));
 sky130_fd_sc_hd__o21ba_1 _41416_ (.A1(_13049_),
    .A2(_13062_),
    .B1_N(_13048_),
    .X(_14137_));
 sky130_fd_sc_hd__a21boi_1 _41417_ (.A1(_14135_),
    .A2(_14136_),
    .B1_N(_14137_),
    .Y(_14138_));
 sky130_fd_sc_hd__and3b_1 _41418_ (.A_N(_14137_),
    .B(_14135_),
    .C(_14136_),
    .X(_14139_));
 sky130_fd_sc_hd__a2111oi_1 _41419_ (.A1(_11981_),
    .A2(_13168_),
    .B1(_14138_),
    .C1(_14139_),
    .D1(_13167_),
    .Y(_14140_));
 sky130_fd_sc_hd__a21oi_1 _41420_ (.A1(_11981_),
    .A2(_13168_),
    .B1(_13167_),
    .Y(_14142_));
 sky130_fd_sc_hd__o21ba_1 _41421_ (.A1(_14138_),
    .A2(_14139_),
    .B1_N(_14142_),
    .X(_14143_));
 sky130_fd_sc_hd__nor2_1 _41422_ (.A(_14140_),
    .B(_14143_),
    .Y(_14144_));
 sky130_fd_sc_hd__nand2_1 _41423_ (.A(_13171_),
    .B(_13176_),
    .Y(_14145_));
 sky130_fd_sc_hd__xnor2_1 _41424_ (.A(_14144_),
    .B(_14145_),
    .Y(_14146_));
 sky130_fd_sc_hd__nor2_1 _41425_ (.A(_14120_),
    .B(_14146_),
    .Y(_14147_));
 sky130_fd_sc_hd__and2_1 _41426_ (.A(_14120_),
    .B(_14146_),
    .X(_14148_));
 sky130_fd_sc_hd__a211oi_4 _41427_ (.A1(_13091_),
    .A2(_13093_),
    .B1(_14147_),
    .C1(_14148_),
    .Y(_14149_));
 sky130_fd_sc_hd__o221a_2 _41428_ (.A1(_13037_),
    .A2(_13092_),
    .B1(_14147_),
    .B2(_14148_),
    .C1(_13091_),
    .X(_14150_));
 sky130_fd_sc_hd__nor3_2 _41429_ (.A(_14089_),
    .B(_14149_),
    .C(_14150_),
    .Y(_14151_));
 sky130_fd_sc_hd__o221a_1 _41430_ (.A1(_13181_),
    .A2(_13149_),
    .B1(_14150_),
    .B2(_14149_),
    .C1(_13180_),
    .X(_14153_));
 sky130_fd_sc_hd__nor2_2 _41431_ (.A(_14151_),
    .B(_14153_),
    .Y(_14154_));
 sky130_fd_sc_hd__inv_2 _41432_ (.A(_14154_),
    .Y(_14155_));
 sky130_fd_sc_hd__o21ai_2 _41433_ (.A1(_14084_),
    .A2(_14088_),
    .B1(_14155_),
    .Y(_14156_));
 sky130_fd_sc_hd__a21o_1 _41434_ (.A1(_14081_),
    .A2(_14082_),
    .B1(_14083_),
    .X(_14157_));
 sky130_fd_sc_hd__o211ai_4 _41435_ (.A1(_14085_),
    .A2(_14087_),
    .B1(_14154_),
    .C1(_14157_),
    .Y(_14158_));
 sky130_fd_sc_hd__nand3_1 _41436_ (.A(_13929_),
    .B(_14156_),
    .C(_14158_),
    .Y(_14159_));
 sky130_fd_sc_hd__o21ai_1 _41437_ (.A1(_14084_),
    .A2(_14088_),
    .B1(_14154_),
    .Y(_14160_));
 sky130_fd_sc_hd__a32oi_2 _41438_ (.A1(_12893_),
    .A2(_13098_),
    .A3(_13099_),
    .B1(_13197_),
    .B2(_13189_),
    .Y(_14161_));
 sky130_fd_sc_hd__o221ai_2 _41439_ (.A1(_14151_),
    .A2(_14153_),
    .B1(_14085_),
    .B2(_14087_),
    .C1(_14157_),
    .Y(_14162_));
 sky130_fd_sc_hd__nand3_2 _41440_ (.A(_14160_),
    .B(_14161_),
    .C(_14162_),
    .Y(_14164_));
 sky130_fd_sc_hd__o21ba_1 _41441_ (.A1(_13115_),
    .A2(_13111_),
    .B1_N(_13110_),
    .X(_14165_));
 sky130_fd_sc_hd__nor2_2 _41442_ (.A(_13209_),
    .B(_14165_),
    .Y(_14166_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41443_ (.A(_13205_),
    .X(_14167_));
 sky130_fd_sc_hd__and3b_1 _41444_ (.A_N(_14167_),
    .B(_14165_),
    .C(_09455_),
    .X(_14168_));
 sky130_fd_sc_hd__a21oi_1 _41445_ (.A1(_13118_),
    .A2(_13147_),
    .B1(_13146_),
    .Y(_14169_));
 sky130_fd_sc_hd__o21a_1 _41446_ (.A1(_14166_),
    .A2(_14168_),
    .B1(_14169_),
    .X(_14170_));
 sky130_fd_sc_hd__nor3_1 _41447_ (.A(_14169_),
    .B(_14166_),
    .C(_14168_),
    .Y(_14171_));
 sky130_fd_sc_hd__a2111o_2 _41448_ (.A1(_12008_),
    .A2(_12021_),
    .B1(_13209_),
    .C1(_14170_),
    .D1(_14171_),
    .X(_14172_));
 sky130_fd_sc_hd__o21bai_2 _41449_ (.A1(_14170_),
    .A2(_14171_),
    .B1_N(_13210_),
    .Y(_14173_));
 sky130_fd_sc_hd__o211a_1 _41450_ (.A1(_13213_),
    .A2(_13214_),
    .B1(_14172_),
    .C1(_14173_),
    .X(_14175_));
 sky130_fd_sc_hd__a211oi_1 _41451_ (.A1(_14172_),
    .A2(_14173_),
    .B1(_13213_),
    .C1(_13214_),
    .Y(_14176_));
 sky130_fd_sc_hd__or2_1 _41452_ (.A(_14175_),
    .B(_14176_),
    .X(_14177_));
 sky130_fd_sc_hd__o21a_1 _41453_ (.A1(_13101_),
    .A2(_13184_),
    .B1(_13186_),
    .X(_14178_));
 sky130_fd_sc_hd__xnor2_2 _41454_ (.A(_14177_),
    .B(_14178_),
    .Y(_14179_));
 sky130_fd_sc_hd__xor2_2 _41455_ (.A(_13220_),
    .B(_14179_),
    .X(_14180_));
 sky130_fd_sc_hd__a21o_1 _41456_ (.A1(_14159_),
    .A2(_14164_),
    .B1(_14180_),
    .X(_14181_));
 sky130_fd_sc_hd__nand3_2 _41457_ (.A(_14159_),
    .B(_14164_),
    .C(_14180_),
    .Y(_14182_));
 sky130_fd_sc_hd__a21o_1 _41458_ (.A1(_13227_),
    .A2(_13223_),
    .B1(_13199_),
    .X(_14183_));
 sky130_fd_sc_hd__a21oi_2 _41459_ (.A1(_14181_),
    .A2(_14182_),
    .B1(_14183_),
    .Y(_14184_));
 sky130_fd_sc_hd__and3_1 _41460_ (.A(_14183_),
    .B(_14181_),
    .C(_14182_),
    .X(_14186_));
 sky130_fd_sc_hd__a21oi_2 _41461_ (.A1(_13203_),
    .A2(_13221_),
    .B1(_13237_),
    .Y(_14187_));
 sky130_fd_sc_hd__o21ai_1 _41462_ (.A1(_14184_),
    .A2(_14186_),
    .B1(_14187_),
    .Y(_14188_));
 sky130_fd_sc_hd__a21oi_1 _41463_ (.A1(_13227_),
    .A2(_13223_),
    .B1(_13199_),
    .Y(_14189_));
 sky130_fd_sc_hd__nand2_1 _41464_ (.A(_14181_),
    .B(_14182_),
    .Y(_14190_));
 sky130_fd_sc_hd__a21oi_1 _41465_ (.A1(_14190_),
    .A2(_14189_),
    .B1(_14187_),
    .Y(_14191_));
 sky130_fd_sc_hd__o21ai_2 _41466_ (.A1(_14189_),
    .A2(_14190_),
    .B1(_14191_),
    .Y(_14192_));
 sky130_fd_sc_hd__o21ai_1 _41467_ (.A1(_11728_),
    .A2(_12091_),
    .B1(_13232_),
    .Y(_14193_));
 sky130_fd_sc_hd__and2_1 _41468_ (.A(_13241_),
    .B(_14193_),
    .X(_14194_));
 sky130_fd_sc_hd__a21boi_2 _41469_ (.A1(_14188_),
    .A2(_14192_),
    .B1_N(_14194_),
    .Y(_14195_));
 sky130_fd_sc_hd__clkbuf_2 _41470_ (.A(_14195_),
    .X(_14197_));
 sky130_fd_sc_hd__nand3b_1 _41471_ (.A_N(_14194_),
    .B(_14188_),
    .C(_14192_),
    .Y(_14198_));
 sky130_fd_sc_hd__clkbuf_2 _41472_ (.A(_14198_),
    .X(_14199_));
 sky130_fd_sc_hd__inv_2 _41473_ (.A(_14199_),
    .Y(_14200_));
 sky130_fd_sc_hd__buf_6 _41474_ (.A(_12892_),
    .X(_14201_));
 sky130_fd_sc_hd__o22ai_2 _41475_ (.A1(_14197_),
    .A2(_14200_),
    .B1(_13252_),
    .B2(_14201_),
    .Y(_14202_));
 sky130_fd_sc_hd__inv_2 _41476_ (.A(_13249_),
    .Y(_14203_));
 sky130_fd_sc_hd__a21o_1 _41477_ (.A1(_11588_),
    .A2(_12727_),
    .B1(_12723_),
    .X(_14204_));
 sky130_fd_sc_hd__o22ai_1 _41478_ (.A1(_13244_),
    .A2(_13254_),
    .B1(_13252_),
    .B2(_14201_),
    .Y(_14205_));
 sky130_fd_sc_hd__inv_2 _41479_ (.A(_14195_),
    .Y(_14206_));
 sky130_fd_sc_hd__nand2_1 _41480_ (.A(_14206_),
    .B(_14199_),
    .Y(_14208_));
 sky130_fd_sc_hd__inv_2 _41481_ (.A(_14208_),
    .Y(_14209_));
 sky130_fd_sc_hd__nand2_2 _41482_ (.A(_14205_),
    .B(_14209_),
    .Y(_14210_));
 sky130_fd_sc_hd__o211a_1 _41483_ (.A1(_14202_),
    .A2(_14203_),
    .B1(_14204_),
    .C1(_14210_),
    .X(_14211_));
 sky130_fd_sc_hd__o221ai_2 _41484_ (.A1(_14197_),
    .A2(_14200_),
    .B1(_13252_),
    .B2(_14201_),
    .C1(_13249_),
    .Y(_14212_));
 sky130_fd_sc_hd__a21oi_1 _41485_ (.A1(_14210_),
    .A2(_14212_),
    .B1(_14204_),
    .Y(_14213_));
 sky130_fd_sc_hd__o21ai_1 _41486_ (.A1(_14211_),
    .A2(_14213_),
    .B1(_12127_),
    .Y(_14214_));
 sky130_fd_sc_hd__clkbuf_2 _41487_ (.A(_13800_),
    .X(_14215_));
 sky130_fd_sc_hd__o221ai_4 _41488_ (.A1(_13270_),
    .A2(_14215_),
    .B1(_14203_),
    .B2(_14202_),
    .C1(_14210_),
    .Y(_14216_));
 sky130_fd_sc_hd__a21o_1 _41489_ (.A1(_14210_),
    .A2(_14212_),
    .B1(_14204_),
    .X(_14217_));
 sky130_fd_sc_hd__nand3_1 _41490_ (.A(_10935_),
    .B(_14216_),
    .C(_14217_),
    .Y(_14219_));
 sky130_fd_sc_hd__nor2_1 _41491_ (.A(_13798_),
    .B(_13804_),
    .Y(_14220_));
 sky130_fd_sc_hd__nand3_1 _41492_ (.A(_14214_),
    .B(_14219_),
    .C(_14220_),
    .Y(_14221_));
 sky130_fd_sc_hd__clkbuf_2 _41493_ (.A(_14221_),
    .X(_14222_));
 sky130_fd_sc_hd__nand3_1 _41494_ (.A(_14217_),
    .B(_12127_),
    .C(_14216_),
    .Y(_14223_));
 sky130_fd_sc_hd__o21bai_1 _41495_ (.A1(_14211_),
    .A2(_14213_),
    .B1_N(_12127_),
    .Y(_14224_));
 sky130_fd_sc_hd__o211ai_2 _41496_ (.A1(_13798_),
    .A2(_13804_),
    .B1(_14223_),
    .C1(_14224_),
    .Y(_14225_));
 sky130_fd_sc_hd__buf_1 _41497_ (.A(_14225_),
    .X(_14226_));
 sky130_fd_sc_hd__nand2_1 _41498_ (.A(_14222_),
    .B(_14226_),
    .Y(_14227_));
 sky130_fd_sc_hd__a21oi_2 _41499_ (.A1(_13272_),
    .A2(_12880_),
    .B1(_13266_),
    .Y(_14228_));
 sky130_fd_sc_hd__nand2_1 _41500_ (.A(_14227_),
    .B(_14228_),
    .Y(_14230_));
 sky130_fd_sc_hd__nor2_1 _41501_ (.A(_12885_),
    .B(_13268_),
    .Y(_14231_));
 sky130_fd_sc_hd__o211ai_1 _41502_ (.A1(_13266_),
    .A2(_14231_),
    .B1(_14222_),
    .C1(_14226_),
    .Y(_14232_));
 sky130_fd_sc_hd__inv_2 _41503_ (.A(_13280_),
    .Y(_14233_));
 sky130_fd_sc_hd__a21o_1 _41504_ (.A1(_13283_),
    .A2(_13277_),
    .B1(_14233_),
    .X(_14234_));
 sky130_fd_sc_hd__a21oi_1 _41505_ (.A1(_14230_),
    .A2(_14232_),
    .B1(_14234_),
    .Y(_14235_));
 sky130_fd_sc_hd__o211a_2 _41506_ (.A1(_13266_),
    .A2(_14231_),
    .B1(_14221_),
    .C1(_14225_),
    .X(_14236_));
 sky130_fd_sc_hd__a221oi_4 _41507_ (.A1(_13281_),
    .A2(_13282_),
    .B1(_14227_),
    .B2(_14228_),
    .C1(_14236_),
    .Y(_14237_));
 sky130_fd_sc_hd__o22ai_2 _41508_ (.A1(_13927_),
    .A2(_13928_),
    .B1(_14235_),
    .B2(_14237_),
    .Y(_14238_));
 sky130_fd_sc_hd__o21ai_1 _41509_ (.A1(_14233_),
    .A2(_13288_),
    .B1(_14230_),
    .Y(_14239_));
 sky130_fd_sc_hd__nor2_1 _41510_ (.A(_13927_),
    .B(_13928_),
    .Y(_14241_));
 sky130_fd_sc_hd__inv_2 _41511_ (.A(_14228_),
    .Y(_14242_));
 sky130_fd_sc_hd__a21oi_1 _41512_ (.A1(_14222_),
    .A2(_14226_),
    .B1(_14242_),
    .Y(_14243_));
 sky130_fd_sc_hd__o21bai_1 _41513_ (.A1(_14243_),
    .A2(_14236_),
    .B1_N(_14234_),
    .Y(_14244_));
 sky130_fd_sc_hd__o211ai_2 _41514_ (.A1(_14236_),
    .A2(_14239_),
    .B1(_14241_),
    .C1(_14244_),
    .Y(_14245_));
 sky130_fd_sc_hd__a21o_1 _41515_ (.A1(_13810_),
    .A2(_13714_),
    .B1(_13808_),
    .X(_14246_));
 sky130_fd_sc_hd__a21oi_2 _41516_ (.A1(_14238_),
    .A2(_14245_),
    .B1(_14246_),
    .Y(_14247_));
 sky130_fd_sc_hd__buf_1 _41517_ (.A(_14244_),
    .X(_14248_));
 sky130_fd_sc_hd__nand2_1 _41518_ (.A(_14248_),
    .B(_14241_),
    .Y(_14249_));
 sky130_fd_sc_hd__o221a_1 _41519_ (.A1(_13808_),
    .A2(_13813_),
    .B1(_14237_),
    .B2(_14249_),
    .C1(_14238_),
    .X(_14250_));
 sky130_fd_sc_hd__o21ai_1 _41520_ (.A1(_12879_),
    .A2(_12883_),
    .B1(_13290_),
    .Y(_14252_));
 sky130_fd_sc_hd__and2_1 _41521_ (.A(_13287_),
    .B(_14252_),
    .X(_14253_));
 sky130_fd_sc_hd__o21ai_1 _41522_ (.A1(_14247_),
    .A2(_14250_),
    .B1(_14253_),
    .Y(_14254_));
 sky130_fd_sc_hd__clkbuf_2 _41523_ (.A(_14254_),
    .X(_14255_));
 sky130_fd_sc_hd__nand2_1 _41524_ (.A(_13287_),
    .B(_14252_),
    .Y(_14256_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41525_ (.A(_02015_),
    .X(_14257_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41526_ (.A(_00395_),
    .X(_14258_));
 sky130_fd_sc_hd__clkbuf_2 _41527_ (.A(_03565_),
    .X(_14259_));
 sky130_fd_sc_hd__xnor2_1 _41528_ (.A(_14259_),
    .B(_12881_),
    .Y(_14260_));
 sky130_fd_sc_hd__or3_1 _41529_ (.A(_14257_),
    .B(_14258_),
    .C(_14260_),
    .X(_14261_));
 sky130_fd_sc_hd__o21ai_1 _41530_ (.A1(_14257_),
    .A2(_14258_),
    .B1(_14260_),
    .Y(_14263_));
 sky130_fd_sc_hd__o211ai_1 _41531_ (.A1(_14233_),
    .A2(_13288_),
    .B1(_14230_),
    .C1(_14232_),
    .Y(_14264_));
 sky130_fd_sc_hd__a22oi_1 _41532_ (.A1(_14261_),
    .A2(_14263_),
    .B1(_14248_),
    .B2(_14264_),
    .Y(_14265_));
 sky130_fd_sc_hd__o211a_1 _41533_ (.A1(_14236_),
    .A2(_14239_),
    .B1(_14241_),
    .C1(_14248_),
    .X(_14266_));
 sky130_fd_sc_hd__o21bai_1 _41534_ (.A1(_14265_),
    .A2(_14266_),
    .B1_N(_14246_),
    .Y(_14267_));
 sky130_fd_sc_hd__nand3_2 _41535_ (.A(_14246_),
    .B(_14238_),
    .C(_14245_),
    .Y(_14268_));
 sky130_fd_sc_hd__nand3_1 _41536_ (.A(_14256_),
    .B(_14267_),
    .C(_14268_),
    .Y(_14269_));
 sky130_fd_sc_hd__clkbuf_2 _41537_ (.A(_14269_),
    .X(_14270_));
 sky130_fd_sc_hd__a211o_1 _41538_ (.A1(_12495_),
    .A2(_12385_),
    .B1(_13703_),
    .C1(net73),
    .X(_14271_));
 sky130_fd_sc_hd__o31ai_2 _41539_ (.A1(_13423_),
    .A2(_13424_),
    .A3(_13706_),
    .B1(_14271_),
    .Y(_14272_));
 sky130_fd_sc_hd__o21bai_2 _41540_ (.A1(_13508_),
    .A2(_13484_),
    .B1_N(_13507_),
    .Y(_14274_));
 sky130_fd_sc_hd__nand3_1 _41541_ (.A(_08417_),
    .B(_13490_),
    .C(_12391_),
    .Y(_14275_));
 sky130_fd_sc_hd__o21ai_1 _41542_ (.A1(_13490_),
    .A2(_11209_),
    .B1(_14275_),
    .Y(_14276_));
 sky130_fd_sc_hd__o21ai_1 _41543_ (.A1(_11206_),
    .A2(_13488_),
    .B1(_13495_),
    .Y(_14277_));
 sky130_fd_sc_hd__xnor2_1 _41544_ (.A(_14276_),
    .B(_14277_),
    .Y(_14278_));
 sky130_fd_sc_hd__a21oi_1 _41545_ (.A1(_13497_),
    .A2(_13498_),
    .B1(_14278_),
    .Y(_14279_));
 sky130_fd_sc_hd__and3_1 _41546_ (.A(_13497_),
    .B(_13498_),
    .C(_14278_),
    .X(_14280_));
 sky130_fd_sc_hd__nor3_1 _41547_ (.A(_14279_),
    .B(_12393_),
    .C(_14280_),
    .Y(_14281_));
 sky130_fd_sc_hd__o21ai_1 _41548_ (.A1(_14280_),
    .A2(_14279_),
    .B1(_12393_),
    .Y(_14282_));
 sky130_fd_sc_hd__and2b_1 _41549_ (.A_N(_14281_),
    .B(_14282_),
    .X(_14283_));
 sky130_fd_sc_hd__and2_1 _41550_ (.A(_14283_),
    .B(_13503_),
    .X(_14285_));
 sky130_fd_sc_hd__nor2_1 _41551_ (.A(_13503_),
    .B(_14283_),
    .Y(_14286_));
 sky130_fd_sc_hd__nor2_1 _41552_ (.A(_14285_),
    .B(_14286_),
    .Y(_14287_));
 sky130_fd_sc_hd__xor2_1 _41553_ (.A(_14274_),
    .B(_14287_),
    .X(_14288_));
 sky130_fd_sc_hd__a21boi_1 _41554_ (.A1(_12423_),
    .A2(_13437_),
    .B1_N(_13440_),
    .Y(_14289_));
 sky130_fd_sc_hd__clkbuf_2 _41555_ (.A(_12432_),
    .X(_14290_));
 sky130_fd_sc_hd__o21a_1 _41556_ (.A1(_13428_),
    .A2(_12425_),
    .B1(_13426_),
    .X(_14291_));
 sky130_fd_sc_hd__a21oi_1 _41557_ (.A1(_12419_),
    .A2(_13428_),
    .B1(_14291_),
    .Y(_14292_));
 sky130_fd_sc_hd__a21oi_2 _41558_ (.A1(_12419_),
    .A2(_14291_),
    .B1(_14292_),
    .Y(_14293_));
 sky130_fd_sc_hd__buf_1 _41559_ (.A(_12425_),
    .X(_14294_));
 sky130_fd_sc_hd__buf_1 _41560_ (.A(_13428_),
    .X(_14296_));
 sky130_fd_sc_hd__a211oi_1 _41561_ (.A1(_13426_),
    .A2(_14294_),
    .B1(_14296_),
    .C1(_12419_),
    .Y(_14297_));
 sky130_fd_sc_hd__o221ai_2 _41562_ (.A1(_14290_),
    .A2(_11277_),
    .B1(_14293_),
    .B2(_14297_),
    .C1(_13434_),
    .Y(_14298_));
 sky130_fd_sc_hd__or4_1 _41563_ (.A(_12421_),
    .B(_14290_),
    .C(_11274_),
    .D(_11275_),
    .X(_14299_));
 sky130_fd_sc_hd__a211oi_1 _41564_ (.A1(_14299_),
    .A2(_13434_),
    .B1(_14293_),
    .C1(_14297_),
    .Y(_14300_));
 sky130_fd_sc_hd__a31o_1 _41565_ (.A1(_11269_),
    .A2(_12428_),
    .A3(_14298_),
    .B1(_14300_),
    .X(_14301_));
 sky130_fd_sc_hd__o21bai_1 _41566_ (.A1(_13433_),
    .A2(_14298_),
    .B1_N(_14301_),
    .Y(_14302_));
 sky130_fd_sc_hd__and2_1 _41567_ (.A(_14289_),
    .B(_14302_),
    .X(_14303_));
 sky130_fd_sc_hd__nor2_1 _41568_ (.A(_14302_),
    .B(_14289_),
    .Y(_14304_));
 sky130_fd_sc_hd__nor2_1 _41569_ (.A(_14303_),
    .B(_14304_),
    .Y(_14305_));
 sky130_fd_sc_hd__a21boi_2 _41570_ (.A1(_13444_),
    .A2(_13448_),
    .B1_N(_14305_),
    .Y(_14307_));
 sky130_fd_sc_hd__o211a_1 _41571_ (.A1(_14303_),
    .A2(_14304_),
    .B1(_13444_),
    .C1(_13448_),
    .X(_14308_));
 sky130_fd_sc_hd__o31ai_1 _41572_ (.A1(_11233_),
    .A2(_12470_),
    .A3(_13472_),
    .B1(_13473_),
    .Y(_14309_));
 sky130_fd_sc_hd__clkbuf_2 _41573_ (.A(_13465_),
    .X(_14310_));
 sky130_fd_sc_hd__nand2_1 _41574_ (.A(_08456_),
    .B(_13458_),
    .Y(_14311_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41575_ (.A(_10038_),
    .X(_14312_));
 sky130_fd_sc_hd__buf_1 _41576_ (.A(_11236_),
    .X(_14313_));
 sky130_fd_sc_hd__nand2_1 _41577_ (.A(_13455_),
    .B(_14313_),
    .Y(_14314_));
 sky130_fd_sc_hd__o22ai_1 _41578_ (.A1(_14314_),
    .A2(_13465_),
    .B1(_14313_),
    .B2(_13454_),
    .Y(_14315_));
 sky130_fd_sc_hd__buf_1 _41579_ (.A(_14315_),
    .X(_14316_));
 sky130_fd_sc_hd__a21bo_1 _41580_ (.A1(_14311_),
    .A2(_14312_),
    .B1_N(_14316_),
    .X(_14318_));
 sky130_fd_sc_hd__clkbuf_2 _41581_ (.A(_08456_),
    .X(_14319_));
 sky130_fd_sc_hd__a211o_1 _41582_ (.A1(_14319_),
    .A2(_13458_),
    .B1(_14315_),
    .C1(_10045_),
    .X(_14320_));
 sky130_fd_sc_hd__and4_1 _41583_ (.A(_13457_),
    .B(_14318_),
    .C(_14320_),
    .D(_13465_),
    .X(_14321_));
 sky130_fd_sc_hd__a22oi_2 _41584_ (.A1(_14310_),
    .A2(_13457_),
    .B1(_14318_),
    .B2(_14320_),
    .Y(_14322_));
 sky130_fd_sc_hd__o2111ai_2 _41585_ (.A1(_11233_),
    .A2(_14310_),
    .B1(_13464_),
    .C1(_13463_),
    .D1(_13462_),
    .Y(_14323_));
 sky130_fd_sc_hd__o211ai_2 _41586_ (.A1(_14321_),
    .A2(_14322_),
    .B1(_13462_),
    .C1(_14323_),
    .Y(_14324_));
 sky130_fd_sc_hd__a211o_1 _41587_ (.A1(_13462_),
    .A2(_14323_),
    .B1(_14321_),
    .C1(_14322_),
    .X(_14325_));
 sky130_fd_sc_hd__o311a_1 _41588_ (.A1(_11233_),
    .A2(_14310_),
    .A3(_12469_),
    .B1(_14324_),
    .C1(_14325_),
    .X(_14326_));
 sky130_fd_sc_hd__a21oi_1 _41589_ (.A1(_14325_),
    .A2(_14324_),
    .B1(_13466_),
    .Y(_14327_));
 sky130_fd_sc_hd__or2_1 _41590_ (.A(_14326_),
    .B(_14327_),
    .X(_14329_));
 sky130_fd_sc_hd__nor2_1 _41591_ (.A(_14309_),
    .B(_14329_),
    .Y(_14330_));
 sky130_fd_sc_hd__and2_1 _41592_ (.A(_14309_),
    .B(_14329_),
    .X(_14331_));
 sky130_fd_sc_hd__or2_1 _41593_ (.A(_14330_),
    .B(_14331_),
    .X(_14332_));
 sky130_fd_sc_hd__a21boi_1 _41594_ (.A1(_13452_),
    .A2(_13478_),
    .B1_N(_13477_),
    .Y(_14333_));
 sky130_fd_sc_hd__xor2_1 _41595_ (.A(_14332_),
    .B(_14333_),
    .X(_14334_));
 sky130_fd_sc_hd__or2b_1 _41596_ (.A(_14308_),
    .B_N(_14334_),
    .X(_14335_));
 sky130_fd_sc_hd__o21bai_1 _41597_ (.A1(_14307_),
    .A2(_14308_),
    .B1_N(_14334_),
    .Y(_14336_));
 sky130_fd_sc_hd__o21a_1 _41598_ (.A1(_14307_),
    .A2(_14335_),
    .B1(_14336_),
    .X(_14337_));
 sky130_fd_sc_hd__or2_1 _41599_ (.A(_14288_),
    .B(_14337_),
    .X(_14338_));
 sky130_fd_sc_hd__nand2_1 _41600_ (.A(_14288_),
    .B(_14337_),
    .Y(_14340_));
 sky130_fd_sc_hd__a2bb2o_4 _41601_ (.A1_N(_13662_),
    .A2_N(_13697_),
    .B1(_13628_),
    .B2(_13661_),
    .X(_14341_));
 sky130_fd_sc_hd__a21oi_1 _41602_ (.A1(_14338_),
    .A2(_14340_),
    .B1(_14341_),
    .Y(_14342_));
 sky130_fd_sc_hd__nand3_1 _41603_ (.A(_14341_),
    .B(_14338_),
    .C(_14340_),
    .Y(_14343_));
 sky130_fd_sc_hd__or2b_1 _41604_ (.A(_14342_),
    .B_N(_14343_),
    .X(_14344_));
 sky130_fd_sc_hd__and2_1 _41605_ (.A(_13448_),
    .B(_13450_),
    .X(_14345_));
 sky130_fd_sc_hd__a21oi_2 _41606_ (.A1(_14345_),
    .A2(_13480_),
    .B1(_13511_),
    .Y(_14346_));
 sky130_fd_sc_hd__nand2_1 _41607_ (.A(_14344_),
    .B(_14346_),
    .Y(_14347_));
 sky130_fd_sc_hd__or2_1 _41608_ (.A(_14346_),
    .B(_14344_),
    .X(_14348_));
 sky130_fd_sc_hd__and2_1 _41609_ (.A(_14347_),
    .B(_14348_),
    .X(_14349_));
 sky130_fd_sc_hd__o21a_1 _41610_ (.A1(_13597_),
    .A2(_13698_),
    .B1(_13598_),
    .X(_14351_));
 sky130_fd_sc_hd__and3_1 _41611_ (.A(_13524_),
    .B(_13519_),
    .C(_09924_),
    .X(_14352_));
 sky130_fd_sc_hd__buf_1 _41612_ (.A(_09924_),
    .X(_14353_));
 sky130_fd_sc_hd__nor2_1 _41613_ (.A(_14353_),
    .B(_13519_),
    .Y(_14354_));
 sky130_fd_sc_hd__o22ai_1 _41614_ (.A1(_08598_),
    .A2(_12329_),
    .B1(_14352_),
    .B2(_14354_),
    .Y(_14355_));
 sky130_fd_sc_hd__or4_1 _41615_ (.A(_08598_),
    .B(_14354_),
    .C(_12329_),
    .D(_14352_),
    .X(_14356_));
 sky130_fd_sc_hd__or4bb_1 _41616_ (.A(_13527_),
    .B(_13529_),
    .C_N(_14355_),
    .D_N(_14356_),
    .X(_14357_));
 sky130_fd_sc_hd__a2bb2o_1 _41617_ (.A1_N(_13527_),
    .A2_N(net175),
    .B1(_14355_),
    .B2(_14356_),
    .X(_14358_));
 sky130_fd_sc_hd__and3_1 _41618_ (.A(_14357_),
    .B(_14358_),
    .C(_13530_),
    .X(_14359_));
 sky130_fd_sc_hd__a21oi_2 _41619_ (.A1(_14357_),
    .A2(_14358_),
    .B1(_13530_),
    .Y(_14360_));
 sky130_fd_sc_hd__o21a_1 _41620_ (.A1(_14359_),
    .A2(_14360_),
    .B1(_13535_),
    .X(_14362_));
 sky130_fd_sc_hd__inv_2 _41621_ (.A(_14362_),
    .Y(_14363_));
 sky130_fd_sc_hd__a21o_1 _41622_ (.A1(_12337_),
    .A2(_13538_),
    .B1(_13536_),
    .X(_14364_));
 sky130_fd_sc_hd__o311ai_4 _41623_ (.A1(_13535_),
    .A2(_14359_),
    .A3(_14360_),
    .B1(_14364_),
    .C1(_13563_),
    .Y(_14365_));
 sky130_fd_sc_hd__and3_1 _41624_ (.A(_14364_),
    .B(_13563_),
    .C(_14362_),
    .X(_14366_));
 sky130_fd_sc_hd__a21o_1 _41625_ (.A1(_14363_),
    .A2(_14365_),
    .B1(_14366_),
    .X(_14367_));
 sky130_fd_sc_hd__clkbuf_2 _41626_ (.A(_11168_),
    .X(_14368_));
 sky130_fd_sc_hd__clkbuf_2 _41627_ (.A(_13543_),
    .X(_14369_));
 sky130_fd_sc_hd__and3b_1 _41628_ (.A_N(_13545_),
    .B(_13543_),
    .C(_13552_),
    .X(_14370_));
 sky130_fd_sc_hd__nor3_1 _41629_ (.A(_14368_),
    .B(_13549_),
    .C(_14370_),
    .Y(_14371_));
 sky130_fd_sc_hd__o21a_1 _41630_ (.A1(_13549_),
    .A2(_14370_),
    .B1(_14368_),
    .X(_14373_));
 sky130_fd_sc_hd__o21ba_1 _41631_ (.A1(_14371_),
    .A2(_14373_),
    .B1_N(_13546_),
    .X(_14374_));
 sky130_fd_sc_hd__a41o_1 _41632_ (.A1(_11158_),
    .A2(_14368_),
    .A3(_13545_),
    .A4(_14369_),
    .B1(_14374_),
    .X(_14375_));
 sky130_fd_sc_hd__o21ba_1 _41633_ (.A1(_12355_),
    .A2(_13554_),
    .B1_N(_13551_),
    .X(_14376_));
 sky130_fd_sc_hd__or2_1 _41634_ (.A(_14375_),
    .B(_14376_),
    .X(_14377_));
 sky130_fd_sc_hd__nand2_1 _41635_ (.A(_14376_),
    .B(_14375_),
    .Y(_14378_));
 sky130_fd_sc_hd__o211a_1 _41636_ (.A1(_13556_),
    .A2(_13560_),
    .B1(_14377_),
    .C1(_14378_),
    .X(_14379_));
 sky130_fd_sc_hd__a211oi_1 _41637_ (.A1(_14377_),
    .A2(_14378_),
    .B1(_13556_),
    .C1(_13560_),
    .Y(_14380_));
 sky130_fd_sc_hd__or2_1 _41638_ (.A(_14379_),
    .B(_14380_),
    .X(_14381_));
 sky130_fd_sc_hd__nand2_1 _41639_ (.A(_14367_),
    .B(_14381_),
    .Y(_14382_));
 sky130_fd_sc_hd__a211o_1 _41640_ (.A1(_14363_),
    .A2(_14365_),
    .B1(_14366_),
    .C1(_14381_),
    .X(_14384_));
 sky130_fd_sc_hd__a21oi_2 _41641_ (.A1(_13591_),
    .A2(_13589_),
    .B1(_13586_),
    .Y(_14385_));
 sky130_fd_sc_hd__clkbuf_2 _41642_ (.A(_12311_),
    .X(_14386_));
 sky130_fd_sc_hd__buf_1 _41643_ (.A(_09969_),
    .X(_14387_));
 sky130_fd_sc_hd__o21a_1 _41644_ (.A1(_13568_),
    .A2(_11110_),
    .B1(_13567_),
    .X(_14388_));
 sky130_fd_sc_hd__a21oi_1 _41645_ (.A1(_09969_),
    .A2(_13568_),
    .B1(_14388_),
    .Y(_14389_));
 sky130_fd_sc_hd__a21oi_1 _41646_ (.A1(_14387_),
    .A2(_14388_),
    .B1(_14389_),
    .Y(_14390_));
 sky130_fd_sc_hd__buf_1 _41647_ (.A(_11110_),
    .X(_14391_));
 sky130_fd_sc_hd__buf_1 _41648_ (.A(_13568_),
    .X(_14392_));
 sky130_fd_sc_hd__a211oi_1 _41649_ (.A1(_13567_),
    .A2(_14391_),
    .B1(_14392_),
    .C1(_14387_),
    .Y(_14393_));
 sky130_fd_sc_hd__o221ai_2 _41650_ (.A1(_14386_),
    .A2(_11102_),
    .B1(_14390_),
    .B2(_14393_),
    .C1(_13576_),
    .Y(_14395_));
 sky130_fd_sc_hd__or4_1 _41651_ (.A(_13573_),
    .B(_12311_),
    .C(_11099_),
    .D(_11100_),
    .X(_14396_));
 sky130_fd_sc_hd__a211oi_1 _41652_ (.A1(_14396_),
    .A2(_13576_),
    .B1(_14390_),
    .C1(_14393_),
    .Y(_14397_));
 sky130_fd_sc_hd__a31o_1 _41653_ (.A1(_09971_),
    .A2(_12307_),
    .A3(_14395_),
    .B1(_14397_),
    .X(_14398_));
 sky130_fd_sc_hd__o21bai_1 _41654_ (.A1(_13575_),
    .A2(_14395_),
    .B1_N(_14398_),
    .Y(_14399_));
 sky130_fd_sc_hd__o41a_1 _41655_ (.A1(_05739_),
    .A2(_07210_),
    .A3(_09962_),
    .A4(_13584_),
    .B1(_13583_),
    .X(_14400_));
 sky130_fd_sc_hd__or2_1 _41656_ (.A(_14399_),
    .B(_14400_),
    .X(_14401_));
 sky130_fd_sc_hd__nand2_1 _41657_ (.A(_14400_),
    .B(_14399_),
    .Y(_14402_));
 sky130_fd_sc_hd__nand2_2 _41658_ (.A(_14401_),
    .B(_14402_),
    .Y(_14403_));
 sky130_fd_sc_hd__xnor2_2 _41659_ (.A(_14385_),
    .B(_14403_),
    .Y(_14404_));
 sky130_fd_sc_hd__nand3_1 _41660_ (.A(_14382_),
    .B(_14384_),
    .C(_14404_),
    .Y(_14406_));
 sky130_fd_sc_hd__a21o_1 _41661_ (.A1(_14382_),
    .A2(_14384_),
    .B1(_14404_),
    .X(_14407_));
 sky130_fd_sc_hd__and2_1 _41662_ (.A(_13564_),
    .B(_13595_),
    .X(_14408_));
 sky130_fd_sc_hd__a21oi_4 _41663_ (.A1(_14406_),
    .A2(_14407_),
    .B1(_14408_),
    .Y(_14409_));
 sky130_fd_sc_hd__o2bb2a_1 _41664_ (.A1_N(_13630_),
    .A2_N(_13654_),
    .B1(_13653_),
    .B2(_13631_),
    .X(_14410_));
 sky130_fd_sc_hd__a21o_1 _41665_ (.A1(_04043_),
    .A2(_05697_),
    .B1(_12188_),
    .X(_14411_));
 sky130_fd_sc_hd__a21oi_1 _41666_ (.A1(_07425_),
    .A2(_13646_),
    .B1(_04047_),
    .Y(_14412_));
 sky130_fd_sc_hd__a21o_1 _41667_ (.A1(_08741_),
    .A2(_07421_),
    .B1(_14412_),
    .X(_14413_));
 sky130_fd_sc_hd__nand3_1 _41668_ (.A(_08741_),
    .B(_07421_),
    .C(_14412_),
    .Y(_14414_));
 sky130_fd_sc_hd__and3_1 _41669_ (.A(_14413_),
    .B(_14414_),
    .C(_08733_),
    .X(_14415_));
 sky130_fd_sc_hd__a21oi_1 _41670_ (.A1(_14413_),
    .A2(_14414_),
    .B1(_08733_),
    .Y(_14417_));
 sky130_fd_sc_hd__a211o_1 _41671_ (.A1(_13633_),
    .A2(_13643_),
    .B1(_14415_),
    .C1(_14417_),
    .X(_14418_));
 sky130_fd_sc_hd__o221ai_2 _41672_ (.A1(_12183_),
    .A2(_13632_),
    .B1(_14417_),
    .B2(_14415_),
    .C1(_13643_),
    .Y(_14419_));
 sky130_fd_sc_hd__a21o_1 _41673_ (.A1(_12199_),
    .A2(_12181_),
    .B1(_13646_),
    .X(_14420_));
 sky130_fd_sc_hd__o21a_1 _41674_ (.A1(_13635_),
    .A2(_13638_),
    .B1(_14420_),
    .X(_14421_));
 sky130_fd_sc_hd__a21oi_1 _41675_ (.A1(_14418_),
    .A2(_14419_),
    .B1(_14421_),
    .Y(_14422_));
 sky130_fd_sc_hd__and3_1 _41676_ (.A(_14418_),
    .B(_14419_),
    .C(_14421_),
    .X(_14423_));
 sky130_fd_sc_hd__a2111o_2 _41677_ (.A1(_13649_),
    .A2(_13650_),
    .B1(_14422_),
    .C1(_14423_),
    .D1(_13644_),
    .X(_14424_));
 sky130_fd_sc_hd__a21oi_1 _41678_ (.A1(_13649_),
    .A2(_13650_),
    .B1(_13644_),
    .Y(_14425_));
 sky130_fd_sc_hd__o21bai_1 _41679_ (.A1(_14422_),
    .A2(_14423_),
    .B1_N(_14425_),
    .Y(_14426_));
 sky130_fd_sc_hd__nand2_2 _41680_ (.A(_14424_),
    .B(_14426_),
    .Y(_14428_));
 sky130_fd_sc_hd__xor2_1 _41681_ (.A(_14411_),
    .B(_14428_),
    .X(_14429_));
 sky130_fd_sc_hd__xnor2_1 _41682_ (.A(_14410_),
    .B(_14429_),
    .Y(_14430_));
 sky130_fd_sc_hd__a21oi_1 _41683_ (.A1(_13629_),
    .A2(_13659_),
    .B1(_13656_),
    .Y(_14431_));
 sky130_fd_sc_hd__nor2_1 _41684_ (.A(_14430_),
    .B(_14431_),
    .Y(_14432_));
 sky130_fd_sc_hd__nand2_1 _41685_ (.A(_13629_),
    .B(_13659_),
    .Y(_14433_));
 sky130_fd_sc_hd__and3b_1 _41686_ (.A_N(_13656_),
    .B(_14433_),
    .C(_14430_),
    .X(_14434_));
 sky130_fd_sc_hd__o221a_1 _41687_ (.A1(_12223_),
    .A2(_12243_),
    .B1(_13612_),
    .B2(_13615_),
    .C1(_12244_),
    .X(_14435_));
 sky130_fd_sc_hd__o41ai_2 _41688_ (.A1(_11013_),
    .A2(_12219_),
    .A3(_13600_),
    .A4(_14435_),
    .B1(_13618_),
    .Y(_14436_));
 sky130_fd_sc_hd__clkbuf_2 _41689_ (.A(_13610_),
    .X(_14437_));
 sky130_fd_sc_hd__buf_1 _41690_ (.A(_12232_),
    .X(_14439_));
 sky130_fd_sc_hd__nand2_1 _41691_ (.A(_14439_),
    .B(_13605_),
    .Y(_14440_));
 sky130_fd_sc_hd__nand2_1 _41692_ (.A(_09764_),
    .B(_12225_),
    .Y(_14441_));
 sky130_fd_sc_hd__o22ai_1 _41693_ (.A1(_14441_),
    .A2(_13610_),
    .B1(_12225_),
    .B2(_13601_),
    .Y(_14442_));
 sky130_fd_sc_hd__buf_1 _41694_ (.A(_14442_),
    .X(_14443_));
 sky130_fd_sc_hd__a21bo_1 _41695_ (.A1(_14440_),
    .A2(_12234_),
    .B1_N(_14443_),
    .X(_14444_));
 sky130_fd_sc_hd__a211o_1 _41696_ (.A1(_14439_),
    .A2(_13605_),
    .B1(_14442_),
    .C1(_12226_),
    .X(_14445_));
 sky130_fd_sc_hd__and4_1 _41697_ (.A(_13604_),
    .B(_14444_),
    .C(_14445_),
    .D(_14437_),
    .X(_14446_));
 sky130_fd_sc_hd__a22oi_2 _41698_ (.A1(_14437_),
    .A2(_13604_),
    .B1(_14444_),
    .B2(_14445_),
    .Y(_14447_));
 sky130_fd_sc_hd__o2111ai_2 _41699_ (.A1(_11012_),
    .A2(_14437_),
    .B1(_13609_),
    .C1(_12222_),
    .D1(_13608_),
    .Y(_14448_));
 sky130_fd_sc_hd__o211ai_2 _41700_ (.A1(_14446_),
    .A2(_14447_),
    .B1(_13608_),
    .C1(_14448_),
    .Y(_14450_));
 sky130_fd_sc_hd__a211o_1 _41701_ (.A1(_13608_),
    .A2(_14448_),
    .B1(_14446_),
    .C1(_14447_),
    .X(_14451_));
 sky130_fd_sc_hd__o311a_1 _41702_ (.A1(_12219_),
    .A2(_14437_),
    .A3(_12227_),
    .B1(_14450_),
    .C1(_14451_),
    .X(_14452_));
 sky130_fd_sc_hd__a21oi_1 _41703_ (.A1(_14451_),
    .A2(_14450_),
    .B1(_13611_),
    .Y(_14453_));
 sky130_fd_sc_hd__or2_1 _41704_ (.A(_14452_),
    .B(_14453_),
    .X(_14454_));
 sky130_fd_sc_hd__xnor2_1 _41705_ (.A(_14436_),
    .B(_14454_),
    .Y(_14455_));
 sky130_fd_sc_hd__a21oi_1 _41706_ (.A1(_13623_),
    .A2(_13627_),
    .B1(_14455_),
    .Y(_14456_));
 sky130_fd_sc_hd__nand3_1 _41707_ (.A(_13623_),
    .B(_13627_),
    .C(_14455_),
    .Y(_14457_));
 sky130_fd_sc_hd__and2b_1 _41708_ (.A_N(_14456_),
    .B(_14457_),
    .X(_14458_));
 sky130_fd_sc_hd__o21bai_2 _41709_ (.A1(_14432_),
    .A2(_14434_),
    .B1_N(_14458_),
    .Y(_14459_));
 sky130_fd_sc_hd__a21o_1 _41710_ (.A1(_13688_),
    .A2(_12260_),
    .B1(_07350_),
    .X(_14461_));
 sky130_fd_sc_hd__clkbuf_2 _41711_ (.A(_11048_),
    .X(_14462_));
 sky130_fd_sc_hd__a21oi_1 _41712_ (.A1(_13688_),
    .A2(_14462_),
    .B1(_13664_),
    .Y(_14463_));
 sky130_fd_sc_hd__a21oi_1 _41713_ (.A1(_12266_),
    .A2(_14461_),
    .B1(_14463_),
    .Y(_14464_));
 sky130_fd_sc_hd__and3b_1 _41714_ (.A_N(_11049_),
    .B(_11050_),
    .C(_13667_),
    .X(_14465_));
 sky130_fd_sc_hd__mux2_1 _41715_ (.A0(_11048_),
    .A1(_07336_),
    .S(_09846_),
    .X(_14466_));
 sky130_fd_sc_hd__or3_1 _41716_ (.A(_07332_),
    .B(_07333_),
    .C(_14466_),
    .X(_14467_));
 sky130_fd_sc_hd__o21ai_1 _41717_ (.A1(_07332_),
    .A2(_07333_),
    .B1(_14466_),
    .Y(_14468_));
 sky130_fd_sc_hd__clkbuf_2 _41718_ (.A(_11050_),
    .X(_14469_));
 sky130_fd_sc_hd__nand4_2 _41719_ (.A(_14467_),
    .B(_14468_),
    .C(_11049_),
    .D(_14469_),
    .Y(_14470_));
 sky130_fd_sc_hd__a22o_1 _41720_ (.A1(_11049_),
    .A2(_14469_),
    .B1(_14467_),
    .B2(_14468_),
    .X(_14472_));
 sky130_fd_sc_hd__o211a_1 _41721_ (.A1(_14465_),
    .A2(_13675_),
    .B1(_14470_),
    .C1(_14472_),
    .X(_14473_));
 sky130_fd_sc_hd__a211oi_1 _41722_ (.A1(_14470_),
    .A2(_14472_),
    .B1(_14465_),
    .C1(_13675_),
    .Y(_14474_));
 sky130_fd_sc_hd__nor2_1 _41723_ (.A(_14473_),
    .B(_14474_),
    .Y(_14475_));
 sky130_fd_sc_hd__xnor2_1 _41724_ (.A(_14464_),
    .B(_14475_),
    .Y(_14476_));
 sky130_fd_sc_hd__or3_2 _41725_ (.A(_13676_),
    .B(_13681_),
    .C(_14476_),
    .X(_14477_));
 sky130_fd_sc_hd__o21ai_1 _41726_ (.A1(_13676_),
    .A2(_13681_),
    .B1(_14476_),
    .Y(_14478_));
 sky130_fd_sc_hd__o221a_1 _41727_ (.A1(_11069_),
    .A2(_13664_),
    .B1(_04099_),
    .B2(_07350_),
    .C1(_13688_),
    .X(_14479_));
 sky130_fd_sc_hd__nand3_1 _41728_ (.A(_14477_),
    .B(_14478_),
    .C(_14479_),
    .Y(_14480_));
 sky130_fd_sc_hd__a21o_1 _41729_ (.A1(_14477_),
    .A2(_14478_),
    .B1(_14479_),
    .X(_14481_));
 sky130_fd_sc_hd__and2_1 _41730_ (.A(_14480_),
    .B(_14481_),
    .X(_14483_));
 sky130_fd_sc_hd__o21a_1 _41731_ (.A1(_13684_),
    .A2(_13687_),
    .B1(_14483_),
    .X(_14484_));
 sky130_fd_sc_hd__a211oi_1 _41732_ (.A1(_13689_),
    .A2(_13686_),
    .B1(_14483_),
    .C1(_13684_),
    .Y(_14485_));
 sky130_fd_sc_hd__nor2_1 _41733_ (.A(_14484_),
    .B(_14485_),
    .Y(_14486_));
 sky130_fd_sc_hd__a21oi_2 _41734_ (.A1(_13696_),
    .A2(_13694_),
    .B1(_13693_),
    .Y(_14487_));
 sky130_fd_sc_hd__xor2_2 _41735_ (.A(_14486_),
    .B(_14487_),
    .X(_14488_));
 sky130_fd_sc_hd__nand2_4 _41736_ (.A(_14459_),
    .B(_14488_),
    .Y(_14489_));
 sky130_fd_sc_hd__inv_2 _41737_ (.A(_14489_),
    .Y(_14490_));
 sky130_fd_sc_hd__or3b_4 _41738_ (.A(_14432_),
    .B(_14434_),
    .C_N(_14458_),
    .X(_14491_));
 sky130_fd_sc_hd__a21oi_1 _41739_ (.A1(_14459_),
    .A2(_14491_),
    .B1(_14488_),
    .Y(_14492_));
 sky130_fd_sc_hd__a21o_1 _41740_ (.A1(_14490_),
    .A2(_14491_),
    .B1(_14492_),
    .X(_14494_));
 sky130_fd_sc_hd__and3_2 _41741_ (.A(_14407_),
    .B(_14408_),
    .C(_14406_),
    .X(_14495_));
 sky130_fd_sc_hd__nor3_4 _41742_ (.A(_14409_),
    .B(_14494_),
    .C(_14495_),
    .Y(_14496_));
 sky130_fd_sc_hd__o21a_1 _41743_ (.A1(_14409_),
    .A2(_14495_),
    .B1(_14494_),
    .X(_14497_));
 sky130_fd_sc_hd__or3_4 _41744_ (.A(_14351_),
    .B(_14496_),
    .C(_14497_),
    .X(_14498_));
 sky130_fd_sc_hd__o221ai_4 _41745_ (.A1(_13597_),
    .A2(_13698_),
    .B1(_14496_),
    .B2(_14497_),
    .C1(_13598_),
    .Y(_14499_));
 sky130_fd_sc_hd__nand2_1 _41746_ (.A(_14498_),
    .B(net72),
    .Y(_14500_));
 sky130_fd_sc_hd__nor2_1 _41747_ (.A(_14349_),
    .B(_14500_),
    .Y(_14501_));
 sky130_fd_sc_hd__and2_1 _41748_ (.A(_14500_),
    .B(_14349_),
    .X(_14502_));
 sky130_fd_sc_hd__nor4_1 _41749_ (.A(_13700_),
    .B(_13704_),
    .C(_14501_),
    .D(_14502_),
    .Y(_14503_));
 sky130_fd_sc_hd__o22a_1 _41750_ (.A1(_13700_),
    .A2(_13704_),
    .B1(_14501_),
    .B2(_14502_),
    .X(_14505_));
 sky130_fd_sc_hd__nor2_1 _41751_ (.A(_14503_),
    .B(_14505_),
    .Y(_14506_));
 sky130_fd_sc_hd__o21ai_4 _41752_ (.A1(_13309_),
    .A2(_13360_),
    .B1(_13417_),
    .Y(_14507_));
 sky130_fd_sc_hd__nor2_1 _41753_ (.A(_13366_),
    .B(_05413_),
    .Y(_14508_));
 sky130_fd_sc_hd__nand2_1 _41754_ (.A(_05413_),
    .B(_13366_),
    .Y(_14509_));
 sky130_fd_sc_hd__and2b_1 _41755_ (.A_N(_14508_),
    .B(_14509_),
    .X(_14510_));
 sky130_fd_sc_hd__and3_1 _41756_ (.A(_11382_),
    .B(_13369_),
    .C(_14510_),
    .X(_14511_));
 sky130_fd_sc_hd__buf_1 _41757_ (.A(_11382_),
    .X(_14512_));
 sky130_fd_sc_hd__a21oi_1 _41758_ (.A1(_14512_),
    .A2(_13369_),
    .B1(_14510_),
    .Y(_14513_));
 sky130_fd_sc_hd__o21ai_1 _41759_ (.A1(_14511_),
    .A2(_14513_),
    .B1(_13367_),
    .Y(_14514_));
 sky130_fd_sc_hd__inv_2 _41760_ (.A(_13369_),
    .Y(_14516_));
 sky130_fd_sc_hd__a31o_1 _41761_ (.A1(_14512_),
    .A2(_12544_),
    .A3(_14516_),
    .B1(_13374_),
    .X(_14517_));
 sky130_fd_sc_hd__and2_1 _41762_ (.A(_14514_),
    .B(_14517_),
    .X(_14518_));
 sky130_fd_sc_hd__nor2_1 _41763_ (.A(_14514_),
    .B(_14517_),
    .Y(_14519_));
 sky130_fd_sc_hd__or2_1 _41764_ (.A(_14518_),
    .B(_14519_),
    .X(_14520_));
 sky130_fd_sc_hd__inv_2 _41765_ (.A(_14520_),
    .Y(_14521_));
 sky130_fd_sc_hd__o21a_1 _41766_ (.A1(_13380_),
    .A2(_13384_),
    .B1(_14521_),
    .X(_14522_));
 sky130_fd_sc_hd__nor3_1 _41767_ (.A(_13380_),
    .B(_13384_),
    .C(_14521_),
    .Y(_14523_));
 sky130_fd_sc_hd__or2_1 _41768_ (.A(_14522_),
    .B(_14523_),
    .X(_14524_));
 sky130_fd_sc_hd__o21ba_1 _41769_ (.A1(_13384_),
    .A2(_14521_),
    .B1_N(_13377_),
    .X(_14525_));
 sky130_fd_sc_hd__a21oi_4 _41770_ (.A1(_13377_),
    .A2(_14524_),
    .B1(_14525_),
    .Y(_14527_));
 sky130_fd_sc_hd__a21o_1 _41771_ (.A1(_13395_),
    .A2(_12539_),
    .B1(_13409_),
    .X(_14528_));
 sky130_fd_sc_hd__or3_1 _41772_ (.A(_08902_),
    .B(_11410_),
    .C(_11414_),
    .X(_14529_));
 sky130_fd_sc_hd__o21ai_1 _41773_ (.A1(_08902_),
    .A2(_11414_),
    .B1(_11410_),
    .Y(_14530_));
 sky130_fd_sc_hd__nand2_1 _41774_ (.A(_14529_),
    .B(_14530_),
    .Y(_14531_));
 sky130_fd_sc_hd__nand2_1 _41775_ (.A(_13396_),
    .B(_14531_),
    .Y(_14532_));
 sky130_fd_sc_hd__or3_1 _41776_ (.A(_13399_),
    .B(_14532_),
    .C(_13401_),
    .X(_14533_));
 sky130_fd_sc_hd__a2bb2o_1 _41777_ (.A1_N(_13399_),
    .A2_N(_13401_),
    .B1(_14531_),
    .B2(_13396_),
    .X(_14534_));
 sky130_fd_sc_hd__and2_1 _41778_ (.A(_14533_),
    .B(_14534_),
    .X(_14535_));
 sky130_fd_sc_hd__o31a_1 _41779_ (.A1(_13401_),
    .A2(_13402_),
    .A3(_13404_),
    .B1(_14535_),
    .X(_14536_));
 sky130_fd_sc_hd__nor3b_2 _41780_ (.A(_13404_),
    .B(_14535_),
    .C_N(_13403_),
    .Y(_14538_));
 sky130_fd_sc_hd__o2bb2ai_4 _41781_ (.A1_N(_13407_),
    .A2_N(_14528_),
    .B1(_14536_),
    .B2(_14538_),
    .Y(_14539_));
 sky130_fd_sc_hd__a2111o_2 _41782_ (.A1(_12531_),
    .A2(_13406_),
    .B1(_13410_),
    .C1(_14536_),
    .D1(_14538_),
    .X(_14540_));
 sky130_fd_sc_hd__nand3_1 _41783_ (.A(_11442_),
    .B(_06941_),
    .C(\delay_line[29][14] ),
    .Y(_14541_));
 sky130_fd_sc_hd__a22o_1 _41784_ (.A1(_14541_),
    .A2(_11443_),
    .B1(_13390_),
    .B2(_13391_),
    .X(_14542_));
 sky130_fd_sc_hd__a21boi_4 _41785_ (.A1(_14539_),
    .A2(_14540_),
    .B1_N(_14542_),
    .Y(_14543_));
 sky130_fd_sc_hd__clkbuf_2 _41786_ (.A(_14542_),
    .X(_14544_));
 sky130_fd_sc_hd__nand3b_2 _41787_ (.A_N(_14544_),
    .B(_14539_),
    .C(_14540_),
    .Y(_14545_));
 sky130_fd_sc_hd__and2b_1 _41788_ (.A_N(_14543_),
    .B(_14545_),
    .X(_14546_));
 sky130_fd_sc_hd__or2_1 _41789_ (.A(_14527_),
    .B(_14546_),
    .X(_14547_));
 sky130_fd_sc_hd__nand2_1 _41790_ (.A(_14527_),
    .B(_14546_),
    .Y(_14549_));
 sky130_fd_sc_hd__buf_1 _41791_ (.A(_13318_),
    .X(_14550_));
 sky130_fd_sc_hd__a21oi_1 _41792_ (.A1(_14550_),
    .A2(_05500_),
    .B1(_07042_),
    .Y(_14551_));
 sky130_fd_sc_hd__o21ai_1 _41793_ (.A1(_05497_),
    .A2(_05499_),
    .B1(_14550_),
    .Y(_14552_));
 sky130_fd_sc_hd__o21ai_1 _41794_ (.A1(_12568_),
    .A2(_14552_),
    .B1(_13322_),
    .Y(_14553_));
 sky130_fd_sc_hd__a311o_1 _41795_ (.A1(_14550_),
    .A2(_05499_),
    .A3(_07039_),
    .B1(_14551_),
    .C1(_14553_),
    .X(_14554_));
 sky130_fd_sc_hd__a31o_1 _41796_ (.A1(_14550_),
    .A2(_05499_),
    .A3(_07039_),
    .B1(_14551_),
    .X(_14555_));
 sky130_fd_sc_hd__nand2_1 _41797_ (.A(_14555_),
    .B(_14553_),
    .Y(_14556_));
 sky130_fd_sc_hd__and2_1 _41798_ (.A(_14554_),
    .B(_14556_),
    .X(_14557_));
 sky130_fd_sc_hd__xor2_1 _41799_ (.A(_13325_),
    .B(_14557_),
    .X(_14558_));
 sky130_fd_sc_hd__nor3b_1 _41800_ (.A(_13331_),
    .B(_13330_),
    .C_N(_14558_),
    .Y(_14560_));
 sky130_fd_sc_hd__o21ba_1 _41801_ (.A1(_13331_),
    .A2(_13330_),
    .B1_N(_14558_),
    .X(_14561_));
 sky130_fd_sc_hd__or4bb_1 _41802_ (.A(_13342_),
    .B(_13343_),
    .C_N(_12579_),
    .D_N(_13334_),
    .X(_14562_));
 sky130_fd_sc_hd__and2_1 _41803_ (.A(_12590_),
    .B(_13344_),
    .X(_14563_));
 sky130_fd_sc_hd__or2_1 _41804_ (.A(_05529_),
    .B(_13340_),
    .X(_14564_));
 sky130_fd_sc_hd__a21o_1 _41805_ (.A1(_10146_),
    .A2(_13337_),
    .B1(_11337_),
    .X(_14565_));
 sky130_fd_sc_hd__a22o_1 _41806_ (.A1(_12584_),
    .A2(_08802_),
    .B1(_14564_),
    .B2(_14565_),
    .X(_14566_));
 sky130_fd_sc_hd__o31a_1 _41807_ (.A1(_05529_),
    .A2(_07015_),
    .A3(_08803_),
    .B1(_14566_),
    .X(_14567_));
 sky130_fd_sc_hd__o21a_1 _41808_ (.A1(_13343_),
    .A2(_14563_),
    .B1(_14567_),
    .X(_14568_));
 sky130_fd_sc_hd__a311oi_1 _41809_ (.A1(_13341_),
    .A2(_13338_),
    .A3(_13340_),
    .B1(_14567_),
    .C1(_14563_),
    .Y(_14569_));
 sky130_fd_sc_hd__or3_1 _41810_ (.A(_11336_),
    .B(_14568_),
    .C(_14569_),
    .X(_14571_));
 sky130_fd_sc_hd__clkbuf_2 _41811_ (.A(_11336_),
    .X(_14572_));
 sky130_fd_sc_hd__o21ai_1 _41812_ (.A1(_14568_),
    .A2(_14569_),
    .B1(_14572_),
    .Y(_14573_));
 sky130_fd_sc_hd__nand2_1 _41813_ (.A(_14571_),
    .B(_14573_),
    .Y(_14574_));
 sky130_fd_sc_hd__a21oi_1 _41814_ (.A1(_13347_),
    .A2(_14562_),
    .B1(_14574_),
    .Y(_14575_));
 sky130_fd_sc_hd__and3_1 _41815_ (.A(_13347_),
    .B(_14574_),
    .C(_14562_),
    .X(_14576_));
 sky130_fd_sc_hd__nor2_1 _41816_ (.A(_14575_),
    .B(_14576_),
    .Y(_14577_));
 sky130_fd_sc_hd__inv_2 _41817_ (.A(_13349_),
    .Y(_14578_));
 sky130_fd_sc_hd__o21a_1 _41818_ (.A1(_14578_),
    .A2(_13353_),
    .B1(_13351_),
    .X(_14579_));
 sky130_fd_sc_hd__xor2_1 _41819_ (.A(_14577_),
    .B(_14579_),
    .X(_14580_));
 sky130_fd_sc_hd__o21a_1 _41820_ (.A1(_14560_),
    .A2(_14561_),
    .B1(_14580_),
    .X(_14582_));
 sky130_fd_sc_hd__nor3_1 _41821_ (.A(_14580_),
    .B(_14560_),
    .C(_14561_),
    .Y(_14583_));
 sky130_fd_sc_hd__nor2_1 _41822_ (.A(_14582_),
    .B(_14583_),
    .Y(_14584_));
 sky130_fd_sc_hd__o21a_1 _41823_ (.A1(_12558_),
    .A2(_13310_),
    .B1(_08784_),
    .X(_14585_));
 sky130_fd_sc_hd__or3_2 _41824_ (.A(_13311_),
    .B(_14585_),
    .C(_13315_),
    .X(_14586_));
 sky130_fd_sc_hd__xnor2_1 _41825_ (.A(_14584_),
    .B(_14586_),
    .Y(_14587_));
 sky130_fd_sc_hd__o211ai_2 _41826_ (.A1(_13333_),
    .A2(_13356_),
    .B1(_13359_),
    .C1(_14587_),
    .Y(_14588_));
 sky130_fd_sc_hd__o21ai_1 _41827_ (.A1(_13333_),
    .A2(_13356_),
    .B1(_13359_),
    .Y(_14589_));
 sky130_fd_sc_hd__or2b_1 _41828_ (.A(_14587_),
    .B_N(_14589_),
    .X(_14590_));
 sky130_fd_sc_hd__nand2_1 _41829_ (.A(_14588_),
    .B(_14590_),
    .Y(_14591_));
 sky130_fd_sc_hd__a21bo_1 _41830_ (.A1(_14547_),
    .A2(_14549_),
    .B1_N(_14591_),
    .X(_14593_));
 sky130_fd_sc_hd__nand3b_1 _41831_ (.A_N(_14591_),
    .B(_14547_),
    .C(_14549_),
    .Y(_14594_));
 sky130_fd_sc_hd__o211a_1 _41832_ (.A1(_13513_),
    .A2(_13514_),
    .B1(_14593_),
    .C1(_14594_),
    .X(_14595_));
 sky130_fd_sc_hd__a211oi_1 _41833_ (.A1(_14593_),
    .A2(_14594_),
    .B1(_13513_),
    .C1(_13514_),
    .Y(_14596_));
 sky130_fd_sc_hd__nor2_1 _41834_ (.A(_14595_),
    .B(_14596_),
    .Y(_14597_));
 sky130_fd_sc_hd__xnor2_2 _41835_ (.A(_14507_),
    .B(_14597_),
    .Y(_14598_));
 sky130_fd_sc_hd__xnor2_1 _41836_ (.A(_14506_),
    .B(_14598_),
    .Y(_14599_));
 sky130_fd_sc_hd__xnor2_1 _41837_ (.A(_14272_),
    .B(_14599_),
    .Y(_14600_));
 sky130_fd_sc_hd__a21bo_1 _41838_ (.A1(_13806_),
    .A2(_13782_),
    .B1_N(_13783_),
    .X(_14601_));
 sky130_fd_sc_hd__nand3_1 _41839_ (.A(_13422_),
    .B(_13419_),
    .C(_13421_),
    .Y(_14602_));
 sky130_fd_sc_hd__nand2_1 _41840_ (.A(_11580_),
    .B(_13793_),
    .Y(_14604_));
 sky130_fd_sc_hd__clkbuf_2 _41841_ (.A(_13785_),
    .X(_14605_));
 sky130_fd_sc_hd__nand2_1 _41842_ (.A(_05319_),
    .B(_05314_),
    .Y(_14606_));
 sky130_fd_sc_hd__a2bb2o_1 _41843_ (.A1_N(_13789_),
    .A2_N(_13787_),
    .B1(_14606_),
    .B2(_11568_),
    .X(_14607_));
 sky130_fd_sc_hd__nor2_1 _41844_ (.A(_14605_),
    .B(_14607_),
    .Y(_14608_));
 sky130_fd_sc_hd__and2_1 _41845_ (.A(_14605_),
    .B(_14607_),
    .X(_14609_));
 sky130_fd_sc_hd__o21ai_1 _41846_ (.A1(_14608_),
    .A2(_14609_),
    .B1(_11580_),
    .Y(_14610_));
 sky130_fd_sc_hd__or3_1 _41847_ (.A(_12696_),
    .B(_14608_),
    .C(_14609_),
    .X(_14611_));
 sky130_fd_sc_hd__a22oi_2 _41848_ (.A1(_13792_),
    .A2(_14604_),
    .B1(_14610_),
    .B2(_14611_),
    .Y(_14612_));
 sky130_fd_sc_hd__and4_1 _41849_ (.A(_13792_),
    .B(_14604_),
    .C(_14610_),
    .D(_14611_),
    .X(_14613_));
 sky130_fd_sc_hd__o22a_1 _41850_ (.A1(_13800_),
    .A2(_13802_),
    .B1(_14612_),
    .B2(_14613_),
    .X(_14615_));
 sky130_fd_sc_hd__nor4_1 _41851_ (.A(_14215_),
    .B(_13802_),
    .C(_14612_),
    .D(_14613_),
    .Y(_14616_));
 sky130_fd_sc_hd__or2_2 _41852_ (.A(_14615_),
    .B(_14616_),
    .X(_14617_));
 sky130_fd_sc_hd__nand2_2 _41853_ (.A(_13776_),
    .B(_13780_),
    .Y(_14618_));
 sky130_fd_sc_hd__a21oi_1 _41854_ (.A1(_13769_),
    .A2(_13761_),
    .B1(_13773_),
    .Y(_14619_));
 sky130_fd_sc_hd__a21oi_1 _41855_ (.A1(_12653_),
    .A2(_12655_),
    .B1(_13732_),
    .Y(_14620_));
 sky130_fd_sc_hd__a22o_1 _41856_ (.A1(_09582_),
    .A2(_05203_),
    .B1(_13718_),
    .B2(_12633_),
    .X(_14621_));
 sky130_fd_sc_hd__a2bb2o_1 _41857_ (.A1_N(_13722_),
    .A2_N(_13725_),
    .B1(_14621_),
    .B2(_13721_),
    .X(_14622_));
 sky130_fd_sc_hd__nand2_1 _41858_ (.A(_13721_),
    .B(_14621_),
    .Y(_14623_));
 sky130_fd_sc_hd__or3_1 _41859_ (.A(_13722_),
    .B(_14623_),
    .C(_13725_),
    .X(_14624_));
 sky130_fd_sc_hd__nand2_1 _41860_ (.A(_14622_),
    .B(_14624_),
    .Y(_14626_));
 sky130_fd_sc_hd__o21bai_2 _41861_ (.A1(net151),
    .A2(_14620_),
    .B1_N(_14626_),
    .Y(_14627_));
 sky130_fd_sc_hd__nand3b_1 _41862_ (.A_N(net151),
    .B(_13733_),
    .C(_14626_),
    .Y(_14628_));
 sky130_fd_sc_hd__a21oi_1 _41863_ (.A1(_14627_),
    .A2(_14628_),
    .B1(_13727_),
    .Y(_14629_));
 sky130_fd_sc_hd__a21bo_1 _41864_ (.A1(_13733_),
    .A2(_14626_),
    .B1_N(_13727_),
    .X(_14630_));
 sky130_fd_sc_hd__or3b_1 _41865_ (.A(_13738_),
    .B(_13739_),
    .C_N(_13740_),
    .X(_14631_));
 sky130_fd_sc_hd__o21ai_1 _41866_ (.A1(_11496_),
    .A2(_08331_),
    .B1(_13740_),
    .Y(_14632_));
 sky130_fd_sc_hd__o211ai_2 _41867_ (.A1(_09633_),
    .A2(_13738_),
    .B1(_13739_),
    .C1(_14632_),
    .Y(_14633_));
 sky130_fd_sc_hd__a221oi_1 _41868_ (.A1(_14631_),
    .A2(_14633_),
    .B1(_13750_),
    .B2(_13742_),
    .C1(_13748_),
    .Y(_14634_));
 sky130_fd_sc_hd__nand2_1 _41869_ (.A(_14631_),
    .B(_14633_),
    .Y(_14635_));
 sky130_fd_sc_hd__a21oi_1 _41870_ (.A1(_13750_),
    .A2(_13742_),
    .B1(_13748_),
    .Y(_14637_));
 sky130_fd_sc_hd__nor2_1 _41871_ (.A(_14635_),
    .B(_14637_),
    .Y(_14638_));
 sky130_fd_sc_hd__nor2_1 _41872_ (.A(_14634_),
    .B(_14638_),
    .Y(_14639_));
 sky130_fd_sc_hd__xor2_1 _41873_ (.A(_13752_),
    .B(_14639_),
    .X(_14640_));
 sky130_fd_sc_hd__a21oi_1 _41874_ (.A1(_12673_),
    .A2(_13754_),
    .B1(_13758_),
    .Y(_14641_));
 sky130_fd_sc_hd__or2_1 _41875_ (.A(_14640_),
    .B(_14641_),
    .X(_14642_));
 sky130_fd_sc_hd__nand2_1 _41876_ (.A(_14641_),
    .B(_14640_),
    .Y(_14643_));
 sky130_fd_sc_hd__and2_1 _41877_ (.A(_14642_),
    .B(_14643_),
    .X(_14644_));
 sky130_fd_sc_hd__nand3b_1 _41878_ (.A_N(_14629_),
    .B(_14630_),
    .C(_14644_),
    .Y(_14645_));
 sky130_fd_sc_hd__a21boi_1 _41879_ (.A1(_13733_),
    .A2(_14626_),
    .B1_N(_13727_),
    .Y(_14646_));
 sky130_fd_sc_hd__o21bai_1 _41880_ (.A1(_14629_),
    .A2(_14646_),
    .B1_N(_14644_),
    .Y(_14648_));
 sky130_fd_sc_hd__a21bo_1 _41881_ (.A1(_06786_),
    .A2(_08295_),
    .B1_N(_11476_),
    .X(_14649_));
 sky130_fd_sc_hd__o211a_1 _41882_ (.A1(_11477_),
    .A2(_06780_),
    .B1(_06785_),
    .C1(_12623_),
    .X(_14650_));
 sky130_fd_sc_hd__a21o_1 _41883_ (.A1(_08292_),
    .A2(_14649_),
    .B1(_14650_),
    .X(_14651_));
 sky130_fd_sc_hd__and2_1 _41884_ (.A(_08292_),
    .B(_14649_),
    .X(_14652_));
 sky130_fd_sc_hd__o21ai_1 _41885_ (.A1(_14650_),
    .A2(_13767_),
    .B1(_14652_),
    .Y(_14653_));
 sky130_fd_sc_hd__o21a_1 _41886_ (.A1(_13767_),
    .A2(_14651_),
    .B1(_14653_),
    .X(_14654_));
 sky130_fd_sc_hd__a21o_1 _41887_ (.A1(_14645_),
    .A2(_14648_),
    .B1(_14654_),
    .X(_14655_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41888_ (.A(_14645_),
    .X(_14656_));
 sky130_fd_sc_hd__nand3_1 _41889_ (.A(_14654_),
    .B(_14648_),
    .C(_14656_),
    .Y(_14657_));
 sky130_fd_sc_hd__inv_2 _41890_ (.A(_13386_),
    .Y(_14659_));
 sky130_fd_sc_hd__o32a_2 _41891_ (.A1(_13392_),
    .A2(_13410_),
    .A3(_13411_),
    .B1(_13413_),
    .B2(_14659_),
    .X(_14660_));
 sky130_fd_sc_hd__a21bo_1 _41892_ (.A1(_14655_),
    .A2(_14657_),
    .B1_N(_14660_),
    .X(_14661_));
 sky130_fd_sc_hd__a21oi_1 _41893_ (.A1(_14656_),
    .A2(_14648_),
    .B1(_14654_),
    .Y(_14662_));
 sky130_fd_sc_hd__nor2_1 _41894_ (.A(_14660_),
    .B(_14662_),
    .Y(_14663_));
 sky130_fd_sc_hd__buf_1 _41895_ (.A(_14657_),
    .X(_14664_));
 sky130_fd_sc_hd__nand2_1 _41896_ (.A(_14663_),
    .B(_14664_),
    .Y(_14665_));
 sky130_fd_sc_hd__nand3b_4 _41897_ (.A_N(_14619_),
    .B(_14661_),
    .C(_14665_),
    .Y(_14666_));
 sky130_fd_sc_hd__a21bo_2 _41898_ (.A1(_14661_),
    .A2(_14665_),
    .B1_N(_14619_),
    .X(_14667_));
 sky130_fd_sc_hd__and3_1 _41899_ (.A(_14618_),
    .B(_14666_),
    .C(_14667_),
    .X(_14668_));
 sky130_fd_sc_hd__a21oi_4 _41900_ (.A1(_14666_),
    .A2(_14667_),
    .B1(_14618_),
    .Y(_14670_));
 sky130_fd_sc_hd__nor2_2 _41901_ (.A(_14668_),
    .B(_14670_),
    .Y(_14671_));
 sky130_fd_sc_hd__xor2_1 _41902_ (.A(_14617_),
    .B(_14671_),
    .X(_14672_));
 sky130_fd_sc_hd__nand3_2 _41903_ (.A(_13421_),
    .B(_14602_),
    .C(_14672_),
    .Y(_14673_));
 sky130_fd_sc_hd__a21o_1 _41904_ (.A1(_13421_),
    .A2(_14602_),
    .B1(_14672_),
    .X(_14674_));
 sky130_fd_sc_hd__nand2_1 _41905_ (.A(_14673_),
    .B(_14674_),
    .Y(_14675_));
 sky130_fd_sc_hd__xor2_1 _41906_ (.A(_14601_),
    .B(_14675_),
    .X(_14676_));
 sky130_fd_sc_hd__xnor2_1 _41907_ (.A(_14600_),
    .B(_14676_),
    .Y(_14677_));
 sky130_fd_sc_hd__o311a_1 _41908_ (.A1(_13712_),
    .A2(_13811_),
    .A3(_13813_),
    .B1(_14677_),
    .C1(_13711_),
    .X(_14678_));
 sky130_fd_sc_hd__o31a_1 _41909_ (.A1(_13811_),
    .A2(_13813_),
    .A3(_13712_),
    .B1(_13711_),
    .X(_14679_));
 sky130_fd_sc_hd__nor2_1 _41910_ (.A(_14679_),
    .B(_14677_),
    .Y(_14681_));
 sky130_fd_sc_hd__nor2_1 _41911_ (.A(_14678_),
    .B(_14681_),
    .Y(_14682_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _41912_ (.A(_14682_),
    .X(_14683_));
 sky130_fd_sc_hd__a21oi_2 _41913_ (.A1(_14255_),
    .A2(_14270_),
    .B1(_14683_),
    .Y(_14684_));
 sky130_fd_sc_hd__o21ai_1 _41914_ (.A1(_13815_),
    .A2(_13816_),
    .B1(_13819_),
    .Y(_14685_));
 sky130_fd_sc_hd__nand3_1 _41915_ (.A(_14255_),
    .B(_14270_),
    .C(_14683_),
    .Y(_14686_));
 sky130_fd_sc_hd__nand2_1 _41916_ (.A(_14685_),
    .B(_14686_),
    .Y(_14687_));
 sky130_fd_sc_hd__a21oi_1 _41917_ (.A1(_14267_),
    .A2(_14268_),
    .B1(_14256_),
    .Y(_14688_));
 sky130_fd_sc_hd__nand2_1 _41918_ (.A(_14256_),
    .B(_14268_),
    .Y(_14689_));
 sky130_fd_sc_hd__nor2_1 _41919_ (.A(_14247_),
    .B(_14689_),
    .Y(_14690_));
 sky130_fd_sc_hd__o21ai_1 _41920_ (.A1(_14688_),
    .A2(_14690_),
    .B1(_14683_),
    .Y(_14692_));
 sky130_fd_sc_hd__o21a_1 _41921_ (.A1(_13815_),
    .A2(_13816_),
    .B1(_13819_),
    .X(_14693_));
 sky130_fd_sc_hd__nand3b_1 _41922_ (.A_N(_14682_),
    .B(_14255_),
    .C(_14270_),
    .Y(_14694_));
 sky130_fd_sc_hd__nand3_2 _41923_ (.A(_14692_),
    .B(_14693_),
    .C(_14694_),
    .Y(_14695_));
 sky130_fd_sc_hd__o21ai_1 _41924_ (.A1(_14684_),
    .A2(_14687_),
    .B1(_14695_),
    .Y(_14696_));
 sky130_fd_sc_hd__nand2_1 _41925_ (.A(_13304_),
    .B(_13303_),
    .Y(_14697_));
 sky130_fd_sc_hd__a31o_1 _41926_ (.A1(_12783_),
    .A2(_14257_),
    .A3(_14258_),
    .B1(_13292_),
    .X(_14698_));
 sky130_fd_sc_hd__xnor2_1 _41927_ (.A(_13846_),
    .B(_14698_),
    .Y(_14699_));
 sky130_fd_sc_hd__o31a_1 _41928_ (.A1(_12783_),
    .A2(_10947_),
    .A3(_10324_),
    .B1(_13850_),
    .X(_14700_));
 sky130_fd_sc_hd__xnor2_1 _41929_ (.A(_14699_),
    .B(_14700_),
    .Y(_14701_));
 sky130_fd_sc_hd__xor2_4 _41930_ (.A(_08967_),
    .B(_13833_),
    .X(_14703_));
 sky130_fd_sc_hd__nand2_2 _41931_ (.A(_13838_),
    .B(_13839_),
    .Y(_14704_));
 sky130_fd_sc_hd__a21oi_4 _41932_ (.A1(_09006_),
    .A2(_03031_),
    .B1(_04527_),
    .Y(_14705_));
 sky130_fd_sc_hd__nor2_2 _41933_ (.A(_07550_),
    .B(_07516_),
    .Y(_14706_));
 sky130_fd_sc_hd__and2_1 _41934_ (.A(_07550_),
    .B(_07516_),
    .X(_14707_));
 sky130_fd_sc_hd__or2_2 _41935_ (.A(_14706_),
    .B(_14707_),
    .X(_14708_));
 sky130_fd_sc_hd__xor2_4 _41936_ (.A(_14705_),
    .B(_14708_),
    .X(_14709_));
 sky130_fd_sc_hd__xor2_4 _41937_ (.A(_14704_),
    .B(_14709_),
    .X(_14710_));
 sky130_fd_sc_hd__xnor2_4 _41938_ (.A(_14703_),
    .B(_14710_),
    .Y(_14711_));
 sky130_fd_sc_hd__nand2_1 _41939_ (.A(_14701_),
    .B(_14711_),
    .Y(_14712_));
 sky130_fd_sc_hd__or2_1 _41940_ (.A(_14701_),
    .B(_14711_),
    .X(_14714_));
 sky130_fd_sc_hd__nand2_1 _41941_ (.A(_14712_),
    .B(_14714_),
    .Y(_14715_));
 sky130_fd_sc_hd__a21oi_1 _41942_ (.A1(_13307_),
    .A2(_14697_),
    .B1(_14715_),
    .Y(_14716_));
 sky130_fd_sc_hd__buf_1 _41943_ (.A(_14716_),
    .X(_14717_));
 sky130_fd_sc_hd__o21ai_2 _41944_ (.A1(_13853_),
    .A2(_13854_),
    .B1(_13858_),
    .Y(_14718_));
 sky130_fd_sc_hd__inv_2 _41945_ (.A(_14718_),
    .Y(_14719_));
 sky130_fd_sc_hd__a31o_1 _41946_ (.A1(_13307_),
    .A2(_14715_),
    .A3(_14697_),
    .B1(_14719_),
    .X(_14720_));
 sky130_fd_sc_hd__and3_1 _41947_ (.A(_13307_),
    .B(_14715_),
    .C(_14697_),
    .X(_14721_));
 sky130_fd_sc_hd__nor2_1 _41948_ (.A(_14716_),
    .B(_14721_),
    .Y(_14722_));
 sky130_fd_sc_hd__o22a_1 _41949_ (.A1(_14717_),
    .A2(_14720_),
    .B1(_14718_),
    .B2(_14722_),
    .X(_14723_));
 sky130_fd_sc_hd__nand2_1 _41950_ (.A(_14696_),
    .B(_14723_),
    .Y(_14725_));
 sky130_fd_sc_hd__a21boi_1 _41951_ (.A1(_13869_),
    .A2(_13826_),
    .B1_N(_13820_),
    .Y(_14726_));
 sky130_fd_sc_hd__o22ai_1 _41952_ (.A1(_14717_),
    .A2(_14720_),
    .B1(_14718_),
    .B2(_14722_),
    .Y(_14727_));
 sky130_fd_sc_hd__o211ai_1 _41953_ (.A1(_14684_),
    .A2(_14687_),
    .B1(_14695_),
    .C1(_14727_),
    .Y(_14728_));
 sky130_fd_sc_hd__nand3_2 _41954_ (.A(_14725_),
    .B(_14726_),
    .C(_14728_),
    .Y(_14729_));
 sky130_fd_sc_hd__a21bo_1 _41955_ (.A1(_13869_),
    .A2(_13827_),
    .B1_N(_13821_),
    .X(_14730_));
 sky130_fd_sc_hd__o221a_1 _41956_ (.A1(_13853_),
    .A2(_13854_),
    .B1(_14717_),
    .B2(_14721_),
    .C1(_13858_),
    .X(_14731_));
 sky130_fd_sc_hd__nor2_1 _41957_ (.A(_14717_),
    .B(_14720_),
    .Y(_14732_));
 sky130_fd_sc_hd__o21ai_1 _41958_ (.A1(_14731_),
    .A2(_14732_),
    .B1(_14696_),
    .Y(_14733_));
 sky130_fd_sc_hd__o211ai_2 _41959_ (.A1(_14684_),
    .A2(_14687_),
    .B1(_14695_),
    .C1(_14723_),
    .Y(_14734_));
 sky130_fd_sc_hd__nand3_2 _41960_ (.A(_14730_),
    .B(_14733_),
    .C(_14734_),
    .Y(_14736_));
 sky130_fd_sc_hd__nand2_1 _41961_ (.A(_13864_),
    .B(_13863_),
    .Y(_14737_));
 sky130_fd_sc_hd__a21oi_4 _41962_ (.A1(_13892_),
    .A2(_13876_),
    .B1(_13891_),
    .Y(_14738_));
 sky130_fd_sc_hd__inv_2 _41963_ (.A(_14738_),
    .Y(_14739_));
 sky130_fd_sc_hd__or2_1 _41964_ (.A(_01420_),
    .B(_04582_),
    .X(_14740_));
 sky130_fd_sc_hd__nor2_1 _41965_ (.A(_13879_),
    .B(_14740_),
    .Y(_14741_));
 sky130_fd_sc_hd__o21a_1 _41966_ (.A1(_01420_),
    .A2(_04582_),
    .B1(_13879_),
    .X(_14742_));
 sky130_fd_sc_hd__a211o_1 _41967_ (.A1(_25240_),
    .A2(_04473_),
    .B1(_14741_),
    .C1(_14742_),
    .X(_14743_));
 sky130_fd_sc_hd__o211ai_2 _41968_ (.A1(_14741_),
    .A2(_14742_),
    .B1(_07597_),
    .C1(_04572_),
    .Y(_14744_));
 sky130_fd_sc_hd__and4_1 _41969_ (.A(_14743_),
    .B(_14744_),
    .C(_08966_),
    .D(_12762_),
    .X(_14745_));
 sky130_fd_sc_hd__a22oi_1 _41970_ (.A1(_10296_),
    .A2(_12762_),
    .B1(_14743_),
    .B2(_14744_),
    .Y(_14747_));
 sky130_fd_sc_hd__nor2_1 _41971_ (.A(_14745_),
    .B(_14747_),
    .Y(_14748_));
 sky130_fd_sc_hd__xnor2_1 _41972_ (.A(_13881_),
    .B(_14748_),
    .Y(_14749_));
 sky130_fd_sc_hd__nand3_1 _41973_ (.A(_13842_),
    .B(_13857_),
    .C(_14749_),
    .Y(_14750_));
 sky130_fd_sc_hd__a21o_1 _41974_ (.A1(_13842_),
    .A2(_13857_),
    .B1(_14749_),
    .X(_14751_));
 sky130_fd_sc_hd__nand2_1 _41975_ (.A(_14750_),
    .B(_14751_),
    .Y(_14752_));
 sky130_fd_sc_hd__a21o_1 _41976_ (.A1(_13884_),
    .A2(_13886_),
    .B1(_14752_),
    .X(_14753_));
 sky130_fd_sc_hd__nand3_1 _41977_ (.A(_13884_),
    .B(_13886_),
    .C(_14752_),
    .Y(_14754_));
 sky130_fd_sc_hd__and2_2 _41978_ (.A(_14753_),
    .B(_14754_),
    .X(_14755_));
 sky130_fd_sc_hd__and2_1 _41979_ (.A(_14739_),
    .B(_14755_),
    .X(_14756_));
 sky130_fd_sc_hd__nor2_1 _41980_ (.A(_14755_),
    .B(_14739_),
    .Y(_14758_));
 sky130_fd_sc_hd__or2_1 _41981_ (.A(_14756_),
    .B(_14758_),
    .X(_14759_));
 sky130_fd_sc_hd__a21o_1 _41982_ (.A1(_13861_),
    .A2(_14737_),
    .B1(_14759_),
    .X(_14760_));
 sky130_fd_sc_hd__nand3_2 _41983_ (.A(_13861_),
    .B(_14737_),
    .C(_14759_),
    .Y(_14761_));
 sky130_fd_sc_hd__a21oi_1 _41984_ (.A1(_14760_),
    .A2(_14761_),
    .B1(_13895_),
    .Y(_14762_));
 sky130_fd_sc_hd__nand3_1 _41985_ (.A(_14760_),
    .B(_14761_),
    .C(_13895_),
    .Y(_14763_));
 sky130_fd_sc_hd__and2b_1 _41986_ (.A_N(_14762_),
    .B(_14763_),
    .X(_14764_));
 sky130_fd_sc_hd__a21oi_2 _41987_ (.A1(_14729_),
    .A2(_14736_),
    .B1(_14764_),
    .Y(_14765_));
 sky130_fd_sc_hd__and3_1 _41988_ (.A(_14729_),
    .B(_14736_),
    .C(_14764_),
    .X(_14766_));
 sky130_fd_sc_hd__nand2_1 _41989_ (.A(_13821_),
    .B(_13827_),
    .Y(_14767_));
 sky130_fd_sc_hd__a22oi_1 _41990_ (.A1(_12810_),
    .A2(_12805_),
    .B1(_13872_),
    .B2(_14767_),
    .Y(_14769_));
 sky130_fd_sc_hd__a22o_1 _41991_ (.A1(_13868_),
    .A2(_14769_),
    .B1(_13875_),
    .B2(_13903_),
    .X(_14770_));
 sky130_fd_sc_hd__o21bai_2 _41992_ (.A1(_14765_),
    .A2(_14766_),
    .B1_N(_14770_),
    .Y(_14771_));
 sky130_fd_sc_hd__a21o_1 _41993_ (.A1(_14729_),
    .A2(_14736_),
    .B1(_14764_),
    .X(_14772_));
 sky130_fd_sc_hd__nand3_1 _41994_ (.A(_14729_),
    .B(_14736_),
    .C(_14764_),
    .Y(_14773_));
 sky130_fd_sc_hd__nand3_1 _41995_ (.A(_14770_),
    .B(_14772_),
    .C(_14773_),
    .Y(_14774_));
 sky130_fd_sc_hd__a21oi_2 _41996_ (.A1(_12838_),
    .A2(_13901_),
    .B1(_13898_),
    .Y(_14775_));
 sky130_fd_sc_hd__a21oi_1 _41997_ (.A1(_14771_),
    .A2(_14774_),
    .B1(_14775_),
    .Y(_14776_));
 sky130_fd_sc_hd__nand2_1 _41998_ (.A(_14770_),
    .B(_14773_),
    .Y(_14777_));
 sky130_fd_sc_hd__o211a_1 _41999_ (.A1(_14765_),
    .A2(_14777_),
    .B1(_14775_),
    .C1(_14771_),
    .X(_14778_));
 sky130_fd_sc_hd__a32oi_4 _42000_ (.A1(_13905_),
    .A2(_13906_),
    .A3(_13904_),
    .B1(_13912_),
    .B2(_13913_),
    .Y(_14780_));
 sky130_fd_sc_hd__o21ai_1 _42001_ (.A1(_14776_),
    .A2(_14778_),
    .B1(_14780_),
    .Y(_14781_));
 sky130_fd_sc_hd__a21oi_1 _42002_ (.A1(_14772_),
    .A2(_14773_),
    .B1(_14770_),
    .Y(_14782_));
 sky130_fd_sc_hd__nor2_1 _42003_ (.A(_14765_),
    .B(_14777_),
    .Y(_14783_));
 sky130_fd_sc_hd__o21bai_1 _42004_ (.A1(_14782_),
    .A2(_14783_),
    .B1_N(_14775_),
    .Y(_14784_));
 sky130_fd_sc_hd__o211ai_1 _42005_ (.A1(_14765_),
    .A2(_14777_),
    .B1(_14775_),
    .C1(_14771_),
    .Y(_14785_));
 sky130_fd_sc_hd__nand3b_1 _42006_ (.A_N(_14780_),
    .B(_14784_),
    .C(_14785_),
    .Y(_14786_));
 sky130_fd_sc_hd__nand2_2 _42007_ (.A(_14781_),
    .B(_14786_),
    .Y(_14787_));
 sky130_fd_sc_hd__a21bo_1 _42008_ (.A1(_13917_),
    .A2(_13925_),
    .B1_N(_13918_),
    .X(_14788_));
 sky130_fd_sc_hd__xnor2_4 _42009_ (.A(_14787_),
    .B(_14788_),
    .Y(_00015_));
 sky130_fd_sc_hd__a31oi_2 _42010_ (.A1(_13307_),
    .A2(_14715_),
    .A3(_14697_),
    .B1(_14719_),
    .Y(_14790_));
 sky130_fd_sc_hd__a21o_2 _42011_ (.A1(_13881_),
    .A2(_14748_),
    .B1(_14745_),
    .X(_14791_));
 sky130_fd_sc_hd__and2_1 _42012_ (.A(_14704_),
    .B(_14709_),
    .X(_14792_));
 sky130_fd_sc_hd__a21oi_1 _42013_ (.A1(_14703_),
    .A2(_14710_),
    .B1(_14792_),
    .Y(_14793_));
 sky130_fd_sc_hd__o211a_1 _42014_ (.A1(_14741_),
    .A2(_14742_),
    .B1(_07597_),
    .C1(_04572_),
    .X(_14794_));
 sky130_fd_sc_hd__a31o_1 _42015_ (.A1(_10467_),
    .A2(_25256_),
    .A3(_14740_),
    .B1(_14794_),
    .X(_14795_));
 sky130_fd_sc_hd__clkbuf_2 _42016_ (.A(_03003_),
    .X(_14796_));
 sky130_fd_sc_hd__o221a_1 _42017_ (.A1(_01420_),
    .A2(_04582_),
    .B1(_03002_),
    .B2(_14796_),
    .C1(_07507_),
    .X(_14797_));
 sky130_fd_sc_hd__a21oi_1 _42018_ (.A1(_14740_),
    .A2(_07507_),
    .B1(_03005_),
    .Y(_14798_));
 sky130_fd_sc_hd__a211oi_1 _42019_ (.A1(_04572_),
    .A2(_04575_),
    .B1(_14797_),
    .C1(_14798_),
    .Y(_14799_));
 sky130_fd_sc_hd__o211a_1 _42020_ (.A1(_14797_),
    .A2(_14798_),
    .B1(_04473_),
    .C1(_04575_),
    .X(_14801_));
 sky130_fd_sc_hd__and4bb_1 _42021_ (.A_N(_14799_),
    .B_N(_14801_),
    .C(_08966_),
    .D(_13833_),
    .X(_14802_));
 sky130_fd_sc_hd__o2bb2a_1 _42022_ (.A1_N(_08966_),
    .A2_N(_13833_),
    .B1(_14799_),
    .B2(_14801_),
    .X(_14803_));
 sky130_fd_sc_hd__nor2_1 _42023_ (.A(_14802_),
    .B(_14803_),
    .Y(_14804_));
 sky130_fd_sc_hd__xnor2_1 _42024_ (.A(_14795_),
    .B(_14804_),
    .Y(_14805_));
 sky130_fd_sc_hd__and2_1 _42025_ (.A(_14793_),
    .B(_14805_),
    .X(_14806_));
 sky130_fd_sc_hd__nor2_1 _42026_ (.A(_14805_),
    .B(_14793_),
    .Y(_14807_));
 sky130_fd_sc_hd__nor2_2 _42027_ (.A(_14806_),
    .B(_14807_),
    .Y(_14808_));
 sky130_fd_sc_hd__xnor2_2 _42028_ (.A(_14791_),
    .B(_14808_),
    .Y(_14809_));
 sky130_fd_sc_hd__and3_1 _42029_ (.A(_14751_),
    .B(_14753_),
    .C(_14809_),
    .X(_14810_));
 sky130_fd_sc_hd__a21oi_4 _42030_ (.A1(_14751_),
    .A2(_14753_),
    .B1(_14809_),
    .Y(_14812_));
 sky130_fd_sc_hd__or2_2 _42031_ (.A(_14810_),
    .B(_14812_),
    .X(_14813_));
 sky130_fd_sc_hd__inv_2 _42032_ (.A(_14813_),
    .Y(_14814_));
 sky130_fd_sc_hd__o21a_1 _42033_ (.A1(_14716_),
    .A2(_14790_),
    .B1(_14814_),
    .X(_14815_));
 sky130_fd_sc_hd__a21oi_2 _42034_ (.A1(_14755_),
    .A2(_14739_),
    .B1(_14815_),
    .Y(_14816_));
 sky130_fd_sc_hd__o31a_1 _42035_ (.A1(_14717_),
    .A2(_14790_),
    .A3(_14814_),
    .B1(_14816_),
    .X(_14817_));
 sky130_fd_sc_hd__nand3b_2 _42036_ (.A_N(_14716_),
    .B(_14720_),
    .C(_14813_),
    .Y(_14818_));
 sky130_fd_sc_hd__inv_2 _42037_ (.A(_14818_),
    .Y(_14819_));
 sky130_fd_sc_hd__o211a_1 _42038_ (.A1(_14819_),
    .A2(_14815_),
    .B1(_14755_),
    .C1(_14739_),
    .X(_14820_));
 sky130_fd_sc_hd__a31oi_1 _42039_ (.A1(_14254_),
    .A2(_14269_),
    .A3(_14682_),
    .B1(_14681_),
    .Y(_14821_));
 sky130_fd_sc_hd__and2b_1 _42040_ (.A_N(_14527_),
    .B(_14545_),
    .X(_14823_));
 sky130_fd_sc_hd__o21ai_1 _42041_ (.A1(_11524_),
    .A2(_12633_),
    .B1(_09582_),
    .Y(_14824_));
 sky130_fd_sc_hd__xnor2_1 _42042_ (.A(_12640_),
    .B(_14824_),
    .Y(_14825_));
 sky130_fd_sc_hd__xnor2_2 _42043_ (.A(_14622_),
    .B(_14825_),
    .Y(_14826_));
 sky130_fd_sc_hd__a21oi_1 _42044_ (.A1(_14627_),
    .A2(_14630_),
    .B1(_14826_),
    .Y(_14827_));
 sky130_fd_sc_hd__and3_1 _42045_ (.A(_14627_),
    .B(_14630_),
    .C(_14826_),
    .X(_14828_));
 sky130_fd_sc_hd__o211ai_1 _42046_ (.A1(_13736_),
    .A2(_13737_),
    .B1(_13751_),
    .C1(_14639_),
    .Y(_14829_));
 sky130_fd_sc_hd__o21ai_2 _42047_ (.A1(_13738_),
    .A2(_13739_),
    .B1(_13740_),
    .Y(_14830_));
 sky130_fd_sc_hd__o211a_1 _42048_ (.A1(_13738_),
    .A2(_13739_),
    .B1(_13740_),
    .C1(_09610_),
    .X(_14831_));
 sky130_fd_sc_hd__a21o_1 _42049_ (.A1(_12664_),
    .A2(_14830_),
    .B1(_14831_),
    .X(_14832_));
 sky130_fd_sc_hd__xor2_1 _42050_ (.A(_14638_),
    .B(_14832_),
    .X(_14834_));
 sky130_fd_sc_hd__a21oi_1 _42051_ (.A1(_14829_),
    .A2(_14642_),
    .B1(_14834_),
    .Y(_14835_));
 sky130_fd_sc_hd__and3_1 _42052_ (.A(_14829_),
    .B(_14642_),
    .C(_14834_),
    .X(_14836_));
 sky130_fd_sc_hd__nor2_1 _42053_ (.A(_14835_),
    .B(_14836_),
    .Y(_14837_));
 sky130_fd_sc_hd__o21bai_1 _42054_ (.A1(_14827_),
    .A2(_14828_),
    .B1_N(_14837_),
    .Y(_14838_));
 sky130_fd_sc_hd__a21o_1 _42055_ (.A1(_14627_),
    .A2(_14630_),
    .B1(_14826_),
    .X(_14839_));
 sky130_fd_sc_hd__nand3b_1 _42056_ (.A_N(_14828_),
    .B(_14837_),
    .C(_14839_),
    .Y(_14840_));
 sky130_fd_sc_hd__nand2_1 _42057_ (.A(_11476_),
    .B(_08289_),
    .Y(_14841_));
 sky130_fd_sc_hd__a22oi_4 _42058_ (.A1(_14841_),
    .A2(_08295_),
    .B1(_13767_),
    .B2(_14652_),
    .Y(_14842_));
 sky130_fd_sc_hd__a21oi_1 _42059_ (.A1(_14838_),
    .A2(_14840_),
    .B1(_14842_),
    .Y(_14843_));
 sky130_fd_sc_hd__nand3_1 _42060_ (.A(_14840_),
    .B(_14842_),
    .C(_14838_),
    .Y(_14845_));
 sky130_fd_sc_hd__inv_2 _42061_ (.A(_14845_),
    .Y(_14846_));
 sky130_fd_sc_hd__nor4_1 _42062_ (.A(_14543_),
    .B(_14823_),
    .C(_14843_),
    .D(_14846_),
    .Y(_14847_));
 sky130_fd_sc_hd__o22a_1 _42063_ (.A1(_14543_),
    .A2(_14823_),
    .B1(_14843_),
    .B2(_14846_),
    .X(_14848_));
 sky130_fd_sc_hd__a211oi_1 _42064_ (.A1(_14656_),
    .A2(_14664_),
    .B1(_14847_),
    .C1(_14848_),
    .Y(_14849_));
 sky130_fd_sc_hd__o211a_1 _42065_ (.A1(_14847_),
    .A2(_14848_),
    .B1(_14656_),
    .C1(_14664_),
    .X(_14850_));
 sky130_fd_sc_hd__nor2_2 _42066_ (.A(_14849_),
    .B(_14850_),
    .Y(_14851_));
 sky130_fd_sc_hd__inv_2 _42067_ (.A(_14661_),
    .Y(_14852_));
 sky130_fd_sc_hd__a2bb2o_2 _42068_ (.A1_N(_14619_),
    .A2_N(_14852_),
    .B1(_14663_),
    .B2(_14664_),
    .X(_14853_));
 sky130_fd_sc_hd__nand2_1 _42069_ (.A(_14851_),
    .B(_14853_),
    .Y(_14854_));
 sky130_fd_sc_hd__or2_1 _42070_ (.A(_14853_),
    .B(_14851_),
    .X(_14856_));
 sky130_fd_sc_hd__clkbuf_2 _42071_ (.A(_11583_),
    .X(_14857_));
 sky130_fd_sc_hd__a2111oi_1 _42072_ (.A1(_11568_),
    .A2(_14606_),
    .B1(_13791_),
    .C1(_14605_),
    .D1(_14857_),
    .Y(_14858_));
 sky130_fd_sc_hd__a21oi_2 _42073_ (.A1(_14857_),
    .A2(_14609_),
    .B1(net88),
    .Y(_14859_));
 sky130_fd_sc_hd__xor2_4 _42074_ (.A(_13803_),
    .B(_14859_),
    .X(_14860_));
 sky130_fd_sc_hd__clkbuf_2 _42075_ (.A(_14860_),
    .X(_14861_));
 sky130_fd_sc_hd__and3_1 _42076_ (.A(_14854_),
    .B(_14856_),
    .C(_14861_),
    .X(_14862_));
 sky130_fd_sc_hd__a21oi_1 _42077_ (.A1(_14854_),
    .A2(_14856_),
    .B1(_14861_),
    .Y(_14863_));
 sky130_fd_sc_hd__a21o_1 _42078_ (.A1(_14597_),
    .A2(_14507_),
    .B1(_14595_),
    .X(_14864_));
 sky130_fd_sc_hd__o21a_2 _42079_ (.A1(_14862_),
    .A2(_14863_),
    .B1(_14864_),
    .X(_14865_));
 sky130_fd_sc_hd__nor3_1 _42080_ (.A(_14863_),
    .B(_14864_),
    .C(_14862_),
    .Y(_14867_));
 sky130_fd_sc_hd__nand3_4 _42081_ (.A(_14618_),
    .B(_14666_),
    .C(_14667_),
    .Y(_14868_));
 sky130_fd_sc_hd__a21oi_1 _42082_ (.A1(_14617_),
    .A2(_14868_),
    .B1(_14670_),
    .Y(_14869_));
 sky130_fd_sc_hd__o21ba_1 _42083_ (.A1(_14865_),
    .A2(_14867_),
    .B1_N(_14869_),
    .X(_14870_));
 sky130_fd_sc_hd__a2111oi_1 _42084_ (.A1(_14617_),
    .A2(_14868_),
    .B1(_14670_),
    .C1(_14865_),
    .D1(_14867_),
    .Y(_14871_));
 sky130_fd_sc_hd__a21oi_1 _42085_ (.A1(_14577_),
    .A2(_14579_),
    .B1(_14575_),
    .Y(_14872_));
 sky130_fd_sc_hd__nand2_1 _42086_ (.A(_14567_),
    .B(_14563_),
    .Y(_14873_));
 sky130_fd_sc_hd__or3_1 _42087_ (.A(_05529_),
    .B(_07015_),
    .C(_11336_),
    .X(_14874_));
 sky130_fd_sc_hd__nor2_1 _42088_ (.A(_07013_),
    .B(_11349_),
    .Y(_14875_));
 sky130_fd_sc_hd__and2_1 _42089_ (.A(_07013_),
    .B(_08802_),
    .X(_14876_));
 sky130_fd_sc_hd__a211oi_2 _42090_ (.A1(_14564_),
    .A2(_14874_),
    .B1(_14875_),
    .C1(_14876_),
    .Y(_14878_));
 sky130_fd_sc_hd__o221a_1 _42091_ (.A1(_14875_),
    .A2(_14876_),
    .B1(_05529_),
    .B2(_13340_),
    .C1(_14874_),
    .X(_14879_));
 sky130_fd_sc_hd__or4bb_1 _42092_ (.A(_14878_),
    .B(_14879_),
    .C_N(_13343_),
    .D_N(_14567_),
    .X(_14880_));
 sky130_fd_sc_hd__a2bb2o_1 _42093_ (.A1_N(_14878_),
    .A2_N(_14879_),
    .B1(_13343_),
    .B2(_14567_),
    .X(_14881_));
 sky130_fd_sc_hd__and3_1 _42094_ (.A(_14880_),
    .B(_14881_),
    .C(_13336_),
    .X(_14882_));
 sky130_fd_sc_hd__a21oi_1 _42095_ (.A1(_14880_),
    .A2(_14881_),
    .B1(_13336_),
    .Y(_14883_));
 sky130_fd_sc_hd__a211o_1 _42096_ (.A1(_14571_),
    .A2(_14873_),
    .B1(_14882_),
    .C1(_14883_),
    .X(_14884_));
 sky130_fd_sc_hd__o211ai_1 _42097_ (.A1(_14882_),
    .A2(_14883_),
    .B1(_14571_),
    .C1(_14873_),
    .Y(_14885_));
 sky130_fd_sc_hd__and3_1 _42098_ (.A(_14872_),
    .B(_14884_),
    .C(_14885_),
    .X(_14886_));
 sky130_fd_sc_hd__a21oi_1 _42099_ (.A1(_14885_),
    .A2(_14884_),
    .B1(_14872_),
    .Y(_14887_));
 sky130_fd_sc_hd__or2_1 _42100_ (.A(_14886_),
    .B(_14887_),
    .X(_14889_));
 sky130_fd_sc_hd__o31ai_1 _42101_ (.A1(_13325_),
    .A2(_13331_),
    .A3(_13330_),
    .B1(_14557_),
    .Y(_14890_));
 sky130_fd_sc_hd__and2_1 _42102_ (.A(_07039_),
    .B(_13318_),
    .X(_14891_));
 sky130_fd_sc_hd__a2bb2o_1 _42103_ (.A1_N(_05498_),
    .A2_N(_05495_),
    .B1(_00971_),
    .B2(_05508_),
    .X(_14892_));
 sky130_fd_sc_hd__o21a_1 _42104_ (.A1(_05497_),
    .A2(_14891_),
    .B1(_14892_),
    .X(_14893_));
 sky130_fd_sc_hd__xnor2_1 _42105_ (.A(_08828_),
    .B(_14891_),
    .Y(_14894_));
 sky130_fd_sc_hd__xnor2_1 _42106_ (.A(_14893_),
    .B(_14894_),
    .Y(_14895_));
 sky130_fd_sc_hd__xor2_1 _42107_ (.A(_14556_),
    .B(_14895_),
    .X(_14896_));
 sky130_fd_sc_hd__and2_1 _42108_ (.A(_14890_),
    .B(_14896_),
    .X(_14897_));
 sky130_fd_sc_hd__nor2_1 _42109_ (.A(_14896_),
    .B(_14890_),
    .Y(_14898_));
 sky130_fd_sc_hd__or3_1 _42110_ (.A(_14889_),
    .B(_14897_),
    .C(_14898_),
    .X(_14900_));
 sky130_fd_sc_hd__o21ai_1 _42111_ (.A1(_14897_),
    .A2(_14898_),
    .B1(_14889_),
    .Y(_14901_));
 sky130_fd_sc_hd__and3_1 _42112_ (.A(_14900_),
    .B(_13310_),
    .C(_14901_),
    .X(_14902_));
 sky130_fd_sc_hd__buf_1 _42113_ (.A(_13310_),
    .X(_14903_));
 sky130_fd_sc_hd__a21oi_1 _42114_ (.A1(_14901_),
    .A2(_14900_),
    .B1(_14903_),
    .Y(_14904_));
 sky130_fd_sc_hd__a21oi_1 _42115_ (.A1(_14586_),
    .A2(_14584_),
    .B1(_14582_),
    .Y(_14905_));
 sky130_fd_sc_hd__o21a_1 _42116_ (.A1(_14902_),
    .A2(_14904_),
    .B1(_14905_),
    .X(_14906_));
 sky130_fd_sc_hd__nor3_1 _42117_ (.A(_14905_),
    .B(_14902_),
    .C(_14904_),
    .Y(_14907_));
 sky130_fd_sc_hd__or2_1 _42118_ (.A(_14906_),
    .B(_14907_),
    .X(_14908_));
 sky130_fd_sc_hd__o211a_1 _42119_ (.A1(net164),
    .A2(_12528_),
    .B1(_13403_),
    .C1(_14535_),
    .X(_14909_));
 sky130_fd_sc_hd__inv_2 _42120_ (.A(_14909_),
    .Y(_14911_));
 sky130_fd_sc_hd__a21oi_1 _42121_ (.A1(_10204_),
    .A2(_11423_),
    .B1(_12516_),
    .Y(_14912_));
 sky130_fd_sc_hd__o31a_1 _42122_ (.A1(_11413_),
    .A2(_12513_),
    .A3(_11414_),
    .B1(_11423_),
    .X(_14913_));
 sky130_fd_sc_hd__a22o_1 _42123_ (.A1(_14529_),
    .A2(_14912_),
    .B1(_14531_),
    .B2(_14913_),
    .X(_14914_));
 sky130_fd_sc_hd__xnor2_1 _42124_ (.A(_14534_),
    .B(_14914_),
    .Y(_14915_));
 sky130_fd_sc_hd__a21oi_2 _42125_ (.A1(_14911_),
    .A2(_14539_),
    .B1(_14915_),
    .Y(_14916_));
 sky130_fd_sc_hd__and3_1 _42126_ (.A(_14911_),
    .B(_14539_),
    .C(_14915_),
    .X(_14917_));
 sky130_fd_sc_hd__o21ai_4 _42127_ (.A1(_14916_),
    .A2(_14917_),
    .B1(_14544_),
    .Y(_14918_));
 sky130_fd_sc_hd__or3_4 _42128_ (.A(_14544_),
    .B(_14916_),
    .C(_14917_),
    .X(_14919_));
 sky130_fd_sc_hd__nor2_1 _42129_ (.A(_10245_),
    .B(_14512_),
    .Y(_14920_));
 sky130_fd_sc_hd__and2_1 _42130_ (.A(_10245_),
    .B(_14512_),
    .X(_14922_));
 sky130_fd_sc_hd__o22ai_2 _42131_ (.A1(_14508_),
    .A2(_14511_),
    .B1(_14920_),
    .B2(_14922_),
    .Y(_14923_));
 sky130_fd_sc_hd__or4_1 _42132_ (.A(_14508_),
    .B(_14511_),
    .C(_14920_),
    .D(_14922_),
    .X(_14924_));
 sky130_fd_sc_hd__and3_1 _42133_ (.A(_14518_),
    .B(_14923_),
    .C(_14924_),
    .X(_14925_));
 sky130_fd_sc_hd__a21oi_1 _42134_ (.A1(_14923_),
    .A2(_14924_),
    .B1(_14518_),
    .Y(_14926_));
 sky130_fd_sc_hd__nor2_1 _42135_ (.A(_14925_),
    .B(_14926_),
    .Y(_14927_));
 sky130_fd_sc_hd__o21a_1 _42136_ (.A1(_14525_),
    .A2(_14522_),
    .B1(_14927_),
    .X(_14928_));
 sky130_fd_sc_hd__nor3_1 _42137_ (.A(_14525_),
    .B(_14522_),
    .C(_14927_),
    .Y(_14929_));
 sky130_fd_sc_hd__nor2_1 _42138_ (.A(_14928_),
    .B(_14929_),
    .Y(_14930_));
 sky130_fd_sc_hd__nand2_2 _42139_ (.A(_14930_),
    .B(_14918_),
    .Y(_14931_));
 sky130_fd_sc_hd__a21boi_1 _42140_ (.A1(_14918_),
    .A2(_14919_),
    .B1_N(_14930_),
    .Y(_14933_));
 sky130_fd_sc_hd__a31oi_4 _42141_ (.A1(_14918_),
    .A2(_14919_),
    .A3(_14931_),
    .B1(_14933_),
    .Y(_14934_));
 sky130_fd_sc_hd__xnor2_2 _42142_ (.A(_14908_),
    .B(_14934_),
    .Y(_14935_));
 sky130_fd_sc_hd__o211ai_2 _42143_ (.A1(_14344_),
    .A2(_14346_),
    .B1(_14343_),
    .C1(_14935_),
    .Y(_14936_));
 sky130_fd_sc_hd__a21o_1 _42144_ (.A1(_14343_),
    .A2(_14348_),
    .B1(_14935_),
    .X(_14937_));
 sky130_fd_sc_hd__nand2_1 _42145_ (.A(_14590_),
    .B(_14594_),
    .Y(_14938_));
 sky130_fd_sc_hd__a21o_1 _42146_ (.A1(_14936_),
    .A2(_14937_),
    .B1(_14938_),
    .X(_14939_));
 sky130_fd_sc_hd__nand3_1 _42147_ (.A(_14938_),
    .B(_14936_),
    .C(_14937_),
    .Y(_14940_));
 sky130_fd_sc_hd__nand2_1 _42148_ (.A(_14939_),
    .B(_14940_),
    .Y(_14941_));
 sky130_fd_sc_hd__inv_2 _42149_ (.A(_14382_),
    .Y(_14942_));
 sky130_fd_sc_hd__o21ai_4 _42150_ (.A1(_14404_),
    .A2(_14942_),
    .B1(_14384_),
    .Y(_14944_));
 sky130_fd_sc_hd__buf_1 _42151_ (.A(_08598_),
    .X(_14945_));
 sky130_fd_sc_hd__or3b_1 _42152_ (.A(_07255_),
    .B(_12324_),
    .C_N(_14945_),
    .X(_14946_));
 sky130_fd_sc_hd__buf_1 _42153_ (.A(_13519_),
    .X(_14947_));
 sky130_fd_sc_hd__a21bo_1 _42154_ (.A1(_14946_),
    .A2(_13521_),
    .B1_N(_14947_),
    .X(_14948_));
 sky130_fd_sc_hd__nor2_1 _42155_ (.A(_14945_),
    .B(_14353_),
    .Y(_14949_));
 sky130_fd_sc_hd__a211o_1 _42156_ (.A1(_12324_),
    .A2(_14949_),
    .B1(_14947_),
    .C1(_12327_),
    .X(_14950_));
 sky130_fd_sc_hd__o311a_1 _42157_ (.A1(_13521_),
    .A2(_14945_),
    .A3(_14353_),
    .B1(_14948_),
    .C1(_14950_),
    .X(_14951_));
 sky130_fd_sc_hd__a21boi_1 _42158_ (.A1(_14357_),
    .A2(_13530_),
    .B1_N(_14358_),
    .Y(_14952_));
 sky130_fd_sc_hd__xnor2_1 _42159_ (.A(_14951_),
    .B(_14952_),
    .Y(_14953_));
 sky130_fd_sc_hd__a21o_1 _42160_ (.A1(_14363_),
    .A2(_14365_),
    .B1(_14953_),
    .X(_14955_));
 sky130_fd_sc_hd__nand3_2 _42161_ (.A(_14363_),
    .B(_14365_),
    .C(_14953_),
    .Y(_14956_));
 sky130_fd_sc_hd__nor2_1 _42162_ (.A(_14375_),
    .B(_14376_),
    .Y(_14957_));
 sky130_fd_sc_hd__buf_2 _42163_ (.A(_13545_),
    .X(_14958_));
 sky130_fd_sc_hd__xnor2_2 _42164_ (.A(_14958_),
    .B(_13552_),
    .Y(_14959_));
 sky130_fd_sc_hd__a41oi_4 _42165_ (.A1(_11158_),
    .A2(_14368_),
    .A3(_14958_),
    .A4(_14369_),
    .B1(_14373_),
    .Y(_14960_));
 sky130_fd_sc_hd__xor2_2 _42166_ (.A(_14959_),
    .B(_14960_),
    .X(_14961_));
 sky130_fd_sc_hd__o21a_1 _42167_ (.A1(_14957_),
    .A2(_14379_),
    .B1(_14961_),
    .X(_14962_));
 sky130_fd_sc_hd__nor3_1 _42168_ (.A(_14957_),
    .B(_14379_),
    .C(_14961_),
    .Y(_14963_));
 sky130_fd_sc_hd__nor2_2 _42169_ (.A(_14962_),
    .B(_14963_),
    .Y(_14964_));
 sky130_fd_sc_hd__a21o_1 _42170_ (.A1(_14955_),
    .A2(_14956_),
    .B1(_14964_),
    .X(_14966_));
 sky130_fd_sc_hd__nand3_4 _42171_ (.A(_14964_),
    .B(_14955_),
    .C(_14956_),
    .Y(_14967_));
 sky130_fd_sc_hd__o21ai_2 _42172_ (.A1(_14403_),
    .A2(_14385_),
    .B1(_14401_),
    .Y(_14968_));
 sky130_fd_sc_hd__o211a_1 _42173_ (.A1(_13568_),
    .A2(_11110_),
    .B1(_14387_),
    .C1(_13567_),
    .X(_14969_));
 sky130_fd_sc_hd__clkbuf_2 _42174_ (.A(_13567_),
    .X(_14970_));
 sky130_fd_sc_hd__o32a_1 _42175_ (.A1(_14970_),
    .A2(_14392_),
    .A3(_14386_),
    .B1(_14969_),
    .B2(_14389_),
    .X(_14971_));
 sky130_fd_sc_hd__o21ai_1 _42176_ (.A1(_13573_),
    .A2(_14392_),
    .B1(_14391_),
    .Y(_14972_));
 sky130_fd_sc_hd__o21ai_1 _42177_ (.A1(_14392_),
    .A2(_14386_),
    .B1(_13573_),
    .Y(_14973_));
 sky130_fd_sc_hd__a21boi_1 _42178_ (.A1(_14391_),
    .A2(_14972_),
    .B1_N(_14973_),
    .Y(_14974_));
 sky130_fd_sc_hd__nor2_1 _42179_ (.A(_14971_),
    .B(_14974_),
    .Y(_14975_));
 sky130_fd_sc_hd__nand2_1 _42180_ (.A(_14971_),
    .B(_14974_),
    .Y(_14977_));
 sky130_fd_sc_hd__or2b_1 _42181_ (.A(_14975_),
    .B_N(_14977_),
    .X(_14978_));
 sky130_fd_sc_hd__xor2_1 _42182_ (.A(_14969_),
    .B(_14978_),
    .X(_14979_));
 sky130_fd_sc_hd__and2b_1 _42183_ (.A_N(_14979_),
    .B(_14398_),
    .X(_14980_));
 sky130_fd_sc_hd__and2b_1 _42184_ (.A_N(_14398_),
    .B(_14979_),
    .X(_14981_));
 sky130_fd_sc_hd__nor2_1 _42185_ (.A(_14980_),
    .B(_14981_),
    .Y(_14982_));
 sky130_fd_sc_hd__xor2_2 _42186_ (.A(_14968_),
    .B(_14982_),
    .X(_14983_));
 sky130_fd_sc_hd__a21o_1 _42187_ (.A1(_14966_),
    .A2(_14967_),
    .B1(_14983_),
    .X(_14984_));
 sky130_fd_sc_hd__nand3_1 _42188_ (.A(_14966_),
    .B(_14967_),
    .C(_14983_),
    .Y(_14985_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _42189_ (.A(_14985_),
    .X(_14986_));
 sky130_fd_sc_hd__or2b_1 _42190_ (.A(_14410_),
    .B_N(_14429_),
    .X(_14988_));
 sky130_fd_sc_hd__nand3b_1 _42191_ (.A_N(_13656_),
    .B(_14433_),
    .C(_14430_),
    .Y(_14989_));
 sky130_fd_sc_hd__a211o_1 _42192_ (.A1(_04043_),
    .A2(_05697_),
    .B1(_12188_),
    .C1(_14428_),
    .X(_14990_));
 sky130_fd_sc_hd__a211oi_1 _42193_ (.A1(_13633_),
    .A2(_13643_),
    .B1(_14415_),
    .C1(_14417_),
    .Y(_14991_));
 sky130_fd_sc_hd__o22a_1 _42194_ (.A1(_13646_),
    .A2(_12182_),
    .B1(_07419_),
    .B2(_07420_),
    .X(_14992_));
 sky130_fd_sc_hd__or3_1 _42195_ (.A(_04047_),
    .B(_13634_),
    .C(_14992_),
    .X(_14993_));
 sky130_fd_sc_hd__nand4_2 _42196_ (.A(_14413_),
    .B(_14414_),
    .C(_13632_),
    .D(_12179_),
    .Y(_14994_));
 sky130_fd_sc_hd__o21a_1 _42197_ (.A1(_12181_),
    .A2(_07419_),
    .B1(_09798_),
    .X(_14995_));
 sky130_fd_sc_hd__xor2_1 _42198_ (.A(_14994_),
    .B(_14995_),
    .X(_14996_));
 sky130_fd_sc_hd__xnor2_1 _42199_ (.A(_14993_),
    .B(_14996_),
    .Y(_14997_));
 sky130_fd_sc_hd__or3_1 _42200_ (.A(_14991_),
    .B(_14997_),
    .C(_14423_),
    .X(_14999_));
 sky130_fd_sc_hd__o21ai_2 _42201_ (.A1(_14991_),
    .A2(_14423_),
    .B1(_14997_),
    .Y(_15000_));
 sky130_fd_sc_hd__o221a_1 _42202_ (.A1(_12199_),
    .A2(_12181_),
    .B1(_13634_),
    .B2(_05688_),
    .C1(_13646_),
    .X(_15001_));
 sky130_fd_sc_hd__and3_1 _42203_ (.A(_14999_),
    .B(_15000_),
    .C(_15001_),
    .X(_15002_));
 sky130_fd_sc_hd__a21oi_2 _42204_ (.A1(_14999_),
    .A2(_15000_),
    .B1(_15001_),
    .Y(_15003_));
 sky130_fd_sc_hd__a211o_1 _42205_ (.A1(_14424_),
    .A2(_14990_),
    .B1(_15002_),
    .C1(_15003_),
    .X(_15004_));
 sky130_fd_sc_hd__o221ai_4 _42206_ (.A1(_14411_),
    .A2(_14428_),
    .B1(_15002_),
    .B2(_15003_),
    .C1(_14424_),
    .Y(_15005_));
 sky130_fd_sc_hd__nand2_1 _42207_ (.A(_15004_),
    .B(_15005_),
    .Y(_15006_));
 sky130_fd_sc_hd__nand3_1 _42208_ (.A(_14988_),
    .B(_14989_),
    .C(_15006_),
    .Y(_15007_));
 sky130_fd_sc_hd__a21o_1 _42209_ (.A1(_14988_),
    .A2(_14989_),
    .B1(_15006_),
    .X(_15008_));
 sky130_fd_sc_hd__a21bo_1 _42210_ (.A1(_13613_),
    .A2(_14450_),
    .B1_N(_14451_),
    .X(_15010_));
 sky130_fd_sc_hd__buf_1 _42211_ (.A(_12234_),
    .X(_15011_));
 sky130_fd_sc_hd__a41oi_1 _42212_ (.A1(_14439_),
    .A2(_15011_),
    .A3(_13605_),
    .A4(_14443_),
    .B1(_14446_),
    .Y(_15012_));
 sky130_fd_sc_hd__buf_1 _42213_ (.A(_09764_),
    .X(_15013_));
 sky130_fd_sc_hd__buf_1 _42214_ (.A(_12225_),
    .X(_15014_));
 sky130_fd_sc_hd__o21ai_1 _42215_ (.A1(_15013_),
    .A2(_12236_),
    .B1(_15014_),
    .Y(_15015_));
 sky130_fd_sc_hd__or2_1 _42216_ (.A(_12225_),
    .B(_12236_),
    .X(_15016_));
 sky130_fd_sc_hd__o2bb2a_1 _42217_ (.A1_N(_15015_),
    .A2_N(_15016_),
    .B1(_14441_),
    .B2(_12232_),
    .X(_15017_));
 sky130_fd_sc_hd__a21boi_1 _42218_ (.A1(_15011_),
    .A2(_14443_),
    .B1_N(_15017_),
    .Y(_15018_));
 sky130_fd_sc_hd__and3b_1 _42219_ (.A_N(_15017_),
    .B(_15011_),
    .C(_14443_),
    .X(_15019_));
 sky130_fd_sc_hd__or2b_1 _42220_ (.A(_15014_),
    .B_N(_13610_),
    .X(_15021_));
 sky130_fd_sc_hd__o211a_1 _42221_ (.A1(_15018_),
    .A2(_15019_),
    .B1(_15013_),
    .C1(_15021_),
    .X(_15022_));
 sky130_fd_sc_hd__a211oi_1 _42222_ (.A1(_15013_),
    .A2(_15021_),
    .B1(_15018_),
    .C1(_15019_),
    .Y(_15023_));
 sky130_fd_sc_hd__or3_2 _42223_ (.A(_15012_),
    .B(_15022_),
    .C(_15023_),
    .X(_15024_));
 sky130_fd_sc_hd__o21a_1 _42224_ (.A1(_15022_),
    .A2(_15023_),
    .B1(_15012_),
    .X(_15025_));
 sky130_fd_sc_hd__inv_2 _42225_ (.A(_15025_),
    .Y(_15026_));
 sky130_fd_sc_hd__nand4_2 _42226_ (.A(_15024_),
    .B(_13602_),
    .C(_13600_),
    .D(_15026_),
    .Y(_15027_));
 sky130_fd_sc_hd__a32o_1 _42227_ (.A1(_13600_),
    .A2(_12224_),
    .A3(_14437_),
    .B1(_15024_),
    .B2(_15026_),
    .X(_15028_));
 sky130_fd_sc_hd__and3_1 _42228_ (.A(_15010_),
    .B(_15027_),
    .C(_15028_),
    .X(_15029_));
 sky130_fd_sc_hd__a21oi_1 _42229_ (.A1(_15027_),
    .A2(_15028_),
    .B1(_15010_),
    .Y(_15030_));
 sky130_fd_sc_hd__nor2_1 _42230_ (.A(_15029_),
    .B(_15030_),
    .Y(_15032_));
 sky130_fd_sc_hd__a21o_1 _42231_ (.A1(_14436_),
    .A2(_14454_),
    .B1(_14456_),
    .X(_15033_));
 sky130_fd_sc_hd__xor2_1 _42232_ (.A(_15032_),
    .B(_15033_),
    .X(_15034_));
 sky130_fd_sc_hd__a21oi_1 _42233_ (.A1(_15007_),
    .A2(_15008_),
    .B1(_15034_),
    .Y(_15035_));
 sky130_fd_sc_hd__nand3_1 _42234_ (.A(_15008_),
    .B(_15034_),
    .C(_15007_),
    .Y(_15036_));
 sky130_fd_sc_hd__and2b_1 _42235_ (.A_N(_15035_),
    .B(_15036_),
    .X(_15037_));
 sky130_fd_sc_hd__o21a_1 _42236_ (.A1(_14462_),
    .A2(_07330_),
    .B1(_08659_),
    .X(_15038_));
 sky130_fd_sc_hd__or2_1 _42237_ (.A(_15038_),
    .B(_14470_),
    .X(_15039_));
 sky130_fd_sc_hd__nand2_1 _42238_ (.A(_14470_),
    .B(_15038_),
    .Y(_15040_));
 sky130_fd_sc_hd__o22a_1 _42239_ (.A1(_13664_),
    .A2(_13667_),
    .B1(_07330_),
    .B2(_07331_),
    .X(_15041_));
 sky130_fd_sc_hd__or3_1 _42240_ (.A(_04099_),
    .B(_05602_),
    .C(_15041_),
    .X(_15043_));
 sky130_fd_sc_hd__a21oi_1 _42241_ (.A1(_15039_),
    .A2(_15040_),
    .B1(_15043_),
    .Y(_15044_));
 sky130_fd_sc_hd__nand3_1 _42242_ (.A(_15043_),
    .B(_15039_),
    .C(_15040_),
    .Y(_15045_));
 sky130_fd_sc_hd__and2b_1 _42243_ (.A_N(_15044_),
    .B(_15045_),
    .X(_15046_));
 sky130_fd_sc_hd__a21oi_1 _42244_ (.A1(_14464_),
    .A2(_14475_),
    .B1(_14473_),
    .Y(_15047_));
 sky130_fd_sc_hd__xnor2_1 _42245_ (.A(_15046_),
    .B(_15047_),
    .Y(_15048_));
 sky130_fd_sc_hd__a211oi_1 _42246_ (.A1(_04097_),
    .A2(_05606_),
    .B1(_07351_),
    .C1(_15048_),
    .Y(_15049_));
 sky130_fd_sc_hd__o21ai_1 _42247_ (.A1(_13688_),
    .A2(_14462_),
    .B1(_13664_),
    .Y(_15050_));
 sky130_fd_sc_hd__o21a_1 _42248_ (.A1(_07351_),
    .A2(_15050_),
    .B1(_15048_),
    .X(_15051_));
 sky130_fd_sc_hd__a211oi_2 _42249_ (.A1(_14477_),
    .A2(_14480_),
    .B1(_15049_),
    .C1(_15051_),
    .Y(_15052_));
 sky130_fd_sc_hd__o211a_1 _42250_ (.A1(_15049_),
    .A2(_15051_),
    .B1(_14477_),
    .C1(_14480_),
    .X(_15054_));
 sky130_fd_sc_hd__a21o_1 _42251_ (.A1(_14486_),
    .A2(_14487_),
    .B1(_14484_),
    .X(_15055_));
 sky130_fd_sc_hd__o21ai_1 _42252_ (.A1(_15052_),
    .A2(_15054_),
    .B1(_15055_),
    .Y(_15056_));
 sky130_fd_sc_hd__or3_1 _42253_ (.A(_15052_),
    .B(_15054_),
    .C(_15055_),
    .X(_15057_));
 sky130_fd_sc_hd__and2_1 _42254_ (.A(_15056_),
    .B(_15057_),
    .X(_15058_));
 sky130_fd_sc_hd__xnor2_1 _42255_ (.A(_15037_),
    .B(_15058_),
    .Y(_15059_));
 sky130_fd_sc_hd__a21o_1 _42256_ (.A1(_14984_),
    .A2(_14985_),
    .B1(_14944_),
    .X(_15060_));
 sky130_fd_sc_hd__nand2_2 _42257_ (.A(_15059_),
    .B(_15060_),
    .Y(_15061_));
 sky130_fd_sc_hd__a31o_1 _42258_ (.A1(_14944_),
    .A2(_14984_),
    .A3(_14986_),
    .B1(_15061_),
    .X(_15062_));
 sky130_fd_sc_hd__nand3_2 _42259_ (.A(_14944_),
    .B(_14984_),
    .C(_14986_),
    .Y(_15063_));
 sky130_fd_sc_hd__a21o_1 _42260_ (.A1(_15063_),
    .A2(_15060_),
    .B1(_15059_),
    .X(_15065_));
 sky130_fd_sc_hd__o211ai_2 _42261_ (.A1(_14409_),
    .A2(_14496_),
    .B1(_15062_),
    .C1(_15065_),
    .Y(_15066_));
 sky130_fd_sc_hd__inv_2 _42262_ (.A(net68),
    .Y(_15067_));
 sky130_fd_sc_hd__a211oi_4 _42263_ (.A1(_15062_),
    .A2(_15065_),
    .B1(_14409_),
    .C1(_14496_),
    .Y(_15068_));
 sky130_fd_sc_hd__o2bb2a_1 _42264_ (.A1_N(_14288_),
    .A2_N(_14337_),
    .B1(_14335_),
    .B2(_14307_),
    .X(_15069_));
 sky130_fd_sc_hd__and3_1 _42265_ (.A(_08412_),
    .B(_13495_),
    .C(_14275_),
    .X(_15070_));
 sky130_fd_sc_hd__buf_1 _42266_ (.A(_13490_),
    .X(_15071_));
 sky130_fd_sc_hd__a2bb2o_1 _42267_ (.A1_N(_08413_),
    .A2_N(_13494_),
    .B1(_15070_),
    .B2(_15071_),
    .X(_15072_));
 sky130_fd_sc_hd__clkbuf_2 _42268_ (.A(_13488_),
    .X(_15073_));
 sky130_fd_sc_hd__o22a_1 _42269_ (.A1(_15071_),
    .A2(_08417_),
    .B1(_07084_),
    .B2(_13488_),
    .X(_15074_));
 sky130_fd_sc_hd__a21oi_1 _42270_ (.A1(_07084_),
    .A2(_15073_),
    .B1(_15074_),
    .Y(_15076_));
 sky130_fd_sc_hd__xnor2_1 _42271_ (.A(_15072_),
    .B(_15076_),
    .Y(_15077_));
 sky130_fd_sc_hd__xnor2_1 _42272_ (.A(_14275_),
    .B(_15077_),
    .Y(_15078_));
 sky130_fd_sc_hd__nor2_1 _42273_ (.A(_14279_),
    .B(_14281_),
    .Y(_15079_));
 sky130_fd_sc_hd__or2_1 _42274_ (.A(_15078_),
    .B(_15079_),
    .X(_15080_));
 sky130_fd_sc_hd__or3b_1 _42275_ (.A(_14279_),
    .B(_14281_),
    .C_N(_15078_),
    .X(_15081_));
 sky130_fd_sc_hd__a221o_1 _42276_ (.A1(_15080_),
    .A2(_15081_),
    .B1(_14274_),
    .B2(_14287_),
    .C1(_14285_),
    .X(_15082_));
 sky130_fd_sc_hd__a21o_1 _42277_ (.A1(_14274_),
    .A2(_14287_),
    .B1(_14285_),
    .X(_15083_));
 sky130_fd_sc_hd__and2_1 _42278_ (.A(_15080_),
    .B(_15081_),
    .X(_15084_));
 sky130_fd_sc_hd__nand2_1 _42279_ (.A(_15083_),
    .B(_15084_),
    .Y(_15085_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _42280_ (.A(_13426_),
    .X(_15087_));
 sky130_fd_sc_hd__o211a_1 _42281_ (.A1(_14296_),
    .A2(_14294_),
    .B1(_12419_),
    .C1(_15087_),
    .X(_15088_));
 sky130_fd_sc_hd__nor2_1 _42282_ (.A(_14290_),
    .B(_13430_),
    .Y(_15089_));
 sky130_fd_sc_hd__o21ai_1 _42283_ (.A1(_12420_),
    .A2(_14296_),
    .B1(_14294_),
    .Y(_15090_));
 sky130_fd_sc_hd__o21ai_1 _42284_ (.A1(_14296_),
    .A2(_12432_),
    .B1(_12421_),
    .Y(_15091_));
 sky130_fd_sc_hd__a21boi_1 _42285_ (.A1(_14294_),
    .A2(_15090_),
    .B1_N(_15091_),
    .Y(_15092_));
 sky130_fd_sc_hd__o21bai_1 _42286_ (.A1(_14293_),
    .A2(_15089_),
    .B1_N(_15092_),
    .Y(_15093_));
 sky130_fd_sc_hd__or3b_1 _42287_ (.A(_14293_),
    .B(_15089_),
    .C_N(_15092_),
    .X(_15094_));
 sky130_fd_sc_hd__and2_1 _42288_ (.A(_15093_),
    .B(_15094_),
    .X(_15095_));
 sky130_fd_sc_hd__xnor2_1 _42289_ (.A(_15088_),
    .B(_15095_),
    .Y(_15096_));
 sky130_fd_sc_hd__or2b_1 _42290_ (.A(_15096_),
    .B_N(_14301_),
    .X(_15098_));
 sky130_fd_sc_hd__or2b_1 _42291_ (.A(_14301_),
    .B_N(_15096_),
    .X(_15099_));
 sky130_fd_sc_hd__nand2_1 _42292_ (.A(_15098_),
    .B(_15099_),
    .Y(_15100_));
 sky130_fd_sc_hd__o21bai_2 _42293_ (.A1(_14304_),
    .A2(_14307_),
    .B1_N(_15100_),
    .Y(_15101_));
 sky130_fd_sc_hd__and2_1 _42294_ (.A(_15098_),
    .B(_15099_),
    .X(_15102_));
 sky130_fd_sc_hd__or3_1 _42295_ (.A(_14304_),
    .B(_14307_),
    .C(_15102_),
    .X(_15103_));
 sky130_fd_sc_hd__o21bai_1 _42296_ (.A1(_14330_),
    .A2(_14333_),
    .B1_N(_14331_),
    .Y(_15104_));
 sky130_fd_sc_hd__a21bo_1 _42297_ (.A1(_13468_),
    .A2(_14324_),
    .B1_N(_14325_),
    .X(_15105_));
 sky130_fd_sc_hd__a41oi_2 _42298_ (.A1(_14319_),
    .A2(_14312_),
    .A3(_13458_),
    .A4(_14316_),
    .B1(_14321_),
    .Y(_15106_));
 sky130_fd_sc_hd__o21ai_1 _42299_ (.A1(_13455_),
    .A2(_07119_),
    .B1(_14313_),
    .Y(_15107_));
 sky130_fd_sc_hd__or2_1 _42300_ (.A(_14313_),
    .B(_07119_),
    .X(_15109_));
 sky130_fd_sc_hd__o2bb2a_1 _42301_ (.A1_N(_15107_),
    .A2_N(_15109_),
    .B1(_14314_),
    .B2(_14319_),
    .X(_15110_));
 sky130_fd_sc_hd__a21boi_1 _42302_ (.A1(_14312_),
    .A2(_14316_),
    .B1_N(_15110_),
    .Y(_15111_));
 sky130_fd_sc_hd__and3b_1 _42303_ (.A_N(_15110_),
    .B(_14312_),
    .C(_14316_),
    .X(_15112_));
 sky130_fd_sc_hd__buf_1 _42304_ (.A(_13455_),
    .X(_15113_));
 sky130_fd_sc_hd__buf_1 _42305_ (.A(_14313_),
    .X(_15114_));
 sky130_fd_sc_hd__or2b_1 _42306_ (.A(_15114_),
    .B_N(_14310_),
    .X(_15115_));
 sky130_fd_sc_hd__o211a_1 _42307_ (.A1(_15111_),
    .A2(_15112_),
    .B1(_15113_),
    .C1(_15115_),
    .X(_15116_));
 sky130_fd_sc_hd__a211oi_1 _42308_ (.A1(_15113_),
    .A2(_15115_),
    .B1(_15111_),
    .C1(_15112_),
    .Y(_15117_));
 sky130_fd_sc_hd__or3_2 _42309_ (.A(_15106_),
    .B(_15116_),
    .C(_15117_),
    .X(_15118_));
 sky130_fd_sc_hd__o21a_1 _42310_ (.A1(_15116_),
    .A2(_15117_),
    .B1(_15106_),
    .X(_15120_));
 sky130_fd_sc_hd__inv_2 _42311_ (.A(_15120_),
    .Y(_15121_));
 sky130_fd_sc_hd__nand4_2 _42312_ (.A(_15118_),
    .B(_13456_),
    .C(_13463_),
    .D(_15121_),
    .Y(_15122_));
 sky130_fd_sc_hd__a22o_1 _42313_ (.A1(_13463_),
    .A2(_13456_),
    .B1(_15121_),
    .B2(_15118_),
    .X(_15123_));
 sky130_fd_sc_hd__and3_1 _42314_ (.A(_15105_),
    .B(_15122_),
    .C(_15123_),
    .X(_15124_));
 sky130_fd_sc_hd__a21oi_1 _42315_ (.A1(_15122_),
    .A2(_15123_),
    .B1(_15105_),
    .Y(_15125_));
 sky130_fd_sc_hd__nor2_1 _42316_ (.A(_15124_),
    .B(_15125_),
    .Y(_15126_));
 sky130_fd_sc_hd__xor2_1 _42317_ (.A(_15104_),
    .B(_15126_),
    .X(_15127_));
 sky130_fd_sc_hd__a21oi_1 _42318_ (.A1(_15101_),
    .A2(_15103_),
    .B1(_15127_),
    .Y(_15128_));
 sky130_fd_sc_hd__and3_1 _42319_ (.A(_15101_),
    .B(_15103_),
    .C(_15127_),
    .X(_15129_));
 sky130_fd_sc_hd__nor2_1 _42320_ (.A(_15128_),
    .B(_15129_),
    .Y(_15131_));
 sky130_fd_sc_hd__a21o_1 _42321_ (.A1(_15082_),
    .A2(_15085_),
    .B1(_15131_),
    .X(_15132_));
 sky130_fd_sc_hd__nand3_1 _42322_ (.A(_15131_),
    .B(_15085_),
    .C(_15082_),
    .Y(_15133_));
 sky130_fd_sc_hd__nand2_1 _42323_ (.A(_15132_),
    .B(_15133_),
    .Y(_15134_));
 sky130_fd_sc_hd__nand3_1 _42324_ (.A(_14489_),
    .B(_14491_),
    .C(_15134_),
    .Y(_15135_));
 sky130_fd_sc_hd__a21o_1 _42325_ (.A1(_14489_),
    .A2(_14491_),
    .B1(_15134_),
    .X(_15136_));
 sky130_fd_sc_hd__nand2_1 _42326_ (.A(_15135_),
    .B(_15136_),
    .Y(_15137_));
 sky130_fd_sc_hd__xnor2_1 _42327_ (.A(_15069_),
    .B(_15137_),
    .Y(_15138_));
 sky130_fd_sc_hd__nor3_1 _42328_ (.A(_15067_),
    .B(net67),
    .C(_15138_),
    .Y(_15139_));
 sky130_fd_sc_hd__o21a_1 _42329_ (.A1(_15067_),
    .A2(net67),
    .B1(_15138_),
    .X(_15140_));
 sky130_fd_sc_hd__a21boi_1 _42330_ (.A1(_14349_),
    .A2(net72),
    .B1_N(_14498_),
    .Y(_15142_));
 sky130_fd_sc_hd__o21ai_1 _42331_ (.A1(_15139_),
    .A2(_15140_),
    .B1(_15142_),
    .Y(_15143_));
 sky130_fd_sc_hd__or3_1 _42332_ (.A(_15140_),
    .B(_15142_),
    .C(_15139_),
    .X(_15144_));
 sky130_fd_sc_hd__nand2_1 _42333_ (.A(_15143_),
    .B(_15144_),
    .Y(_15145_));
 sky130_fd_sc_hd__xnor2_1 _42334_ (.A(_14941_),
    .B(_15145_),
    .Y(_15146_));
 sky130_fd_sc_hd__o21ba_1 _42335_ (.A1(_14503_),
    .A2(_14598_),
    .B1_N(_14505_),
    .X(_15147_));
 sky130_fd_sc_hd__nand2_1 _42336_ (.A(_15146_),
    .B(_15147_),
    .Y(_15148_));
 sky130_fd_sc_hd__or2_1 _42337_ (.A(_15147_),
    .B(_15146_),
    .X(_15149_));
 sky130_fd_sc_hd__nand2_1 _42338_ (.A(_15148_),
    .B(_15149_),
    .Y(_15150_));
 sky130_fd_sc_hd__o21ai_2 _42339_ (.A1(_14870_),
    .A2(net62),
    .B1(_15150_),
    .Y(_15151_));
 sky130_fd_sc_hd__or3_4 _42340_ (.A(_14870_),
    .B(net62),
    .C(_15150_),
    .X(_15153_));
 sky130_fd_sc_hd__o2bb2a_1 _42341_ (.A1_N(_14272_),
    .A2_N(_14599_),
    .B1(_14600_),
    .B2(_14676_),
    .X(_15154_));
 sky130_fd_sc_hd__a21bo_2 _42342_ (.A1(_15151_),
    .A2(_15153_),
    .B1_N(_15154_),
    .X(_15155_));
 sky130_fd_sc_hd__nand3b_4 _42343_ (.A_N(_15154_),
    .B(_15151_),
    .C(_15153_),
    .Y(_15156_));
 sky130_fd_sc_hd__nand2_1 _42344_ (.A(_15155_),
    .B(_15156_),
    .Y(_15157_));
 sky130_fd_sc_hd__and3_1 _42345_ (.A(_14261_),
    .B(_14263_),
    .C(_14248_),
    .X(_15158_));
 sky130_fd_sc_hd__o21ba_1 _42346_ (.A1(_13803_),
    .A2(_14613_),
    .B1_N(_14612_),
    .X(_15159_));
 sky130_fd_sc_hd__inv_2 _42347_ (.A(_15159_),
    .Y(_15160_));
 sky130_fd_sc_hd__buf_1 _42348_ (.A(_15160_),
    .X(_15161_));
 sky130_fd_sc_hd__buf_2 _42349_ (.A(_13270_),
    .X(_15162_));
 sky130_fd_sc_hd__buf_2 _42350_ (.A(_14215_),
    .X(_15164_));
 sky130_fd_sc_hd__o21a_1 _42351_ (.A1(_13244_),
    .A2(_13254_),
    .B1(_14199_),
    .X(_15165_));
 sky130_fd_sc_hd__nor2_1 _42352_ (.A(_13252_),
    .B(_14197_),
    .Y(_15166_));
 sky130_fd_sc_hd__nand2_1 _42353_ (.A(_15166_),
    .B(_14199_),
    .Y(_15167_));
 sky130_fd_sc_hd__o22ai_2 _42354_ (.A1(_14197_),
    .A2(_15165_),
    .B1(_15167_),
    .B2(_14201_),
    .Y(_15168_));
 sky130_fd_sc_hd__o32a_2 _42355_ (.A1(_13219_),
    .A2(_13216_),
    .A3(_14179_),
    .B1(_14178_),
    .B2(_14177_),
    .X(_15169_));
 sky130_fd_sc_hd__nor2_1 _42356_ (.A(_14155_),
    .B(_14084_),
    .Y(_15170_));
 sky130_fd_sc_hd__nand2_1 _42357_ (.A(_14041_),
    .B(_14080_),
    .Y(_15171_));
 sky130_fd_sc_hd__nand2_1 _42358_ (.A(_14038_),
    .B(_15171_),
    .Y(_15172_));
 sky130_fd_sc_hd__o21ai_1 _42359_ (.A1(_13994_),
    .A2(_13986_),
    .B1(_13997_),
    .Y(_15173_));
 sky130_fd_sc_hd__o311a_2 _42360_ (.A1(_12912_),
    .A2(_11836_),
    .A3(_11837_),
    .B1(_11812_),
    .C1(_13939_),
    .X(_15175_));
 sky130_fd_sc_hd__a21oi_1 _42361_ (.A1(_13957_),
    .A2(_13945_),
    .B1(_15175_),
    .Y(_15176_));
 sky130_fd_sc_hd__a21o_1 _42362_ (.A1(_13944_),
    .A2(_13941_),
    .B1(_13957_),
    .X(_15177_));
 sky130_fd_sc_hd__nand3_2 _42363_ (.A(_13962_),
    .B(_15176_),
    .C(_15177_),
    .Y(_15178_));
 sky130_fd_sc_hd__o21a_1 _42364_ (.A1(_12914_),
    .A2(_13939_),
    .B1(_12895_),
    .X(_15179_));
 sky130_fd_sc_hd__a21oi_1 _42365_ (.A1(_13945_),
    .A2(_13941_),
    .B1(_13957_),
    .Y(_15180_));
 sky130_fd_sc_hd__o22ai_4 _42366_ (.A1(_15175_),
    .A2(_15179_),
    .B1(_15180_),
    .B2(_13951_),
    .Y(_15181_));
 sky130_fd_sc_hd__o211ai_4 _42367_ (.A1(_13968_),
    .A2(_12897_),
    .B1(_15178_),
    .C1(_15181_),
    .Y(_15182_));
 sky130_fd_sc_hd__a31o_1 _42368_ (.A1(_11823_),
    .A2(_11825_),
    .A3(_12900_),
    .B1(_10568_),
    .X(_15183_));
 sky130_fd_sc_hd__a221o_2 _42369_ (.A1(_13942_),
    .A2(_12911_),
    .B1(_15183_),
    .B2(_13946_),
    .C1(_11803_),
    .X(_15184_));
 sky130_fd_sc_hd__nand2_1 _42370_ (.A(_15182_),
    .B(_15184_),
    .Y(_15186_));
 sky130_fd_sc_hd__o211ai_1 _42371_ (.A1(_12896_),
    .A2(_13953_),
    .B1(_13950_),
    .C1(_12944_),
    .Y(_15187_));
 sky130_fd_sc_hd__a21oi_1 _42372_ (.A1(_15187_),
    .A2(_13962_),
    .B1(_13964_),
    .Y(_15188_));
 sky130_fd_sc_hd__a21oi_1 _42373_ (.A1(_13974_),
    .A2(_13966_),
    .B1(_15188_),
    .Y(_15189_));
 sky130_fd_sc_hd__nand2_1 _42374_ (.A(_15186_),
    .B(_15189_),
    .Y(_15190_));
 sky130_fd_sc_hd__a31oi_1 _42375_ (.A1(_15187_),
    .A2(_13962_),
    .A3(_13964_),
    .B1(_12952_),
    .Y(_15191_));
 sky130_fd_sc_hd__o21ai_1 _42376_ (.A1(_15188_),
    .A2(_15191_),
    .B1(_15182_),
    .Y(_15192_));
 sky130_fd_sc_hd__clkbuf_2 _42377_ (.A(_15192_),
    .X(_15193_));
 sky130_fd_sc_hd__a21oi_1 _42378_ (.A1(_15190_),
    .A2(_15193_),
    .B1(_13982_),
    .Y(_15194_));
 sky130_fd_sc_hd__a21o_1 _42379_ (.A1(_13974_),
    .A2(_13971_),
    .B1(_15188_),
    .X(_15195_));
 sky130_fd_sc_hd__inv_2 _42380_ (.A(_15184_),
    .Y(_15197_));
 sky130_fd_sc_hd__a31oi_2 _42381_ (.A1(_13974_),
    .A2(_15178_),
    .A3(_15181_),
    .B1(_15197_),
    .Y(_15198_));
 sky130_fd_sc_hd__o211a_1 _42382_ (.A1(_15195_),
    .A2(_15198_),
    .B1(_13982_),
    .C1(_15193_),
    .X(_15199_));
 sky130_fd_sc_hd__o31a_1 _42383_ (.A1(_13978_),
    .A2(_13975_),
    .A3(_13977_),
    .B1(_13989_),
    .X(_15200_));
 sky130_fd_sc_hd__o21ai_2 _42384_ (.A1(_15194_),
    .A2(_15199_),
    .B1(_15200_),
    .Y(_15201_));
 sky130_fd_sc_hd__a21o_1 _42385_ (.A1(_15190_),
    .A2(_15192_),
    .B1(_13969_),
    .X(_15202_));
 sky130_fd_sc_hd__o211ai_1 _42386_ (.A1(_15195_),
    .A2(_15198_),
    .B1(_13969_),
    .C1(_15193_),
    .Y(_15203_));
 sky130_fd_sc_hd__nand2_1 _42387_ (.A(_13973_),
    .B(_13989_),
    .Y(_15204_));
 sky130_fd_sc_hd__nand3_1 _42388_ (.A(_15202_),
    .B(_15203_),
    .C(_15204_),
    .Y(_15205_));
 sky130_fd_sc_hd__buf_1 _42389_ (.A(_10640_),
    .X(_15206_));
 sky130_fd_sc_hd__a21o_1 _42390_ (.A1(_15201_),
    .A2(_15205_),
    .B1(_15206_),
    .X(_15208_));
 sky130_fd_sc_hd__clkbuf_2 _42391_ (.A(_15205_),
    .X(_15209_));
 sky130_fd_sc_hd__nand3_1 _42392_ (.A(_15201_),
    .B(_15209_),
    .C(_15206_),
    .Y(_15210_));
 sky130_fd_sc_hd__nand3_2 _42393_ (.A(_15173_),
    .B(_15208_),
    .C(_15210_),
    .Y(_15211_));
 sky130_fd_sc_hd__a21oi_1 _42394_ (.A1(_15201_),
    .A2(_15209_),
    .B1(_15206_),
    .Y(_15212_));
 sky130_fd_sc_hd__and3_1 _42395_ (.A(_15201_),
    .B(_15205_),
    .C(_15206_),
    .X(_15213_));
 sky130_fd_sc_hd__o21a_1 _42396_ (.A1(_13994_),
    .A2(_13986_),
    .B1(_13997_),
    .X(_15214_));
 sky130_fd_sc_hd__o21ai_2 _42397_ (.A1(_15212_),
    .A2(_15213_),
    .B1(_15214_),
    .Y(_15215_));
 sky130_fd_sc_hd__buf_1 _42398_ (.A(_14008_),
    .X(_15216_));
 sky130_fd_sc_hd__clkbuf_2 _42399_ (.A(_15216_),
    .X(_15217_));
 sky130_fd_sc_hd__or4b_1 _42400_ (.A(_11905_),
    .B(_03125_),
    .C(_10500_),
    .D_N(_15217_),
    .X(_15219_));
 sky130_fd_sc_hd__o21a_1 _42401_ (.A1(_14012_),
    .A2(_14024_),
    .B1(_15219_),
    .X(_15220_));
 sky130_fd_sc_hd__a21oi_1 _42402_ (.A1(_12994_),
    .A2(_14008_),
    .B1(_14010_),
    .Y(_15221_));
 sky130_fd_sc_hd__a311oi_2 _42403_ (.A1(_14010_),
    .A2(_14007_),
    .A3(_04797_),
    .B1(_10648_),
    .C1(_15221_),
    .Y(_15222_));
 sky130_fd_sc_hd__clkbuf_2 _42404_ (.A(_11772_),
    .X(_15223_));
 sky130_fd_sc_hd__nand2_1 _42405_ (.A(_13006_),
    .B(_15223_),
    .Y(_15224_));
 sky130_fd_sc_hd__xor2_1 _42406_ (.A(_14013_),
    .B(_15224_),
    .X(_15225_));
 sky130_fd_sc_hd__xnor2_1 _42407_ (.A(_15222_),
    .B(_15225_),
    .Y(_15226_));
 sky130_fd_sc_hd__or2_2 _42408_ (.A(_13992_),
    .B(_15226_),
    .X(_15227_));
 sky130_fd_sc_hd__nand2_1 _42409_ (.A(_13992_),
    .B(_15226_),
    .Y(_15228_));
 sky130_fd_sc_hd__nand2_1 _42410_ (.A(_15227_),
    .B(_15228_),
    .Y(_15230_));
 sky130_fd_sc_hd__or2_1 _42411_ (.A(_15220_),
    .B(_15230_),
    .X(_15231_));
 sky130_fd_sc_hd__inv_2 _42412_ (.A(_15231_),
    .Y(_15232_));
 sky130_fd_sc_hd__o211a_1 _42413_ (.A1(_14012_),
    .A2(_14024_),
    .B1(_15219_),
    .C1(_15230_),
    .X(_15233_));
 sky130_fd_sc_hd__o2bb2ai_2 _42414_ (.A1_N(_15211_),
    .A2_N(_15215_),
    .B1(_15232_),
    .B2(_15233_),
    .Y(_15234_));
 sky130_fd_sc_hd__nor2_1 _42415_ (.A(_15232_),
    .B(_15233_),
    .Y(_15235_));
 sky130_fd_sc_hd__nand3_2 _42416_ (.A(_15211_),
    .B(_15215_),
    .C(_15235_),
    .Y(_15236_));
 sky130_fd_sc_hd__nor2_1 _42417_ (.A(_14035_),
    .B(_14036_),
    .Y(_15237_));
 sky130_fd_sc_hd__inv_2 _42418_ (.A(_15237_),
    .Y(_15238_));
 sky130_fd_sc_hd__nand2_1 _42419_ (.A(_14004_),
    .B(_15238_),
    .Y(_15239_));
 sky130_fd_sc_hd__nand2_1 _42420_ (.A(_14000_),
    .B(_15239_),
    .Y(_15241_));
 sky130_fd_sc_hd__a21oi_2 _42421_ (.A1(_15234_),
    .A2(_15236_),
    .B1(_15241_),
    .Y(_15242_));
 sky130_fd_sc_hd__and3_1 _42422_ (.A(_15241_),
    .B(_15234_),
    .C(_15236_),
    .X(_15243_));
 sky130_fd_sc_hd__a21bo_1 _42423_ (.A1(_14018_),
    .A2(_14021_),
    .B1_N(_10527_),
    .X(_15244_));
 sky130_fd_sc_hd__a21o_1 _42424_ (.A1(_14008_),
    .A2(_14043_),
    .B1(_15223_),
    .X(_15245_));
 sky130_fd_sc_hd__o211ai_2 _42425_ (.A1(_14014_),
    .A2(_14015_),
    .B1(_10527_),
    .C1(_12993_),
    .Y(_15246_));
 sky130_fd_sc_hd__a21o_1 _42426_ (.A1(_15246_),
    .A2(_14019_),
    .B1(_13008_),
    .X(_15247_));
 sky130_fd_sc_hd__a22oi_2 _42427_ (.A1(_15244_),
    .A2(_14007_),
    .B1(_15245_),
    .B2(_15247_),
    .Y(_15248_));
 sky130_fd_sc_hd__o2111ai_2 _42428_ (.A1(_15223_),
    .A2(_14043_),
    .B1(_12997_),
    .C1(_15244_),
    .D1(_15247_),
    .Y(_15249_));
 sky130_fd_sc_hd__inv_2 _42429_ (.A(_15249_),
    .Y(_15250_));
 sky130_fd_sc_hd__or3_1 _42430_ (.A(_15248_),
    .B(_14045_),
    .C(_15250_),
    .X(_15252_));
 sky130_fd_sc_hd__o21ai_1 _42431_ (.A1(_15250_),
    .A2(_15248_),
    .B1(_14045_),
    .Y(_15253_));
 sky130_fd_sc_hd__o211a_1 _42432_ (.A1(_14048_),
    .A2(_14050_),
    .B1(_15252_),
    .C1(_15253_),
    .X(_15254_));
 sky130_fd_sc_hd__a211oi_1 _42433_ (.A1(_15252_),
    .A2(_15253_),
    .B1(_14048_),
    .C1(_14050_),
    .Y(_15255_));
 sky130_fd_sc_hd__nor2_1 _42434_ (.A(_15254_),
    .B(_15255_),
    .Y(_15256_));
 sky130_fd_sc_hd__a21bo_1 _42435_ (.A1(_10705_),
    .A2(_11768_),
    .B1_N(_07691_),
    .X(_15257_));
 sky130_fd_sc_hd__nand3_1 _42436_ (.A(_07692_),
    .B(_15257_),
    .C(_11749_),
    .Y(_15258_));
 sky130_fd_sc_hd__or2b_1 _42437_ (.A(_11753_),
    .B_N(_07691_),
    .X(_15259_));
 sky130_fd_sc_hd__and2_1 _42438_ (.A(_07690_),
    .B(_11768_),
    .X(_15260_));
 sky130_fd_sc_hd__o2bb2a_1 _42439_ (.A1_N(_15258_),
    .A2_N(_15259_),
    .B1(_15260_),
    .B2(_14062_),
    .X(_15261_));
 sky130_fd_sc_hd__and4bb_1 _42440_ (.A_N(_15260_),
    .B_N(_14062_),
    .C(_15258_),
    .D(_15259_),
    .X(_15263_));
 sky130_fd_sc_hd__a21oi_1 _42441_ (.A1(_04646_),
    .A2(_09148_),
    .B1(_07675_),
    .Y(_15264_));
 sky130_fd_sc_hd__and3_1 _42442_ (.A(_04646_),
    .B(_07675_),
    .C(_10687_),
    .X(_15265_));
 sky130_fd_sc_hd__o21a_1 _42443_ (.A1(_15264_),
    .A2(_15265_),
    .B1(_10677_),
    .X(_15266_));
 sky130_fd_sc_hd__a211oi_1 _42444_ (.A1(_11738_),
    .A2(_06400_),
    .B1(_15264_),
    .C1(_11748_),
    .Y(_15267_));
 sky130_fd_sc_hd__and2b_1 _42445_ (.A_N(_03349_),
    .B(_11752_),
    .X(_15268_));
 sky130_fd_sc_hd__and4bb_2 _42446_ (.A_N(_15266_),
    .B_N(_15267_),
    .C(_13050_),
    .D(_15268_),
    .X(_15269_));
 sky130_fd_sc_hd__o2bb2a_1 _42447_ (.A1_N(_13060_),
    .A2_N(_15268_),
    .B1(_15266_),
    .B2(_15267_),
    .X(_15270_));
 sky130_fd_sc_hd__o22ai_2 _42448_ (.A1(_15261_),
    .A2(_15263_),
    .B1(_15269_),
    .B2(_15270_),
    .Y(_15271_));
 sky130_fd_sc_hd__or4_2 _42449_ (.A(_15261_),
    .B(_15263_),
    .C(_15269_),
    .D(_15270_),
    .X(_15272_));
 sky130_fd_sc_hd__and3_1 _42450_ (.A(_15256_),
    .B(_15271_),
    .C(_15272_),
    .X(_15274_));
 sky130_fd_sc_hd__o2bb2a_1 _42451_ (.A1_N(_15272_),
    .A2_N(_15271_),
    .B1(_15254_),
    .B2(_15255_),
    .X(_15275_));
 sky130_fd_sc_hd__o211a_1 _42452_ (.A1(_15274_),
    .A2(_15275_),
    .B1(_14027_),
    .C1(_14030_),
    .X(_15276_));
 sky130_fd_sc_hd__a211o_1 _42453_ (.A1(_14027_),
    .A2(_14030_),
    .B1(_15274_),
    .C1(_15275_),
    .X(_15277_));
 sky130_fd_sc_hd__nor2_1 _42454_ (.A(_14071_),
    .B(_14072_),
    .Y(_15278_));
 sky130_fd_sc_hd__and3b_1 _42455_ (.A_N(_15276_),
    .B(_15277_),
    .C(_15278_),
    .X(_15279_));
 sky130_fd_sc_hd__and2b_1 _42456_ (.A_N(_15276_),
    .B(_15277_),
    .X(_15280_));
 sky130_fd_sc_hd__nor2_1 _42457_ (.A(_15278_),
    .B(_15280_),
    .Y(_15281_));
 sky130_fd_sc_hd__nor2_1 _42458_ (.A(_15279_),
    .B(_15281_),
    .Y(_15282_));
 sky130_fd_sc_hd__o21bai_1 _42459_ (.A1(_15242_),
    .A2(_15243_),
    .B1_N(_15282_),
    .Y(_15283_));
 sky130_fd_sc_hd__nand3_2 _42460_ (.A(_15241_),
    .B(_15234_),
    .C(_15236_),
    .Y(_15285_));
 sky130_fd_sc_hd__nand3b_1 _42461_ (.A_N(_15242_),
    .B(_15285_),
    .C(_15282_),
    .Y(_15286_));
 sky130_fd_sc_hd__nand3b_4 _42462_ (.A_N(_15172_),
    .B(_15283_),
    .C(_15286_),
    .Y(_15287_));
 sky130_fd_sc_hd__a32oi_4 _42463_ (.A1(_13931_),
    .A2(_13995_),
    .A3(_13999_),
    .B1(_14005_),
    .B2(_15238_),
    .Y(_15288_));
 sky130_fd_sc_hd__nand2_1 _42464_ (.A(_15234_),
    .B(_15236_),
    .Y(_15289_));
 sky130_fd_sc_hd__o2bb2ai_4 _42465_ (.A1_N(_15288_),
    .A2_N(_15289_),
    .B1(_15279_),
    .B2(_15281_),
    .Y(_15290_));
 sky130_fd_sc_hd__o21ai_1 _42466_ (.A1(_15242_),
    .A2(_15243_),
    .B1(_15282_),
    .Y(_15291_));
 sky130_fd_sc_hd__o211ai_4 _42467_ (.A1(_15290_),
    .A2(_15243_),
    .B1(_15172_),
    .C1(_15291_),
    .Y(_15292_));
 sky130_fd_sc_hd__a21boi_1 _42468_ (.A1(_14074_),
    .A2(_14077_),
    .B1_N(_14076_),
    .Y(_15293_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _42469_ (.A(_13112_),
    .X(_15294_));
 sky130_fd_sc_hd__and4b_1 _42470_ (.A_N(_13112_),
    .B(_13205_),
    .C(_09391_),
    .D(_13124_),
    .X(_15296_));
 sky130_fd_sc_hd__a22o_1 _42471_ (.A1(_15294_),
    .A2(_13125_),
    .B1(_15296_),
    .B2(_13113_),
    .X(_15297_));
 sky130_fd_sc_hd__nand2_1 _42472_ (.A(_13139_),
    .B(_13112_),
    .Y(_15298_));
 sky130_fd_sc_hd__clkbuf_2 _42473_ (.A(_13113_),
    .X(_15299_));
 sky130_fd_sc_hd__o22ai_2 _42474_ (.A1(_13121_),
    .A2(_15298_),
    .B1(_15299_),
    .B2(_14109_),
    .Y(_15300_));
 sky130_fd_sc_hd__xnor2_1 _42475_ (.A(_15297_),
    .B(_15300_),
    .Y(_15301_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _42476_ (.A(_12026_),
    .X(_15302_));
 sky130_fd_sc_hd__and3_1 _42477_ (.A(_15302_),
    .B(_12002_),
    .C(_13139_),
    .X(_15303_));
 sky130_fd_sc_hd__nor2_2 _42478_ (.A(_12011_),
    .B(_15302_),
    .Y(_15304_));
 sky130_fd_sc_hd__or3b_1 _42479_ (.A(_12025_),
    .B(_15302_),
    .C_N(_12002_),
    .X(_15305_));
 sky130_fd_sc_hd__or3b_1 _42480_ (.A(_15303_),
    .B(_15304_),
    .C_N(_15305_),
    .X(_15307_));
 sky130_fd_sc_hd__xor2_1 _42481_ (.A(_13113_),
    .B(_15307_),
    .X(_15308_));
 sky130_fd_sc_hd__and3_1 _42482_ (.A(_14124_),
    .B(_14126_),
    .C(_13151_),
    .X(_15309_));
 sky130_fd_sc_hd__o21ai_1 _42483_ (.A1(_14123_),
    .A2(_15309_),
    .B1(_13134_),
    .Y(_15310_));
 sky130_fd_sc_hd__a21oi_1 _42484_ (.A1(_14124_),
    .A2(_13151_),
    .B1(_14123_),
    .Y(_15311_));
 sky130_fd_sc_hd__o211ai_2 _42485_ (.A1(_13156_),
    .A2(net186),
    .B1(_15311_),
    .C1(_13135_),
    .Y(_15312_));
 sky130_fd_sc_hd__o221a_1 _42486_ (.A1(_13135_),
    .A2(_14123_),
    .B1(_15310_),
    .B2(_14104_),
    .C1(_15312_),
    .X(_15313_));
 sky130_fd_sc_hd__nor2_1 _42487_ (.A(_15308_),
    .B(_15313_),
    .Y(_15314_));
 sky130_fd_sc_hd__nand2_1 _42488_ (.A(_15308_),
    .B(_15313_),
    .Y(_15315_));
 sky130_fd_sc_hd__inv_2 _42489_ (.A(_15315_),
    .Y(_15316_));
 sky130_fd_sc_hd__o221a_1 _42490_ (.A1(_13136_),
    .A2(_14104_),
    .B1(_15314_),
    .B2(_15316_),
    .C1(_14112_),
    .X(_15318_));
 sky130_fd_sc_hd__a211o_1 _42491_ (.A1(_14102_),
    .A2(_14112_),
    .B1(_15314_),
    .C1(_15316_),
    .X(_15319_));
 sky130_fd_sc_hd__and2b_1 _42492_ (.A_N(_15318_),
    .B(_15319_),
    .X(_15320_));
 sky130_fd_sc_hd__nand2_1 _42493_ (.A(_15301_),
    .B(_15320_),
    .Y(_15321_));
 sky130_fd_sc_hd__or2_1 _42494_ (.A(_15301_),
    .B(_15320_),
    .X(_15322_));
 sky130_fd_sc_hd__and2_1 _42495_ (.A(_15321_),
    .B(_15322_),
    .X(_15323_));
 sky130_fd_sc_hd__o21ba_1 _42496_ (.A1(_14142_),
    .A2(_14138_),
    .B1_N(_14139_),
    .X(_15324_));
 sky130_fd_sc_hd__o21ai_1 _42497_ (.A1(_14067_),
    .A2(_14059_),
    .B1(_14068_),
    .Y(_15325_));
 sky130_fd_sc_hd__nand2_1 _42498_ (.A(_11753_),
    .B(_14056_),
    .Y(_15326_));
 sky130_fd_sc_hd__a21bo_1 _42499_ (.A1(_14057_),
    .A2(_14058_),
    .B1_N(_15326_),
    .X(_15327_));
 sky130_fd_sc_hd__buf_1 _42500_ (.A(_11969_),
    .X(_15329_));
 sky130_fd_sc_hd__nand2_1 _42501_ (.A(_10802_),
    .B(_10758_),
    .Y(_15330_));
 sky130_fd_sc_hd__and3_1 _42502_ (.A(_11968_),
    .B(_15329_),
    .C(_15330_),
    .X(_15331_));
 sky130_fd_sc_hd__buf_1 _42503_ (.A(_10802_),
    .X(_15332_));
 sky130_fd_sc_hd__and3_1 _42504_ (.A(_11970_),
    .B(_10758_),
    .C(_15332_),
    .X(_15333_));
 sky130_fd_sc_hd__nor3_1 _42505_ (.A(_13051_),
    .B(_15331_),
    .C(_15333_),
    .Y(_15334_));
 sky130_fd_sc_hd__o21a_1 _42506_ (.A1(_15331_),
    .A2(_15333_),
    .B1(_13051_),
    .X(_15335_));
 sky130_fd_sc_hd__nor2_1 _42507_ (.A(_15334_),
    .B(_15335_),
    .Y(_15336_));
 sky130_fd_sc_hd__and2_1 _42508_ (.A(_15327_),
    .B(_15336_),
    .X(_15337_));
 sky130_fd_sc_hd__inv_2 _42509_ (.A(_15337_),
    .Y(_15338_));
 sky130_fd_sc_hd__or2_1 _42510_ (.A(_15336_),
    .B(_15327_),
    .X(_15340_));
 sky130_fd_sc_hd__and3_1 _42511_ (.A(_15338_),
    .B(_14128_),
    .C(_15340_),
    .X(_15341_));
 sky130_fd_sc_hd__a21oi_1 _42512_ (.A1(_15340_),
    .A2(_15338_),
    .B1(_14128_),
    .Y(_15342_));
 sky130_fd_sc_hd__nor2_1 _42513_ (.A(_15341_),
    .B(_15342_),
    .Y(_15343_));
 sky130_fd_sc_hd__xnor2_1 _42514_ (.A(_15325_),
    .B(_15343_),
    .Y(_15344_));
 sky130_fd_sc_hd__and3_1 _42515_ (.A(_14133_),
    .B(_14135_),
    .C(_15344_),
    .X(_15345_));
 sky130_fd_sc_hd__a21oi_1 _42516_ (.A1(_14133_),
    .A2(_14135_),
    .B1(_15344_),
    .Y(_15346_));
 sky130_fd_sc_hd__nor3_1 _42517_ (.A(_15324_),
    .B(_15345_),
    .C(_15346_),
    .Y(_15347_));
 sky130_fd_sc_hd__o21a_1 _42518_ (.A1(_15345_),
    .A2(_15346_),
    .B1(_15324_),
    .X(_15348_));
 sky130_fd_sc_hd__nor2_1 _42519_ (.A(_15347_),
    .B(_15348_),
    .Y(_15349_));
 sky130_fd_sc_hd__xnor2_1 _42520_ (.A(_15323_),
    .B(_15349_),
    .Y(_15351_));
 sky130_fd_sc_hd__nor2_1 _42521_ (.A(_15293_),
    .B(_15351_),
    .Y(_15352_));
 sky130_fd_sc_hd__and2_1 _42522_ (.A(_15351_),
    .B(_15293_),
    .X(_15353_));
 sky130_fd_sc_hd__nor2_2 _42523_ (.A(_15352_),
    .B(_15353_),
    .Y(_15354_));
 sky130_fd_sc_hd__a21oi_1 _42524_ (.A1(_13171_),
    .A2(_13176_),
    .B1(_14144_),
    .Y(_15355_));
 sky130_fd_sc_hd__a21o_1 _42525_ (.A1(_14120_),
    .A2(_14146_),
    .B1(_15355_),
    .X(_15356_));
 sky130_fd_sc_hd__xor2_4 _42526_ (.A(_15354_),
    .B(_15356_),
    .X(_15357_));
 sky130_fd_sc_hd__a21o_1 _42527_ (.A1(_15287_),
    .A2(_15292_),
    .B1(_15357_),
    .X(_15358_));
 sky130_fd_sc_hd__nand3_1 _42528_ (.A(_15287_),
    .B(_15292_),
    .C(_15357_),
    .Y(_15359_));
 sky130_fd_sc_hd__o211ai_2 _42529_ (.A1(_14088_),
    .A2(_15170_),
    .B1(_15358_),
    .C1(_15359_),
    .Y(_15360_));
 sky130_fd_sc_hd__inv_2 _42530_ (.A(_15357_),
    .Y(_15362_));
 sky130_fd_sc_hd__a21o_1 _42531_ (.A1(_15287_),
    .A2(_15292_),
    .B1(_15362_),
    .X(_15363_));
 sky130_fd_sc_hd__nand3_1 _42532_ (.A(_15287_),
    .B(_15292_),
    .C(_15362_),
    .Y(_15364_));
 sky130_fd_sc_hd__o22a_1 _42533_ (.A1(_14085_),
    .A2(_14087_),
    .B1(_14155_),
    .B2(_14084_),
    .X(_15365_));
 sky130_fd_sc_hd__nand3_2 _42534_ (.A(_15363_),
    .B(_15364_),
    .C(_15365_),
    .Y(_15366_));
 sky130_fd_sc_hd__o211ai_4 _42535_ (.A1(_13213_),
    .A2(_13214_),
    .B1(_14172_),
    .C1(_14173_),
    .Y(_15367_));
 sky130_fd_sc_hd__o31ai_2 _42536_ (.A1(_14169_),
    .A2(_14166_),
    .A3(_14168_),
    .B1(_14172_),
    .Y(_15368_));
 sky130_fd_sc_hd__buf_1 _42537_ (.A(\delay_line[1][15] ),
    .X(_15369_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _42538_ (.A(_15369_),
    .X(_15370_));
 sky130_fd_sc_hd__nand3b_1 _42539_ (.A_N(_14091_),
    .B(_14096_),
    .C(_14098_),
    .Y(_15371_));
 sky130_fd_sc_hd__a2bb2o_1 _42540_ (.A1_N(_14167_),
    .A2_N(_15370_),
    .B1(_14098_),
    .B2(_15371_),
    .X(_15373_));
 sky130_fd_sc_hd__or4bb_1 _42541_ (.A(_14167_),
    .B(_15369_),
    .C_N(_14098_),
    .D_N(_15371_),
    .X(_15374_));
 sky130_fd_sc_hd__a221oi_1 _42542_ (.A1(_15373_),
    .A2(_15374_),
    .B1(_14100_),
    .B2(_14116_),
    .C1(_14114_),
    .Y(_15375_));
 sky130_fd_sc_hd__o211a_1 _42543_ (.A1(_14114_),
    .A2(_14118_),
    .B1(_15373_),
    .C1(_15374_),
    .X(_15376_));
 sky130_fd_sc_hd__nor2_1 _42544_ (.A(_15375_),
    .B(_15376_),
    .Y(_15377_));
 sky130_fd_sc_hd__xnor2_1 _42545_ (.A(_14166_),
    .B(_15377_),
    .Y(_15378_));
 sky130_fd_sc_hd__xnor2_1 _42546_ (.A(_15368_),
    .B(_15378_),
    .Y(_15379_));
 sky130_fd_sc_hd__o21ai_2 _42547_ (.A1(_14149_),
    .A2(_14151_),
    .B1(_15379_),
    .Y(_15380_));
 sky130_fd_sc_hd__o21bai_1 _42548_ (.A1(_14089_),
    .A2(_14150_),
    .B1_N(_14149_),
    .Y(_15381_));
 sky130_fd_sc_hd__or2_1 _42549_ (.A(_15381_),
    .B(_15379_),
    .X(_15382_));
 sky130_fd_sc_hd__nand2_2 _42550_ (.A(_15380_),
    .B(_15382_),
    .Y(_15384_));
 sky130_fd_sc_hd__xor2_2 _42551_ (.A(_15367_),
    .B(_15384_),
    .X(_15385_));
 sky130_fd_sc_hd__inv_2 _42552_ (.A(_15385_),
    .Y(_15386_));
 sky130_fd_sc_hd__a21o_1 _42553_ (.A1(_15360_),
    .A2(_15366_),
    .B1(_15386_),
    .X(_15387_));
 sky130_fd_sc_hd__a32oi_4 _42554_ (.A1(_13929_),
    .A2(_14156_),
    .A3(_14158_),
    .B1(_14164_),
    .B2(_14180_),
    .Y(_15388_));
 sky130_fd_sc_hd__clkbuf_2 _42555_ (.A(_15360_),
    .X(_15389_));
 sky130_fd_sc_hd__nand3_1 _42556_ (.A(_15386_),
    .B(_15389_),
    .C(_15366_),
    .Y(_15390_));
 sky130_fd_sc_hd__nand3_1 _42557_ (.A(_15387_),
    .B(_15388_),
    .C(_15390_),
    .Y(_15391_));
 sky130_fd_sc_hd__nand2_1 _42558_ (.A(_15389_),
    .B(_15366_),
    .Y(_15392_));
 sky130_fd_sc_hd__a21oi_1 _42559_ (.A1(_15386_),
    .A2(_15392_),
    .B1(_15388_),
    .Y(_15393_));
 sky130_fd_sc_hd__nand3_1 _42560_ (.A(_15389_),
    .B(_15366_),
    .C(_15385_),
    .Y(_15395_));
 sky130_fd_sc_hd__nand2_2 _42561_ (.A(_15393_),
    .B(_15395_),
    .Y(_15396_));
 sky130_fd_sc_hd__nand2_1 _42562_ (.A(_15391_),
    .B(_15396_),
    .Y(_15397_));
 sky130_fd_sc_hd__nor2_1 _42563_ (.A(_15169_),
    .B(_15397_),
    .Y(_15398_));
 sky130_fd_sc_hd__or2_1 _42564_ (.A(_14189_),
    .B(_14190_),
    .X(_15399_));
 sky130_fd_sc_hd__a22o_1 _42565_ (.A1(_15397_),
    .A2(_15169_),
    .B1(_14192_),
    .B2(_15399_),
    .X(_15400_));
 sky130_fd_sc_hd__nand2_1 _42566_ (.A(_15397_),
    .B(_15169_),
    .Y(_15401_));
 sky130_fd_sc_hd__nand3b_1 _42567_ (.A_N(_15169_),
    .B(_15391_),
    .C(_15396_),
    .Y(_15402_));
 sky130_fd_sc_hd__o21ai_4 _42568_ (.A1(_14187_),
    .A2(_14184_),
    .B1(_15399_),
    .Y(_15403_));
 sky130_fd_sc_hd__a21oi_2 _42569_ (.A1(_15401_),
    .A2(_15402_),
    .B1(_15403_),
    .Y(_15404_));
 sky130_fd_sc_hd__o21ba_1 _42570_ (.A1(_15398_),
    .A2(_15400_),
    .B1_N(_15404_),
    .X(_15406_));
 sky130_fd_sc_hd__nand2_1 _42571_ (.A(_15168_),
    .B(_15406_),
    .Y(_15407_));
 sky130_fd_sc_hd__buf_6 _42572_ (.A(_15407_),
    .X(_15408_));
 sky130_fd_sc_hd__o21bai_2 _42573_ (.A1(_15398_),
    .A2(_15400_),
    .B1_N(_15404_),
    .Y(_15409_));
 sky130_fd_sc_hd__o221ai_2 _42574_ (.A1(_14197_),
    .A2(_15165_),
    .B1(_15167_),
    .B2(_14201_),
    .C1(_15409_),
    .Y(_15410_));
 sky130_fd_sc_hd__clkbuf_2 _42575_ (.A(_15410_),
    .X(_15411_));
 sky130_fd_sc_hd__o211ai_4 _42576_ (.A1(_15162_),
    .A2(_15164_),
    .B1(_15408_),
    .C1(_15411_),
    .Y(_15412_));
 sky130_fd_sc_hd__nand2_1 _42577_ (.A(_15407_),
    .B(_15410_),
    .Y(_15413_));
 sky130_fd_sc_hd__a21oi_2 _42578_ (.A1(_11588_),
    .A2(_12727_),
    .B1(_13270_),
    .Y(_15414_));
 sky130_fd_sc_hd__a21oi_1 _42579_ (.A1(_15413_),
    .A2(_15414_),
    .B1(_10935_),
    .Y(_15415_));
 sky130_fd_sc_hd__a21o_1 _42580_ (.A1(_15408_),
    .A2(_15411_),
    .B1(_14204_),
    .X(_15417_));
 sky130_fd_sc_hd__nand2_1 _42581_ (.A(_15412_),
    .B(_15417_),
    .Y(_15418_));
 sky130_fd_sc_hd__a22oi_2 _42582_ (.A1(_15412_),
    .A2(_15415_),
    .B1(_15418_),
    .B2(_12875_),
    .Y(_15419_));
 sky130_fd_sc_hd__o21ai_1 _42583_ (.A1(_12885_),
    .A2(_14213_),
    .B1(_14216_),
    .Y(_15420_));
 sky130_fd_sc_hd__buf_1 _42584_ (.A(_15420_),
    .X(_15421_));
 sky130_fd_sc_hd__o21ai_1 _42585_ (.A1(_15161_),
    .A2(_15419_),
    .B1(_15421_),
    .Y(_15422_));
 sky130_fd_sc_hd__clkbuf_2 _42586_ (.A(_15415_),
    .X(_15423_));
 sky130_fd_sc_hd__a221oi_4 _42587_ (.A1(_15412_),
    .A2(_15423_),
    .B1(_15418_),
    .B2(_12875_),
    .C1(_15159_),
    .Y(_15424_));
 sky130_fd_sc_hd__a21bo_1 _42588_ (.A1(_14242_),
    .A2(_14222_),
    .B1_N(_14226_),
    .X(_15425_));
 sky130_fd_sc_hd__o21ai_1 _42589_ (.A1(_15414_),
    .A2(_15413_),
    .B1(_15415_),
    .Y(_15426_));
 sky130_fd_sc_hd__o211a_1 _42590_ (.A1(_13270_),
    .A2(_14215_),
    .B1(_15407_),
    .C1(_15411_),
    .X(_15428_));
 sky130_fd_sc_hd__clkbuf_2 _42591_ (.A(_14204_),
    .X(_15429_));
 sky130_fd_sc_hd__a21oi_1 _42592_ (.A1(_15408_),
    .A2(_15411_),
    .B1(_15429_),
    .Y(_15430_));
 sky130_fd_sc_hd__o21ai_1 _42593_ (.A1(_15428_),
    .A2(_15430_),
    .B1(_12885_),
    .Y(_15431_));
 sky130_fd_sc_hd__a21oi_1 _42594_ (.A1(_15426_),
    .A2(_15431_),
    .B1(_15161_),
    .Y(_15432_));
 sky130_fd_sc_hd__inv_2 _42595_ (.A(_15420_),
    .Y(_15433_));
 sky130_fd_sc_hd__o21ai_1 _42596_ (.A1(_15424_),
    .A2(_15432_),
    .B1(_15433_),
    .Y(_15434_));
 sky130_fd_sc_hd__o211ai_1 _42597_ (.A1(_15422_),
    .A2(_15424_),
    .B1(_15425_),
    .C1(_15434_),
    .Y(_15435_));
 sky130_fd_sc_hd__o21ai_1 _42598_ (.A1(_15424_),
    .A2(_15432_),
    .B1(_15421_),
    .Y(_15436_));
 sky130_fd_sc_hd__a21boi_1 _42599_ (.A1(_14242_),
    .A2(_14222_),
    .B1_N(_14226_),
    .Y(_15437_));
 sky130_fd_sc_hd__a21o_1 _42600_ (.A1(_15426_),
    .A2(_15431_),
    .B1(_15160_),
    .X(_15439_));
 sky130_fd_sc_hd__nand2_1 _42601_ (.A(_15419_),
    .B(_15161_),
    .Y(_15440_));
 sky130_fd_sc_hd__nand3_1 _42602_ (.A(_15439_),
    .B(_15433_),
    .C(_15440_),
    .Y(_15441_));
 sky130_fd_sc_hd__nand3_1 _42603_ (.A(_15436_),
    .B(_15437_),
    .C(_15441_),
    .Y(_15442_));
 sky130_fd_sc_hd__or3b_1 _42604_ (.A(_00395_),
    .B(_12153_),
    .C_N(_14259_),
    .X(_15443_));
 sky130_fd_sc_hd__o211a_1 _42605_ (.A1(_02004_),
    .A2(_03560_),
    .B1(_13294_),
    .C1(_15443_),
    .X(_15444_));
 sky130_fd_sc_hd__o21ai_1 _42606_ (.A1(_02004_),
    .A2(_03560_),
    .B1(_15443_),
    .Y(_15445_));
 sky130_fd_sc_hd__and2_1 _42607_ (.A(_12875_),
    .B(_15445_),
    .X(_15446_));
 sky130_fd_sc_hd__or2_1 _42608_ (.A(_15444_),
    .B(_15446_),
    .X(_15447_));
 sky130_fd_sc_hd__a21o_1 _42609_ (.A1(_15435_),
    .A2(_15442_),
    .B1(_15447_),
    .X(_15448_));
 sky130_fd_sc_hd__a21boi_4 _42610_ (.A1(_14601_),
    .A2(_14673_),
    .B1_N(_14674_),
    .Y(_15450_));
 sky130_fd_sc_hd__and3_1 _42611_ (.A(_15421_),
    .B(_15440_),
    .C(_15439_),
    .X(_15451_));
 sky130_fd_sc_hd__nand2_1 _42612_ (.A(_15425_),
    .B(_15434_),
    .Y(_15452_));
 sky130_fd_sc_hd__o211ai_2 _42613_ (.A1(_15451_),
    .A2(_15452_),
    .B1(_15442_),
    .C1(_15447_),
    .Y(_15453_));
 sky130_fd_sc_hd__nand3_4 _42614_ (.A(_15448_),
    .B(_15450_),
    .C(_15453_),
    .Y(_15454_));
 sky130_fd_sc_hd__nor2_1 _42615_ (.A(_15444_),
    .B(_15446_),
    .Y(_15455_));
 sky130_fd_sc_hd__a21o_1 _42616_ (.A1(_15435_),
    .A2(_15442_),
    .B1(_15455_),
    .X(_15456_));
 sky130_fd_sc_hd__a31oi_2 _42617_ (.A1(_15436_),
    .A2(_15437_),
    .A3(_15441_),
    .B1(_15447_),
    .Y(_15457_));
 sky130_fd_sc_hd__o21ai_1 _42618_ (.A1(_15451_),
    .A2(_15452_),
    .B1(_15457_),
    .Y(_15458_));
 sky130_fd_sc_hd__nand3b_1 _42619_ (.A_N(_15450_),
    .B(_15456_),
    .C(_15458_),
    .Y(_15459_));
 sky130_fd_sc_hd__buf_6 _42620_ (.A(_15459_),
    .X(_15461_));
 sky130_fd_sc_hd__o211ai_4 _42621_ (.A1(_14237_),
    .A2(_15158_),
    .B1(_15454_),
    .C1(_15461_),
    .Y(_15462_));
 sky130_fd_sc_hd__a31o_1 _42622_ (.A1(_14261_),
    .A2(_14263_),
    .A3(_14248_),
    .B1(_14237_),
    .X(_15463_));
 sky130_fd_sc_hd__a21o_1 _42623_ (.A1(_15454_),
    .A2(_15461_),
    .B1(_15463_),
    .X(_15464_));
 sky130_fd_sc_hd__nand3_1 _42624_ (.A(_15157_),
    .B(_15462_),
    .C(_15464_),
    .Y(_15465_));
 sky130_fd_sc_hd__o211a_1 _42625_ (.A1(_14237_),
    .A2(_15158_),
    .B1(_15454_),
    .C1(_15459_),
    .X(_15466_));
 sky130_fd_sc_hd__a21oi_2 _42626_ (.A1(_15454_),
    .A2(_15461_),
    .B1(_15463_),
    .Y(_15467_));
 sky130_fd_sc_hd__o21bai_1 _42627_ (.A1(_15466_),
    .A2(_15467_),
    .B1_N(_15157_),
    .Y(_15468_));
 sky130_fd_sc_hd__nand3_1 _42628_ (.A(_14821_),
    .B(_15465_),
    .C(_15468_),
    .Y(_15469_));
 sky130_fd_sc_hd__a31o_1 _42629_ (.A1(_14255_),
    .A2(_14270_),
    .A3(_14683_),
    .B1(_14681_),
    .X(_15470_));
 sky130_fd_sc_hd__o21ai_2 _42630_ (.A1(_15466_),
    .A2(_15467_),
    .B1(_15157_),
    .Y(_15472_));
 sky130_fd_sc_hd__nand4_2 _42631_ (.A(_15155_),
    .B(_15156_),
    .C(_15462_),
    .D(_15464_),
    .Y(_15473_));
 sky130_fd_sc_hd__nand3_1 _42632_ (.A(_15470_),
    .B(_15472_),
    .C(_15473_),
    .Y(_15474_));
 sky130_fd_sc_hd__nand2_1 _42633_ (.A(_15469_),
    .B(_15474_),
    .Y(_15475_));
 sky130_fd_sc_hd__o21ai_1 _42634_ (.A1(_14253_),
    .A2(_14247_),
    .B1(_14268_),
    .Y(_15476_));
 sky130_fd_sc_hd__and3b_1 _42635_ (.A_N(_14259_),
    .B(_13926_),
    .C(_14257_),
    .X(_15477_));
 sky130_fd_sc_hd__o21a_1 _42636_ (.A1(_00399_),
    .A2(_02005_),
    .B1(_12880_),
    .X(_15478_));
 sky130_fd_sc_hd__buf_2 _42637_ (.A(_10436_),
    .X(_15479_));
 sky130_fd_sc_hd__o221ai_2 _42638_ (.A1(_12147_),
    .A2(_13926_),
    .B1(_15477_),
    .B2(_15478_),
    .C1(_15479_),
    .Y(_15480_));
 sky130_fd_sc_hd__or3b_1 _42639_ (.A(_13926_),
    .B(_13844_),
    .C_N(_12783_),
    .X(_15481_));
 sky130_fd_sc_hd__a211o_1 _42640_ (.A1(_15481_),
    .A2(_15479_),
    .B1(_15477_),
    .C1(_15478_),
    .X(_15483_));
 sky130_fd_sc_hd__nand2_1 _42641_ (.A(_15480_),
    .B(_15483_),
    .Y(_15484_));
 sky130_fd_sc_hd__o21a_1 _42642_ (.A1(_12149_),
    .A2(_13292_),
    .B1(_15479_),
    .X(_15485_));
 sky130_fd_sc_hd__xor2_1 _42643_ (.A(_15484_),
    .B(_15485_),
    .X(_15486_));
 sky130_fd_sc_hd__buf_2 _42644_ (.A(_08967_),
    .X(_15487_));
 sky130_fd_sc_hd__xor2_2 _42645_ (.A(_15487_),
    .B(_14706_),
    .X(_15488_));
 sky130_fd_sc_hd__o21ai_1 _42646_ (.A1(_03033_),
    .A2(_08974_),
    .B1(_10429_),
    .Y(_15489_));
 sky130_fd_sc_hd__or3_1 _42647_ (.A(_03033_),
    .B(_09007_),
    .C(_08974_),
    .X(_15490_));
 sky130_fd_sc_hd__buf_2 _42648_ (.A(_09006_),
    .X(_15491_));
 sky130_fd_sc_hd__a21o_1 _42649_ (.A1(_08978_),
    .A2(_15491_),
    .B1(_12782_),
    .X(_15492_));
 sky130_fd_sc_hd__o21ai_1 _42650_ (.A1(_08978_),
    .A2(_15491_),
    .B1(_12782_),
    .Y(_15494_));
 sky130_fd_sc_hd__a22o_1 _42651_ (.A1(_15489_),
    .A2(_15490_),
    .B1(_15492_),
    .B2(_15494_),
    .X(_15495_));
 sky130_fd_sc_hd__nand4_1 _42652_ (.A(_15489_),
    .B(_15490_),
    .C(_15492_),
    .D(_15494_),
    .Y(_15496_));
 sky130_fd_sc_hd__nand2_1 _42653_ (.A(_15495_),
    .B(_15496_),
    .Y(_15497_));
 sky130_fd_sc_hd__a2bb2o_1 _42654_ (.A1_N(_09002_),
    .A2_N(_10321_),
    .B1(_15479_),
    .B2(_10435_),
    .X(_15498_));
 sky130_fd_sc_hd__buf_2 _42655_ (.A(_08978_),
    .X(_15499_));
 sky130_fd_sc_hd__nor2_1 _42656_ (.A(_15491_),
    .B(_12782_),
    .Y(_15500_));
 sky130_fd_sc_hd__a21oi_2 _42657_ (.A1(_10324_),
    .A2(_15499_),
    .B1(_15500_),
    .Y(_15501_));
 sky130_fd_sc_hd__a2bb2o_1 _42658_ (.A1_N(_14705_),
    .A2_N(_14708_),
    .B1(_15498_),
    .B2(_15501_),
    .X(_15502_));
 sky130_fd_sc_hd__xnor2_1 _42659_ (.A(_15497_),
    .B(_15502_),
    .Y(_15503_));
 sky130_fd_sc_hd__xnor2_2 _42660_ (.A(_15488_),
    .B(_15503_),
    .Y(_15505_));
 sky130_fd_sc_hd__nor2_1 _42661_ (.A(_15486_),
    .B(_15505_),
    .Y(_15506_));
 sky130_fd_sc_hd__and2_1 _42662_ (.A(_15486_),
    .B(_15505_),
    .X(_15507_));
 sky130_fd_sc_hd__or2_1 _42663_ (.A(_15506_),
    .B(_15507_),
    .X(_15508_));
 sky130_fd_sc_hd__inv_2 _42664_ (.A(_15508_),
    .Y(_15509_));
 sky130_fd_sc_hd__nand2_1 _42665_ (.A(_15476_),
    .B(_15509_),
    .Y(_15510_));
 sky130_fd_sc_hd__clkbuf_2 _42666_ (.A(_15510_),
    .X(_15511_));
 sky130_fd_sc_hd__o211ai_2 _42667_ (.A1(_14253_),
    .A2(_14247_),
    .B1(_14268_),
    .C1(_15508_),
    .Y(_15512_));
 sky130_fd_sc_hd__o21ai_2 _42668_ (.A1(_14699_),
    .A2(_14700_),
    .B1(_14714_),
    .Y(_15513_));
 sky130_fd_sc_hd__a21oi_1 _42669_ (.A1(_15511_),
    .A2(_15512_),
    .B1(_15513_),
    .Y(_15514_));
 sky130_fd_sc_hd__and3_1 _42670_ (.A(_15513_),
    .B(_15510_),
    .C(_15512_),
    .X(_15516_));
 sky130_fd_sc_hd__nor2_1 _42671_ (.A(_15514_),
    .B(_15516_),
    .Y(_15517_));
 sky130_fd_sc_hd__nand2_1 _42672_ (.A(_15475_),
    .B(_15517_),
    .Y(_15518_));
 sky130_fd_sc_hd__a21o_1 _42673_ (.A1(_14255_),
    .A2(_14270_),
    .B1(_14683_),
    .X(_15519_));
 sky130_fd_sc_hd__a32oi_2 _42674_ (.A1(_14685_),
    .A2(_15519_),
    .A3(_14686_),
    .B1(_14723_),
    .B2(_14695_),
    .Y(_15520_));
 sky130_fd_sc_hd__clkbuf_2 _42675_ (.A(_15469_),
    .X(_15521_));
 sky130_fd_sc_hd__o211ai_1 _42676_ (.A1(_15514_),
    .A2(_15516_),
    .B1(_15521_),
    .C1(_15474_),
    .Y(_15522_));
 sky130_fd_sc_hd__nand3_2 _42677_ (.A(_15518_),
    .B(_15520_),
    .C(_15522_),
    .Y(_15523_));
 sky130_fd_sc_hd__o2bb2ai_1 _42678_ (.A1_N(_14723_),
    .A2_N(_14695_),
    .B1(_14687_),
    .B2(_14684_),
    .Y(_15524_));
 sky130_fd_sc_hd__a21o_1 _42679_ (.A1(_15511_),
    .A2(_15512_),
    .B1(_15513_),
    .X(_15525_));
 sky130_fd_sc_hd__nand3_1 _42680_ (.A(_15513_),
    .B(_15511_),
    .C(_15512_),
    .Y(_15527_));
 sky130_fd_sc_hd__nand4_1 _42681_ (.A(_15521_),
    .B(_15474_),
    .C(_15525_),
    .D(_15527_),
    .Y(_15528_));
 sky130_fd_sc_hd__o2bb2ai_1 _42682_ (.A1_N(_15521_),
    .A2_N(_15474_),
    .B1(_15514_),
    .B2(_15516_),
    .Y(_15529_));
 sky130_fd_sc_hd__nand3_2 _42683_ (.A(_15524_),
    .B(_15528_),
    .C(_15529_),
    .Y(_15530_));
 sky130_fd_sc_hd__o211a_1 _42684_ (.A1(_14817_),
    .A2(_14820_),
    .B1(_15523_),
    .C1(_15530_),
    .X(_15531_));
 sky130_fd_sc_hd__nand2_1 _42685_ (.A(_14729_),
    .B(_14764_),
    .Y(_15532_));
 sky130_fd_sc_hd__nand2_1 _42686_ (.A(_14736_),
    .B(_15532_),
    .Y(_15533_));
 sky130_fd_sc_hd__nand2_1 _42687_ (.A(_15523_),
    .B(_15530_),
    .Y(_15534_));
 sky130_fd_sc_hd__a21oi_1 _42688_ (.A1(_14818_),
    .A2(_14816_),
    .B1(_14820_),
    .Y(_15535_));
 sky130_fd_sc_hd__nand2_1 _42689_ (.A(_15534_),
    .B(_15535_),
    .Y(_15536_));
 sky130_fd_sc_hd__nand2_1 _42690_ (.A(_15533_),
    .B(_15536_),
    .Y(_15538_));
 sky130_fd_sc_hd__a21oi_1 _42691_ (.A1(_13861_),
    .A2(_14737_),
    .B1(_14759_),
    .Y(_15539_));
 sky130_fd_sc_hd__o21a_1 _42692_ (.A1(_13895_),
    .A2(_15539_),
    .B1(_14761_),
    .X(_15540_));
 sky130_fd_sc_hd__a21oi_2 _42693_ (.A1(_14756_),
    .A2(_14818_),
    .B1(_14815_),
    .Y(_15541_));
 sky130_fd_sc_hd__o22a_1 _42694_ (.A1(_15541_),
    .A2(_14815_),
    .B1(_14756_),
    .B2(_14817_),
    .X(_15542_));
 sky130_fd_sc_hd__a21oi_1 _42695_ (.A1(_15523_),
    .A2(_15530_),
    .B1(_15542_),
    .Y(_15543_));
 sky130_fd_sc_hd__o21bai_1 _42696_ (.A1(_15531_),
    .A2(_15543_),
    .B1_N(_15533_),
    .Y(_15544_));
 sky130_fd_sc_hd__clkbuf_2 _42697_ (.A(_15544_),
    .X(_15545_));
 sky130_fd_sc_hd__o211a_1 _42698_ (.A1(_15531_),
    .A2(_15538_),
    .B1(_15540_),
    .C1(_15545_),
    .X(_15546_));
 sky130_fd_sc_hd__o211ai_1 _42699_ (.A1(_14817_),
    .A2(_14820_),
    .B1(_15523_),
    .C1(_15530_),
    .Y(_15547_));
 sky130_fd_sc_hd__nand3_2 _42700_ (.A(_15533_),
    .B(_15547_),
    .C(_15536_),
    .Y(_15549_));
 sky130_fd_sc_hd__a21oi_1 _42701_ (.A1(_15545_),
    .A2(_15549_),
    .B1(_15540_),
    .Y(_15550_));
 sky130_fd_sc_hd__a2bb2o_1 _42702_ (.A1_N(_14765_),
    .A2_N(_14777_),
    .B1(_14775_),
    .B2(_14771_),
    .X(_15551_));
 sky130_fd_sc_hd__o21bai_1 _42703_ (.A1(_15546_),
    .A2(_15550_),
    .B1_N(_15551_),
    .Y(_15552_));
 sky130_fd_sc_hd__o2111ai_1 _42704_ (.A1(_13895_),
    .A2(_15539_),
    .B1(_14761_),
    .C1(_15545_),
    .D1(_15549_),
    .Y(_15553_));
 sky130_fd_sc_hd__a21o_1 _42705_ (.A1(_15545_),
    .A2(_15549_),
    .B1(_15540_),
    .X(_15554_));
 sky130_fd_sc_hd__nand3_1 _42706_ (.A(_15551_),
    .B(_15553_),
    .C(_15554_),
    .Y(_15555_));
 sky130_fd_sc_hd__and2_2 _42707_ (.A(_15552_),
    .B(_15555_),
    .X(_15556_));
 sky130_fd_sc_hd__inv_2 _42708_ (.A(_13916_),
    .Y(_15557_));
 sky130_fd_sc_hd__nand2_1 _42709_ (.A(_13914_),
    .B(_13915_),
    .Y(_15558_));
 sky130_fd_sc_hd__o21ai_1 _42710_ (.A1(_15557_),
    .A2(_15558_),
    .B1(_14786_),
    .Y(_15560_));
 sky130_fd_sc_hd__and4_1 _42711_ (.A(_13917_),
    .B(_13918_),
    .C(_14781_),
    .D(_14786_),
    .X(_15561_));
 sky130_fd_sc_hd__a22o_2 _42712_ (.A1(_14781_),
    .A2(_15560_),
    .B1(_13925_),
    .B2(_15561_),
    .X(_15562_));
 sky130_fd_sc_hd__xor2_4 _42713_ (.A(_15556_),
    .B(_15562_),
    .X(_00016_));
 sky130_fd_sc_hd__a21bo_1 _42714_ (.A1(_15552_),
    .A2(_15562_),
    .B1_N(_15555_),
    .X(_15563_));
 sky130_fd_sc_hd__a32o_1 _42715_ (.A1(_15470_),
    .A2(_15472_),
    .A3(_15473_),
    .B1(_15517_),
    .B2(_15521_),
    .X(_15564_));
 sky130_fd_sc_hd__or3_2 _42716_ (.A(_14259_),
    .B(_14258_),
    .C(_13844_),
    .X(_15565_));
 sky130_fd_sc_hd__buf_2 _42717_ (.A(_15479_),
    .X(_15566_));
 sky130_fd_sc_hd__nor2_1 _42718_ (.A(_12153_),
    .B(_03566_),
    .Y(_15567_));
 sky130_fd_sc_hd__a211o_1 _42719_ (.A1(_15565_),
    .A2(_15566_),
    .B1(_15567_),
    .C1(_15444_),
    .X(_15568_));
 sky130_fd_sc_hd__buf_1 _42720_ (.A(_15566_),
    .X(_15570_));
 sky130_fd_sc_hd__o211ai_2 _42721_ (.A1(_15567_),
    .A2(_15444_),
    .B1(_15565_),
    .C1(_15570_),
    .Y(_15571_));
 sky130_fd_sc_hd__a32o_1 _42722_ (.A1(_12783_),
    .A2(_14257_),
    .A3(_14258_),
    .B1(_15478_),
    .B2(_15565_),
    .X(_15572_));
 sky130_fd_sc_hd__and4_1 _42723_ (.A(_15568_),
    .B(_15571_),
    .C(_15572_),
    .D(_15570_),
    .X(_15573_));
 sky130_fd_sc_hd__clkbuf_2 _42724_ (.A(_15566_),
    .X(_15574_));
 sky130_fd_sc_hd__a22oi_1 _42725_ (.A1(_15572_),
    .A2(_15574_),
    .B1(_15568_),
    .B2(_15571_),
    .Y(_15575_));
 sky130_fd_sc_hd__clkbuf_2 _42726_ (.A(_15487_),
    .X(_15576_));
 sky130_fd_sc_hd__buf_2 _42727_ (.A(_15576_),
    .X(_15577_));
 sky130_fd_sc_hd__a21oi_1 _42728_ (.A1(_10429_),
    .A2(_12764_),
    .B1(_15577_),
    .Y(_15578_));
 sky130_fd_sc_hd__and3_2 _42729_ (.A(_15576_),
    .B(_10429_),
    .C(_12764_),
    .X(_15579_));
 sky130_fd_sc_hd__or3_1 _42730_ (.A(_10321_),
    .B(_09004_),
    .C(_10435_),
    .X(_15581_));
 sky130_fd_sc_hd__o21ai_1 _42731_ (.A1(_10321_),
    .A2(_09004_),
    .B1(_10435_),
    .Y(_15582_));
 sky130_fd_sc_hd__o21a_1 _42732_ (.A1(_15499_),
    .A2(_15491_),
    .B1(_15566_),
    .X(_15583_));
 sky130_fd_sc_hd__and4_1 _42733_ (.A(_15489_),
    .B(_15490_),
    .C(_15492_),
    .D(_15494_),
    .X(_15584_));
 sky130_fd_sc_hd__a211oi_1 _42734_ (.A1(_15581_),
    .A2(_15582_),
    .B1(_15583_),
    .C1(_15584_),
    .Y(_15585_));
 sky130_fd_sc_hd__o211a_1 _42735_ (.A1(_15583_),
    .A2(_15584_),
    .B1(_15581_),
    .C1(_15582_),
    .X(_15586_));
 sky130_fd_sc_hd__nor4_2 _42736_ (.A(_15578_),
    .B(_15579_),
    .C(_15585_),
    .D(_15586_),
    .Y(_15587_));
 sky130_fd_sc_hd__o22a_2 _42737_ (.A1(_15578_),
    .A2(_15579_),
    .B1(_15585_),
    .B2(_15586_),
    .X(_15588_));
 sky130_fd_sc_hd__nor4_1 _42738_ (.A(_15573_),
    .B(_15575_),
    .C(net149),
    .D(_15588_),
    .Y(_15589_));
 sky130_fd_sc_hd__o22a_1 _42739_ (.A1(_15573_),
    .A2(_15575_),
    .B1(net149),
    .B2(_15588_),
    .X(_15590_));
 sky130_fd_sc_hd__or2_1 _42740_ (.A(net144),
    .B(_15590_),
    .X(_15592_));
 sky130_fd_sc_hd__a21o_1 _42741_ (.A1(_15461_),
    .A2(_15462_),
    .B1(_15592_),
    .X(_15593_));
 sky130_fd_sc_hd__o211ai_2 _42742_ (.A1(_15589_),
    .A2(_15590_),
    .B1(_15461_),
    .C1(_15462_),
    .Y(_15594_));
 sky130_fd_sc_hd__a31o_1 _42743_ (.A1(_15480_),
    .A2(_15483_),
    .A3(_15485_),
    .B1(_15506_),
    .X(_15595_));
 sky130_fd_sc_hd__a21oi_2 _42744_ (.A1(_15593_),
    .A2(_15594_),
    .B1(_15595_),
    .Y(_15596_));
 sky130_fd_sc_hd__and3_1 _42745_ (.A(_15595_),
    .B(_15593_),
    .C(_15594_),
    .X(_15597_));
 sky130_fd_sc_hd__o21ai_1 _42746_ (.A1(_15466_),
    .A2(_15467_),
    .B1(_15156_),
    .Y(_15598_));
 sky130_fd_sc_hd__clkbuf_2 _42747_ (.A(_14861_),
    .X(_15599_));
 sky130_fd_sc_hd__o21bai_2 _42748_ (.A1(_14853_),
    .A2(_14851_),
    .B1_N(_15599_),
    .Y(_15600_));
 sky130_fd_sc_hd__nand2_1 _42749_ (.A(_14854_),
    .B(_15600_),
    .Y(_15601_));
 sky130_fd_sc_hd__a21boi_2 _42750_ (.A1(_14938_),
    .A2(_14936_),
    .B1_N(_14937_),
    .Y(_15603_));
 sky130_fd_sc_hd__or2_1 _42751_ (.A(_14543_),
    .B(_14823_),
    .X(_15604_));
 sky130_fd_sc_hd__o311a_1 _42752_ (.A1(_15604_),
    .A2(_14843_),
    .A3(_14846_),
    .B1(_14664_),
    .C1(_14656_),
    .X(_15605_));
 sky130_fd_sc_hd__nor2_2 _42753_ (.A(_14848_),
    .B(_15605_),
    .Y(_15606_));
 sky130_fd_sc_hd__a2bb2o_2 _42754_ (.A1_N(_14622_),
    .A2_N(_14825_),
    .B1(_14824_),
    .B2(_12640_),
    .X(_15607_));
 sky130_fd_sc_hd__and4bb_1 _42755_ (.A_N(_14832_),
    .B_N(_14637_),
    .C(_14633_),
    .D(_14631_),
    .X(_15608_));
 sky130_fd_sc_hd__a211o_1 _42756_ (.A1(_12664_),
    .A2(_14830_),
    .B1(_15608_),
    .C1(_14835_),
    .X(_15609_));
 sky130_fd_sc_hd__o21ai_1 _42757_ (.A1(_15607_),
    .A2(_14827_),
    .B1(_15609_),
    .Y(_15610_));
 sky130_fd_sc_hd__a211oi_2 _42758_ (.A1(_12664_),
    .A2(_14830_),
    .B1(_15608_),
    .C1(_14835_),
    .Y(_15611_));
 sky130_fd_sc_hd__inv_2 _42759_ (.A(_15607_),
    .Y(_15612_));
 sky130_fd_sc_hd__nand3_1 _42760_ (.A(_14839_),
    .B(_15611_),
    .C(_15612_),
    .Y(_15614_));
 sky130_fd_sc_hd__a32o_1 _42761_ (.A1(_13767_),
    .A2(_14649_),
    .A3(_08292_),
    .B1(_14841_),
    .B2(_08295_),
    .X(_15615_));
 sky130_fd_sc_hd__a21oi_1 _42762_ (.A1(_15610_),
    .A2(_15614_),
    .B1(_15615_),
    .Y(_15616_));
 sky130_fd_sc_hd__and3_1 _42763_ (.A(_15615_),
    .B(_15610_),
    .C(_15614_),
    .X(_15617_));
 sky130_fd_sc_hd__o2bb2a_1 _42764_ (.A1_N(_14919_),
    .A2_N(_14931_),
    .B1(_15616_),
    .B2(_15617_),
    .X(_15618_));
 sky130_fd_sc_hd__a21boi_1 _42765_ (.A1(_15615_),
    .A2(_14840_),
    .B1_N(_14838_),
    .Y(_15619_));
 sky130_fd_sc_hd__nand2_1 _42766_ (.A(_14919_),
    .B(_14931_),
    .Y(_15620_));
 sky130_fd_sc_hd__nor3_1 _42767_ (.A(_15620_),
    .B(_15616_),
    .C(_15617_),
    .Y(_15621_));
 sky130_fd_sc_hd__or2_1 _42768_ (.A(_15619_),
    .B(_15621_),
    .X(_15622_));
 sky130_fd_sc_hd__o21ai_1 _42769_ (.A1(_15618_),
    .A2(_15621_),
    .B1(_15619_),
    .Y(_15623_));
 sky130_fd_sc_hd__o21ai_4 _42770_ (.A1(_15618_),
    .A2(_15622_),
    .B1(_15623_),
    .Y(_15625_));
 sky130_fd_sc_hd__xnor2_1 _42771_ (.A(_15606_),
    .B(_15625_),
    .Y(_15626_));
 sky130_fd_sc_hd__xnor2_2 _42772_ (.A(_15599_),
    .B(_15626_),
    .Y(_15627_));
 sky130_fd_sc_hd__xnor2_2 _42773_ (.A(_15603_),
    .B(_15627_),
    .Y(_15628_));
 sky130_fd_sc_hd__xnor2_1 _42774_ (.A(_15601_),
    .B(_15628_),
    .Y(_15629_));
 sky130_fd_sc_hd__and4_2 _42775_ (.A(_09901_),
    .B(_14369_),
    .C(_14958_),
    .D(_14368_),
    .X(_15630_));
 sky130_fd_sc_hd__o21ba_1 _42776_ (.A1(_14958_),
    .A2(_09901_),
    .B1_N(_14369_),
    .X(_15631_));
 sky130_fd_sc_hd__o22a_1 _42777_ (.A1(_14959_),
    .A2(_14960_),
    .B1(_15631_),
    .B2(_14370_),
    .X(_15632_));
 sky130_fd_sc_hd__o21ai_1 _42778_ (.A1(_14957_),
    .A2(_14379_),
    .B1(_14961_),
    .Y(_15633_));
 sky130_fd_sc_hd__o21a_1 _42779_ (.A1(_15630_),
    .A2(_15632_),
    .B1(_15633_),
    .X(_15634_));
 sky130_fd_sc_hd__nor2_1 _42780_ (.A(_15630_),
    .B(_15632_),
    .Y(_15636_));
 sky130_fd_sc_hd__o211a_2 _42781_ (.A1(_14957_),
    .A2(_14379_),
    .B1(_14961_),
    .C1(_15636_),
    .X(_15637_));
 sky130_fd_sc_hd__or2b_1 _42782_ (.A(_14952_),
    .B_N(_14951_),
    .X(_15638_));
 sky130_fd_sc_hd__o21a_1 _42783_ (.A1(_13521_),
    .A2(_14947_),
    .B1(_14945_),
    .X(_15639_));
 sky130_fd_sc_hd__a31oi_1 _42784_ (.A1(_12327_),
    .A2(_14353_),
    .A3(_07251_),
    .B1(_15639_),
    .Y(_15640_));
 sky130_fd_sc_hd__and3_1 _42785_ (.A(_15638_),
    .B(_14956_),
    .C(_15640_),
    .X(_15641_));
 sky130_fd_sc_hd__a21oi_1 _42786_ (.A1(_15638_),
    .A2(_14956_),
    .B1(_15640_),
    .Y(_15642_));
 sky130_fd_sc_hd__nor4_1 _42787_ (.A(_15634_),
    .B(_15637_),
    .C(_15641_),
    .D(_15642_),
    .Y(_15643_));
 sky130_fd_sc_hd__a21o_1 _42788_ (.A1(_14968_),
    .A2(_14982_),
    .B1(_14980_),
    .X(_15644_));
 sky130_fd_sc_hd__xnor2_1 _42789_ (.A(_14970_),
    .B(_14972_),
    .Y(_15645_));
 sky130_fd_sc_hd__a311o_1 _42790_ (.A1(_14387_),
    .A2(_14977_),
    .A3(_14388_),
    .B1(_14975_),
    .C1(_15645_),
    .X(_15647_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _42791_ (.A(_14392_),
    .X(_15648_));
 sky130_fd_sc_hd__o2111a_1 _42792_ (.A1(_15648_),
    .A2(_14391_),
    .B1(_14387_),
    .C1(_14970_),
    .D1(_14977_),
    .X(_15649_));
 sky130_fd_sc_hd__o21ai_2 _42793_ (.A1(_14975_),
    .A2(_15649_),
    .B1(_15645_),
    .Y(_15650_));
 sky130_fd_sc_hd__nand3_2 _42794_ (.A(_15644_),
    .B(_15647_),
    .C(_15650_),
    .Y(_15651_));
 sky130_fd_sc_hd__a221o_1 _42795_ (.A1(_15647_),
    .A2(_15650_),
    .B1(_14968_),
    .B2(_14982_),
    .C1(_14980_),
    .X(_15652_));
 sky130_fd_sc_hd__nand2_2 _42796_ (.A(_15651_),
    .B(_15652_),
    .Y(_15653_));
 sky130_fd_sc_hd__o22a_2 _42797_ (.A1(_15634_),
    .A2(_15637_),
    .B1(_15641_),
    .B2(_15642_),
    .X(_15654_));
 sky130_fd_sc_hd__or2_2 _42798_ (.A(_15653_),
    .B(_15654_),
    .X(_15655_));
 sky130_fd_sc_hd__o21ai_1 _42799_ (.A1(net79),
    .A2(_15654_),
    .B1(_15653_),
    .Y(_15656_));
 sky130_fd_sc_hd__o21ai_4 _42800_ (.A1(net79),
    .A2(_15655_),
    .B1(_15656_),
    .Y(_15658_));
 sky130_fd_sc_hd__a21o_1 _42801_ (.A1(_14967_),
    .A2(_14986_),
    .B1(_15658_),
    .X(_15659_));
 sky130_fd_sc_hd__nand2_1 _42802_ (.A(_14967_),
    .B(_14986_),
    .Y(_15660_));
 sky130_fd_sc_hd__inv_2 _42803_ (.A(_15660_),
    .Y(_15661_));
 sky130_fd_sc_hd__nand2_1 _42804_ (.A(_15658_),
    .B(_15661_),
    .Y(_15662_));
 sky130_fd_sc_hd__nand3_1 _42805_ (.A(_14988_),
    .B(_14989_),
    .C(_15004_),
    .Y(_15663_));
 sky130_fd_sc_hd__buf_1 _42806_ (.A(_12181_),
    .X(_15664_));
 sky130_fd_sc_hd__nand2_1 _42807_ (.A(_14994_),
    .B(_14995_),
    .Y(_15665_));
 sky130_fd_sc_hd__a21o_1 _42808_ (.A1(_14994_),
    .A2(_14993_),
    .B1(_14995_),
    .X(_15666_));
 sky130_fd_sc_hd__a22oi_2 _42809_ (.A1(_15664_),
    .A2(_14992_),
    .B1(_15665_),
    .B2(_15666_),
    .Y(_15667_));
 sky130_fd_sc_hd__buf_1 _42810_ (.A(_13632_),
    .X(_15669_));
 sky130_fd_sc_hd__and3_1 _42811_ (.A(_15664_),
    .B(_12182_),
    .C(_15669_),
    .X(_15670_));
 sky130_fd_sc_hd__nand3_1 _42812_ (.A(_14999_),
    .B(_15000_),
    .C(_15001_),
    .Y(_15671_));
 sky130_fd_sc_hd__o211a_1 _42813_ (.A1(_15667_),
    .A2(_15670_),
    .B1(_15000_),
    .C1(_15671_),
    .X(_15672_));
 sky130_fd_sc_hd__a211o_1 _42814_ (.A1(_15000_),
    .A2(_15671_),
    .B1(_15667_),
    .C1(_15670_),
    .X(_15673_));
 sky130_fd_sc_hd__and2b_1 _42815_ (.A_N(_15672_),
    .B(_15673_),
    .X(_15674_));
 sky130_fd_sc_hd__a21oi_1 _42816_ (.A1(_15005_),
    .A2(_15663_),
    .B1(_15674_),
    .Y(_15675_));
 sky130_fd_sc_hd__inv_2 _42817_ (.A(_15675_),
    .Y(_15676_));
 sky130_fd_sc_hd__nand3_2 _42818_ (.A(_15005_),
    .B(_15663_),
    .C(_15674_),
    .Y(_15677_));
 sky130_fd_sc_hd__buf_2 _42819_ (.A(_15011_),
    .X(_15678_));
 sky130_fd_sc_hd__nor2_1 _42820_ (.A(_15678_),
    .B(_15016_),
    .Y(_15680_));
 sky130_fd_sc_hd__nand2_1 _42821_ (.A(_15011_),
    .B(_15017_),
    .Y(_15681_));
 sky130_fd_sc_hd__o211a_1 _42822_ (.A1(_12224_),
    .A2(_14439_),
    .B1(_15014_),
    .C1(_15681_),
    .X(_15682_));
 sky130_fd_sc_hd__or3_1 _42823_ (.A(_12226_),
    .B(_14443_),
    .C(_15017_),
    .X(_15683_));
 sky130_fd_sc_hd__or2b_1 _42824_ (.A(_15022_),
    .B_N(_15683_),
    .X(_15684_));
 sky130_fd_sc_hd__or3_1 _42825_ (.A(_15680_),
    .B(_15682_),
    .C(_15684_),
    .X(_15685_));
 sky130_fd_sc_hd__o21ai_1 _42826_ (.A1(_15680_),
    .A2(_15682_),
    .B1(_15684_),
    .Y(_15686_));
 sky130_fd_sc_hd__nor2_1 _42827_ (.A(_12224_),
    .B(_15021_),
    .Y(_15687_));
 sky130_fd_sc_hd__and3_1 _42828_ (.A(_15685_),
    .B(_15686_),
    .C(_15687_),
    .X(_15688_));
 sky130_fd_sc_hd__o2bb2a_1 _42829_ (.A1_N(_15685_),
    .A2_N(_15686_),
    .B1(_12224_),
    .B2(_15021_),
    .X(_15689_));
 sky130_fd_sc_hd__o211a_1 _42830_ (.A1(_15688_),
    .A2(_15689_),
    .B1(_15024_),
    .C1(_15027_),
    .X(_15691_));
 sky130_fd_sc_hd__a211oi_1 _42831_ (.A1(_15024_),
    .A2(_15027_),
    .B1(_15688_),
    .C1(_15689_),
    .Y(_15692_));
 sky130_fd_sc_hd__nor2_1 _42832_ (.A(_15691_),
    .B(_15692_),
    .Y(_15693_));
 sky130_fd_sc_hd__a21oi_1 _42833_ (.A1(_15033_),
    .A2(_15032_),
    .B1(_15029_),
    .Y(_15694_));
 sky130_fd_sc_hd__xnor2_1 _42834_ (.A(_15693_),
    .B(_15694_),
    .Y(_15695_));
 sky130_fd_sc_hd__a21o_1 _42835_ (.A1(_15676_),
    .A2(_15677_),
    .B1(_15695_),
    .X(_15696_));
 sky130_fd_sc_hd__nand3_2 _42836_ (.A(_15676_),
    .B(_15677_),
    .C(_15695_),
    .Y(_15697_));
 sky130_fd_sc_hd__inv_2 _42837_ (.A(_15054_),
    .Y(_15698_));
 sky130_fd_sc_hd__a211o_1 _42838_ (.A1(_14486_),
    .A2(_14487_),
    .B1(_15052_),
    .C1(_14484_),
    .X(_15699_));
 sky130_fd_sc_hd__a21o_1 _42839_ (.A1(_14470_),
    .A2(_15043_),
    .B1(_15038_),
    .X(_15700_));
 sky130_fd_sc_hd__a22oi_2 _42840_ (.A1(_14462_),
    .A2(_15041_),
    .B1(_15040_),
    .B2(_15700_),
    .Y(_15702_));
 sky130_fd_sc_hd__o32a_1 _42841_ (.A1(_07351_),
    .A2(_15050_),
    .A3(_15048_),
    .B1(_15047_),
    .B2(_15046_),
    .X(_15703_));
 sky130_fd_sc_hd__o21ai_1 _42842_ (.A1(_07333_),
    .A2(_15702_),
    .B1(_15703_),
    .Y(_15704_));
 sky130_fd_sc_hd__buf_1 _42843_ (.A(_14462_),
    .X(_15705_));
 sky130_fd_sc_hd__buf_1 _42844_ (.A(_13667_),
    .X(_15706_));
 sky130_fd_sc_hd__buf_1 _42845_ (.A(_11049_),
    .X(_15707_));
 sky130_fd_sc_hd__a311o_1 _42846_ (.A1(_15705_),
    .A2(_15706_),
    .A3(_15707_),
    .B1(_15702_),
    .C1(_15703_),
    .X(_15708_));
 sky130_fd_sc_hd__and2_1 _42847_ (.A(_15704_),
    .B(_15708_),
    .X(_15709_));
 sky130_fd_sc_hd__a21o_1 _42848_ (.A1(_15698_),
    .A2(_15699_),
    .B1(_15709_),
    .X(_15710_));
 sky130_fd_sc_hd__o211ai_2 _42849_ (.A1(_15052_),
    .A2(_15055_),
    .B1(_15709_),
    .C1(_15698_),
    .Y(_15711_));
 sky130_fd_sc_hd__and2_1 _42850_ (.A(_15710_),
    .B(_15711_),
    .X(_15713_));
 sky130_fd_sc_hd__a21oi_1 _42851_ (.A1(_15696_),
    .A2(_15697_),
    .B1(_15713_),
    .Y(_15714_));
 sky130_fd_sc_hd__and3_1 _42852_ (.A(_15713_),
    .B(_15696_),
    .C(_15697_),
    .X(_15715_));
 sky130_fd_sc_hd__or2_1 _42853_ (.A(_15714_),
    .B(_15715_),
    .X(_15716_));
 sky130_fd_sc_hd__a21o_1 _42854_ (.A1(_15659_),
    .A2(_15662_),
    .B1(_15716_),
    .X(_15717_));
 sky130_fd_sc_hd__nand3_2 _42855_ (.A(_15659_),
    .B(_15662_),
    .C(_15716_),
    .Y(_15718_));
 sky130_fd_sc_hd__a22oi_2 _42856_ (.A1(_15063_),
    .A2(_15061_),
    .B1(_15717_),
    .B2(_15718_),
    .Y(_15719_));
 sky130_fd_sc_hd__a31o_1 _42857_ (.A1(_15131_),
    .A2(_15085_),
    .A3(_15082_),
    .B1(_15129_),
    .X(_15720_));
 sky130_fd_sc_hd__o21ai_2 _42858_ (.A1(_15035_),
    .A2(_15058_),
    .B1(_15036_),
    .Y(_15721_));
 sky130_fd_sc_hd__nor2_1 _42859_ (.A(_15071_),
    .B(_15073_),
    .Y(_15722_));
 sky130_fd_sc_hd__o32a_1 _42860_ (.A1(_15071_),
    .A2(_07084_),
    .A3(_07080_),
    .B1(_15722_),
    .B2(_08417_),
    .X(_15724_));
 sky130_fd_sc_hd__a21oi_1 _42861_ (.A1(_15080_),
    .A2(_15085_),
    .B1(_15724_),
    .Y(_15725_));
 sky130_fd_sc_hd__o211a_1 _42862_ (.A1(_15078_),
    .A2(_15079_),
    .B1(_15724_),
    .C1(_15085_),
    .X(_15726_));
 sky130_fd_sc_hd__or2_1 _42863_ (.A(_15725_),
    .B(_15726_),
    .X(_15727_));
 sky130_fd_sc_hd__a21bo_1 _42864_ (.A1(_15094_),
    .A2(_15088_),
    .B1_N(_15093_),
    .X(_15728_));
 sky130_fd_sc_hd__xnor2_1 _42865_ (.A(_15087_),
    .B(_15090_),
    .Y(_15729_));
 sky130_fd_sc_hd__nand2_1 _42866_ (.A(_15728_),
    .B(_15729_),
    .Y(_15730_));
 sky130_fd_sc_hd__or2_1 _42867_ (.A(_15729_),
    .B(_15728_),
    .X(_15731_));
 sky130_fd_sc_hd__nand2_1 _42868_ (.A(_15730_),
    .B(_15731_),
    .Y(_15732_));
 sky130_fd_sc_hd__a21o_1 _42869_ (.A1(_15098_),
    .A2(_15101_),
    .B1(_15732_),
    .X(_15733_));
 sky130_fd_sc_hd__nand3_1 _42870_ (.A(_15098_),
    .B(_15101_),
    .C(_15732_),
    .Y(_15735_));
 sky130_fd_sc_hd__buf_1 _42871_ (.A(_14312_),
    .X(_15736_));
 sky130_fd_sc_hd__nor2_1 _42872_ (.A(_15736_),
    .B(_15109_),
    .Y(_15737_));
 sky130_fd_sc_hd__nand2_1 _42873_ (.A(_15736_),
    .B(_15110_),
    .Y(_15738_));
 sky130_fd_sc_hd__o211a_1 _42874_ (.A1(_14319_),
    .A2(_14314_),
    .B1(_15114_),
    .C1(_15738_),
    .X(_15739_));
 sky130_fd_sc_hd__or3_1 _42875_ (.A(_10045_),
    .B(_14316_),
    .C(_15110_),
    .X(_15740_));
 sky130_fd_sc_hd__or2b_1 _42876_ (.A(_15116_),
    .B_N(_15740_),
    .X(_15741_));
 sky130_fd_sc_hd__or3_1 _42877_ (.A(_15737_),
    .B(_15739_),
    .C(_15741_),
    .X(_15742_));
 sky130_fd_sc_hd__o21ai_1 _42878_ (.A1(_15737_),
    .A2(_15739_),
    .B1(_15741_),
    .Y(_15743_));
 sky130_fd_sc_hd__and3b_1 _42879_ (.A_N(_15114_),
    .B(_15113_),
    .C(_14310_),
    .X(_15744_));
 sky130_fd_sc_hd__and3_1 _42880_ (.A(_15742_),
    .B(_15743_),
    .C(_15744_),
    .X(_15746_));
 sky130_fd_sc_hd__a21oi_1 _42881_ (.A1(_15742_),
    .A2(_15743_),
    .B1(_15744_),
    .Y(_15747_));
 sky130_fd_sc_hd__a211oi_1 _42882_ (.A1(_15118_),
    .A2(_15122_),
    .B1(_15746_),
    .C1(_15747_),
    .Y(_15748_));
 sky130_fd_sc_hd__o211a_1 _42883_ (.A1(_15746_),
    .A2(_15747_),
    .B1(_15118_),
    .C1(_15122_),
    .X(_15749_));
 sky130_fd_sc_hd__nor2_1 _42884_ (.A(_15748_),
    .B(_15749_),
    .Y(_15750_));
 sky130_fd_sc_hd__a21oi_1 _42885_ (.A1(_15104_),
    .A2(_15126_),
    .B1(_15124_),
    .Y(_15751_));
 sky130_fd_sc_hd__xnor2_1 _42886_ (.A(_15750_),
    .B(_15751_),
    .Y(_15752_));
 sky130_fd_sc_hd__a21oi_1 _42887_ (.A1(_15733_),
    .A2(_15735_),
    .B1(_15752_),
    .Y(_15753_));
 sky130_fd_sc_hd__nand3_1 _42888_ (.A(_15752_),
    .B(_15733_),
    .C(_15735_),
    .Y(_15754_));
 sky130_fd_sc_hd__and2b_1 _42889_ (.A_N(_15753_),
    .B(_15754_),
    .X(_15755_));
 sky130_fd_sc_hd__xnor2_1 _42890_ (.A(_15727_),
    .B(_15755_),
    .Y(_15757_));
 sky130_fd_sc_hd__xor2_1 _42891_ (.A(net78),
    .B(_15757_),
    .X(_15758_));
 sky130_fd_sc_hd__xor2_2 _42892_ (.A(_15720_),
    .B(_15758_),
    .X(_15759_));
 sky130_fd_sc_hd__nand4_4 _42893_ (.A(_15063_),
    .B(_15061_),
    .C(_15717_),
    .D(_15718_),
    .Y(_15760_));
 sky130_fd_sc_hd__and3b_1 _42894_ (.A_N(net65),
    .B(_15759_),
    .C(_15760_),
    .X(_15761_));
 sky130_fd_sc_hd__inv_2 _42895_ (.A(net65),
    .Y(_15762_));
 sky130_fd_sc_hd__a21oi_1 _42896_ (.A1(_15762_),
    .A2(_15760_),
    .B1(_15759_),
    .Y(_15763_));
 sky130_fd_sc_hd__o21a_1 _42897_ (.A1(net67),
    .A2(_15138_),
    .B1(net68),
    .X(_15764_));
 sky130_fd_sc_hd__o21a_1 _42898_ (.A1(_15761_),
    .A2(_15763_),
    .B1(_15764_),
    .X(_15765_));
 sky130_fd_sc_hd__o32a_2 _42899_ (.A1(_14905_),
    .A2(_14902_),
    .A3(_14904_),
    .B1(_14906_),
    .B2(_14934_),
    .X(_15766_));
 sky130_fd_sc_hd__or2_1 _42900_ (.A(_15069_),
    .B(_15137_),
    .X(_15768_));
 sky130_fd_sc_hd__clkbuf_2 _42901_ (.A(_14903_),
    .X(_15769_));
 sky130_fd_sc_hd__a21boi_2 _42902_ (.A1(_14900_),
    .A2(_15769_),
    .B1_N(_14901_),
    .Y(_15770_));
 sky130_fd_sc_hd__clkbuf_2 _42903_ (.A(_14550_),
    .X(_15771_));
 sky130_fd_sc_hd__a21o_1 _42904_ (.A1(_02223_),
    .A2(_05508_),
    .B1(_15771_),
    .X(_15772_));
 sky130_fd_sc_hd__a2bb2o_1 _42905_ (.A1_N(_14556_),
    .A2_N(_14895_),
    .B1(_15772_),
    .B2(_05501_),
    .X(_15773_));
 sky130_fd_sc_hd__a21o_1 _42906_ (.A1(_14893_),
    .A2(_14894_),
    .B1(_15773_),
    .X(_15774_));
 sky130_fd_sc_hd__o311a_1 _42907_ (.A1(_13325_),
    .A2(_13331_),
    .A3(_13330_),
    .B1(_14557_),
    .C1(_14896_),
    .X(_15775_));
 sky130_fd_sc_hd__clkbuf_2 _42908_ (.A(_13336_),
    .X(_15776_));
 sky130_fd_sc_hd__o211ai_1 _42909_ (.A1(_11337_),
    .A2(_07013_),
    .B1(_12584_),
    .C1(_15776_),
    .Y(_15777_));
 sky130_fd_sc_hd__or3b_1 _42910_ (.A(_14876_),
    .B(_14878_),
    .C_N(_13337_),
    .X(_15779_));
 sky130_fd_sc_hd__a21oi_2 _42911_ (.A1(_15777_),
    .A2(_15779_),
    .B1(_14572_),
    .Y(_15780_));
 sky130_fd_sc_hd__a21boi_2 _42912_ (.A1(_15776_),
    .A2(_14881_),
    .B1_N(_14880_),
    .Y(_15781_));
 sky130_fd_sc_hd__a21o_1 _42913_ (.A1(_14572_),
    .A2(_15779_),
    .B1(_15781_),
    .X(_15782_));
 sky130_fd_sc_hd__and2_1 _42914_ (.A(_14572_),
    .B(_15779_),
    .X(_15783_));
 sky130_fd_sc_hd__o21ai_1 _42915_ (.A1(_15783_),
    .A2(_15780_),
    .B1(_15781_),
    .Y(_15784_));
 sky130_fd_sc_hd__o21a_1 _42916_ (.A1(_15780_),
    .A2(_15782_),
    .B1(_15784_),
    .X(_15785_));
 sky130_fd_sc_hd__a21boi_1 _42917_ (.A1(_14872_),
    .A2(_14884_),
    .B1_N(_14885_),
    .Y(_15786_));
 sky130_fd_sc_hd__xor2_1 _42918_ (.A(_15785_),
    .B(_15786_),
    .X(_15787_));
 sky130_fd_sc_hd__o21ai_1 _42919_ (.A1(_15774_),
    .A2(_15775_),
    .B1(_15787_),
    .Y(_15788_));
 sky130_fd_sc_hd__or3_1 _42920_ (.A(_15775_),
    .B(_15774_),
    .C(_15787_),
    .X(_15790_));
 sky130_fd_sc_hd__a21oi_1 _42921_ (.A1(_15788_),
    .A2(_15790_),
    .B1(_14903_),
    .Y(_15791_));
 sky130_fd_sc_hd__o311a_1 _42922_ (.A1(_15775_),
    .A2(_15774_),
    .A3(_15787_),
    .B1(_14903_),
    .C1(_15788_),
    .X(_15792_));
 sky130_fd_sc_hd__or2_1 _42923_ (.A(_15791_),
    .B(_15792_),
    .X(_15793_));
 sky130_fd_sc_hd__xnor2_2 _42924_ (.A(_15770_),
    .B(_15793_),
    .Y(_15794_));
 sky130_fd_sc_hd__o21ai_1 _42925_ (.A1(_10244_),
    .A2(_13366_),
    .B1(_10245_),
    .Y(_15795_));
 sky130_fd_sc_hd__a32o_1 _42926_ (.A1(_14518_),
    .A2(_14923_),
    .A3(_14924_),
    .B1(_15795_),
    .B2(_14512_),
    .X(_15796_));
 sky130_fd_sc_hd__a211o_2 _42927_ (.A1(_10245_),
    .A2(_14511_),
    .B1(_15796_),
    .C1(_14928_),
    .X(_15797_));
 sky130_fd_sc_hd__o31ai_2 _42928_ (.A1(_11413_),
    .A2(_12513_),
    .A3(_11414_),
    .B1(_11423_),
    .Y(_15798_));
 sky130_fd_sc_hd__nor2_1 _42929_ (.A(_14544_),
    .B(_14916_),
    .Y(_15799_));
 sky130_fd_sc_hd__o21a_1 _42930_ (.A1(_14913_),
    .A2(_14916_),
    .B1(_14544_),
    .X(_15801_));
 sky130_fd_sc_hd__a21oi_2 _42931_ (.A1(_15798_),
    .A2(_15799_),
    .B1(_15801_),
    .Y(_15802_));
 sky130_fd_sc_hd__xor2_4 _42932_ (.A(_15797_),
    .B(_15802_),
    .X(_15803_));
 sky130_fd_sc_hd__xnor2_2 _42933_ (.A(_15794_),
    .B(_15803_),
    .Y(_15804_));
 sky130_fd_sc_hd__a21o_1 _42934_ (.A1(_15136_),
    .A2(_15768_),
    .B1(_15804_),
    .X(_15805_));
 sky130_fd_sc_hd__o211ai_1 _42935_ (.A1(_15137_),
    .A2(_15069_),
    .B1(_15136_),
    .C1(_15804_),
    .Y(_15806_));
 sky130_fd_sc_hd__nand2_1 _42936_ (.A(_15805_),
    .B(_15806_),
    .Y(_15807_));
 sky130_fd_sc_hd__xnor2_1 _42937_ (.A(_15766_),
    .B(_15807_),
    .Y(_15808_));
 sky130_fd_sc_hd__or2_1 _42938_ (.A(_15765_),
    .B(_15808_),
    .X(_15809_));
 sky130_fd_sc_hd__or3_2 _42939_ (.A(_15764_),
    .B(_15761_),
    .C(_15763_),
    .X(_15810_));
 sky130_fd_sc_hd__nand2b_1 _42940_ (.A_N(_15809_),
    .B(_15810_),
    .Y(_15812_));
 sky130_fd_sc_hd__inv_2 _42941_ (.A(_15765_),
    .Y(_15813_));
 sky130_fd_sc_hd__a21bo_1 _42942_ (.A1(_15810_),
    .A2(_15813_),
    .B1_N(_15808_),
    .X(_15814_));
 sky130_fd_sc_hd__o21a_1 _42943_ (.A1(_14941_),
    .A2(_15145_),
    .B1(_15144_),
    .X(_15815_));
 sky130_fd_sc_hd__a21boi_1 _42944_ (.A1(_15812_),
    .A2(_15814_),
    .B1_N(_15815_),
    .Y(_15816_));
 sky130_fd_sc_hd__nand3b_1 _42945_ (.A_N(_15815_),
    .B(_15812_),
    .C(_15814_),
    .Y(_15817_));
 sky130_fd_sc_hd__nand2b_1 _42946_ (.A_N(_15816_),
    .B(_15817_),
    .Y(_15818_));
 sky130_fd_sc_hd__nand2_1 _42947_ (.A(_15629_),
    .B(_15818_),
    .Y(_15819_));
 sky130_fd_sc_hd__or2_1 _42948_ (.A(_15818_),
    .B(_15629_),
    .X(_15820_));
 sky130_fd_sc_hd__and4_2 _42949_ (.A(_15149_),
    .B(_15153_),
    .C(_15819_),
    .D(_15820_),
    .X(_15821_));
 sky130_fd_sc_hd__a22oi_4 _42950_ (.A1(_15149_),
    .A2(_15153_),
    .B1(_15819_),
    .B2(_15820_),
    .Y(_15823_));
 sky130_fd_sc_hd__o211a_1 _42951_ (.A1(_15422_),
    .A2(_15424_),
    .B1(_15425_),
    .C1(_15434_),
    .X(_15824_));
 sky130_fd_sc_hd__a21boi_2 _42952_ (.A1(_15287_),
    .A2(_15357_),
    .B1_N(_15292_),
    .Y(_15825_));
 sky130_fd_sc_hd__a21oi_1 _42953_ (.A1(_15202_),
    .A2(_15203_),
    .B1(_15204_),
    .Y(_15826_));
 sky130_fd_sc_hd__a21oi_1 _42954_ (.A1(_13962_),
    .A2(_15177_),
    .B1(_15176_),
    .Y(_15827_));
 sky130_fd_sc_hd__o21ai_1 _42955_ (.A1(_12952_),
    .A2(_15827_),
    .B1(_15178_),
    .Y(_15828_));
 sky130_fd_sc_hd__a21o_1 _42956_ (.A1(_12925_),
    .A2(_13941_),
    .B1(_15179_),
    .X(_15829_));
 sky130_fd_sc_hd__or3_1 _42957_ (.A(_13968_),
    .B(_12962_),
    .C(_15175_),
    .X(_15830_));
 sky130_fd_sc_hd__o21ai_2 _42958_ (.A1(_12952_),
    .A2(_15829_),
    .B1(_15830_),
    .Y(_15831_));
 sky130_fd_sc_hd__and2_2 _42959_ (.A(_15828_),
    .B(_15831_),
    .X(_15832_));
 sky130_fd_sc_hd__a21oi_2 _42960_ (.A1(_13974_),
    .A2(_15181_),
    .B1(_15831_),
    .Y(_15834_));
 sky130_fd_sc_hd__a22oi_4 _42961_ (.A1(_15182_),
    .A2(_15195_),
    .B1(_15190_),
    .B2(_13982_),
    .Y(_15835_));
 sky130_fd_sc_hd__o31ai_4 _42962_ (.A1(_15832_),
    .A2(_15834_),
    .A3(_15835_),
    .B1(_15184_),
    .Y(_15836_));
 sky130_fd_sc_hd__o211a_1 _42963_ (.A1(_12956_),
    .A2(_15826_),
    .B1(_15205_),
    .C1(_15836_),
    .X(_15837_));
 sky130_fd_sc_hd__nand2_1 _42964_ (.A(_15201_),
    .B(_15206_),
    .Y(_15838_));
 sky130_fd_sc_hd__a21oi_2 _42965_ (.A1(_15209_),
    .A2(_15838_),
    .B1(_15836_),
    .Y(_15839_));
 sky130_fd_sc_hd__and2_1 _42966_ (.A(_12994_),
    .B(_15217_),
    .X(_15840_));
 sky130_fd_sc_hd__or2b_1 _42967_ (.A(_14013_),
    .B_N(_14007_),
    .X(_15841_));
 sky130_fd_sc_hd__clkbuf_2 _42968_ (.A(_15223_),
    .X(_15842_));
 sky130_fd_sc_hd__nor2_1 _42969_ (.A(_15216_),
    .B(_15842_),
    .Y(_15843_));
 sky130_fd_sc_hd__a31o_1 _42970_ (.A1(_13014_),
    .A2(_15841_),
    .A3(_15842_),
    .B1(_15843_),
    .X(_15845_));
 sky130_fd_sc_hd__or3b_1 _42971_ (.A(_14010_),
    .B(_15840_),
    .C_N(_15845_),
    .X(_15846_));
 sky130_fd_sc_hd__a311o_1 _42972_ (.A1(_15842_),
    .A2(_13014_),
    .A3(_15841_),
    .B1(_15843_),
    .C1(_15221_),
    .X(_15847_));
 sky130_fd_sc_hd__nand2_1 _42973_ (.A(_15846_),
    .B(_15847_),
    .Y(_15848_));
 sky130_fd_sc_hd__a32o_1 _42974_ (.A1(_12994_),
    .A2(_15217_),
    .A3(_10648_),
    .B1(_15222_),
    .B2(_15225_),
    .X(_15849_));
 sky130_fd_sc_hd__nor2_1 _42975_ (.A(_15848_),
    .B(_15849_),
    .Y(_15850_));
 sky130_fd_sc_hd__and2_1 _42976_ (.A(_15848_),
    .B(_15849_),
    .X(_15851_));
 sky130_fd_sc_hd__nor2_1 _42977_ (.A(_15850_),
    .B(_15851_),
    .Y(_15852_));
 sky130_fd_sc_hd__inv_2 _42978_ (.A(_15852_),
    .Y(_15853_));
 sky130_fd_sc_hd__o21ai_2 _42979_ (.A1(_15837_),
    .A2(_15839_),
    .B1(_15853_),
    .Y(_15854_));
 sky130_fd_sc_hd__a21o_1 _42980_ (.A1(_15209_),
    .A2(_15838_),
    .B1(_15836_),
    .X(_15856_));
 sky130_fd_sc_hd__nand3b_2 _42981_ (.A_N(_15837_),
    .B(_15856_),
    .C(_15852_),
    .Y(_15857_));
 sky130_fd_sc_hd__nand2_1 _42982_ (.A(_15854_),
    .B(_15857_),
    .Y(_15858_));
 sky130_fd_sc_hd__a21boi_1 _42983_ (.A1(_15215_),
    .A2(_15235_),
    .B1_N(_15211_),
    .Y(_15859_));
 sky130_fd_sc_hd__nand2_1 _42984_ (.A(_15858_),
    .B(_15859_),
    .Y(_15860_));
 sky130_fd_sc_hd__inv_2 _42985_ (.A(_15235_),
    .Y(_15861_));
 sky130_fd_sc_hd__a21oi_1 _42986_ (.A1(_15208_),
    .A2(_15210_),
    .B1(_15173_),
    .Y(_15862_));
 sky130_fd_sc_hd__o21ai_1 _42987_ (.A1(_15861_),
    .A2(_15862_),
    .B1(_15211_),
    .Y(_15863_));
 sky130_fd_sc_hd__nand3_1 _42988_ (.A(_15854_),
    .B(_15857_),
    .C(_15863_),
    .Y(_15864_));
 sky130_fd_sc_hd__clkbuf_2 _42989_ (.A(_15864_),
    .X(_15865_));
 sky130_fd_sc_hd__clkbuf_2 _42990_ (.A(_13060_),
    .X(_15867_));
 sky130_fd_sc_hd__buf_1 _42991_ (.A(_13041_),
    .X(_15868_));
 sky130_fd_sc_hd__and3_1 _42992_ (.A(_07692_),
    .B(_15257_),
    .C(_13041_),
    .X(_15869_));
 sky130_fd_sc_hd__a21oi_1 _42993_ (.A1(_07696_),
    .A2(_15868_),
    .B1(_15842_),
    .Y(_15870_));
 sky130_fd_sc_hd__and3_1 _42994_ (.A(_07696_),
    .B(_15868_),
    .C(_15223_),
    .X(_15871_));
 sky130_fd_sc_hd__a2111oi_1 _42995_ (.A1(_15868_),
    .A2(_15260_),
    .B1(_15869_),
    .C1(_15870_),
    .D1(_15871_),
    .Y(_15872_));
 sky130_fd_sc_hd__and3_1 _42996_ (.A(_07690_),
    .B(_14060_),
    .C(_15868_),
    .X(_15873_));
 sky130_fd_sc_hd__o22a_2 _42997_ (.A1(_15870_),
    .A2(_15871_),
    .B1(_15873_),
    .B2(_15869_),
    .X(_15874_));
 sky130_fd_sc_hd__a311oi_4 _42998_ (.A1(_11752_),
    .A2(_13045_),
    .A3(_15867_),
    .B1(net174),
    .C1(_15874_),
    .Y(_15875_));
 sky130_fd_sc_hd__o211a_1 _42999_ (.A1(_15872_),
    .A2(_15874_),
    .B1(_15867_),
    .C1(_06400_),
    .X(_15876_));
 sky130_fd_sc_hd__buf_1 _43000_ (.A(_13008_),
    .X(_15878_));
 sky130_fd_sc_hd__o21a_1 _43001_ (.A1(_15878_),
    .A2(_14043_),
    .B1(_15216_),
    .X(_15879_));
 sky130_fd_sc_hd__nor3_1 _43002_ (.A(_15216_),
    .B(_15878_),
    .C(_14043_),
    .Y(_15880_));
 sky130_fd_sc_hd__clkbuf_2 _43003_ (.A(_15878_),
    .X(_15881_));
 sky130_fd_sc_hd__a2111oi_1 _43004_ (.A1(_15246_),
    .A2(_14019_),
    .B1(_15879_),
    .C1(_15880_),
    .D1(_15881_),
    .Y(_15882_));
 sky130_fd_sc_hd__o21a_1 _43005_ (.A1(_15879_),
    .A2(_15880_),
    .B1(_15247_),
    .X(_15883_));
 sky130_fd_sc_hd__o21ai_1 _43006_ (.A1(_14045_),
    .A2(_15248_),
    .B1(_15249_),
    .Y(_15884_));
 sky130_fd_sc_hd__or3_1 _43007_ (.A(net162),
    .B(_15883_),
    .C(_15884_),
    .X(_15885_));
 sky130_fd_sc_hd__o21ai_2 _43008_ (.A1(net160),
    .A2(_15883_),
    .B1(_15884_),
    .Y(_15886_));
 sky130_fd_sc_hd__or4bb_1 _43009_ (.A(_15875_),
    .B(_15876_),
    .C_N(_15885_),
    .D_N(_15886_),
    .X(_15887_));
 sky130_fd_sc_hd__inv_2 _43010_ (.A(_15887_),
    .Y(_15889_));
 sky130_fd_sc_hd__a2bb2oi_2 _43011_ (.A1_N(_15875_),
    .A2_N(_15876_),
    .B1(_15885_),
    .B2(_15886_),
    .Y(_15890_));
 sky130_fd_sc_hd__a211o_1 _43012_ (.A1(_15227_),
    .A2(_15231_),
    .B1(_15889_),
    .C1(_15890_),
    .X(_15891_));
 sky130_fd_sc_hd__o221ai_4 _43013_ (.A1(_15230_),
    .A2(_15220_),
    .B1(_15890_),
    .B2(_15889_),
    .C1(_15227_),
    .Y(_15892_));
 sky130_fd_sc_hd__a31o_1 _43014_ (.A1(_15256_),
    .A2(_15271_),
    .A3(_15272_),
    .B1(_15254_),
    .X(_15893_));
 sky130_fd_sc_hd__a21boi_2 _43015_ (.A1(_15891_),
    .A2(_15892_),
    .B1_N(_15893_),
    .Y(_15894_));
 sky130_fd_sc_hd__and4bb_1 _43016_ (.A_N(_15254_),
    .B_N(_15274_),
    .C(_15891_),
    .D(_15892_),
    .X(_15895_));
 sky130_fd_sc_hd__nor2_2 _43017_ (.A(_15894_),
    .B(_15895_),
    .Y(_15896_));
 sky130_fd_sc_hd__nand3_1 _43018_ (.A(_15860_),
    .B(_15865_),
    .C(_15896_),
    .Y(_15897_));
 sky130_fd_sc_hd__o2bb2ai_1 _43019_ (.A1_N(_15860_),
    .A2_N(_15864_),
    .B1(_15894_),
    .B2(_15895_),
    .Y(_15898_));
 sky130_fd_sc_hd__nand4_4 _43020_ (.A(_15285_),
    .B(_15290_),
    .C(_15897_),
    .D(_15898_),
    .Y(_15900_));
 sky130_fd_sc_hd__o21ai_1 _43021_ (.A1(_15282_),
    .A2(_15242_),
    .B1(_15285_),
    .Y(_15901_));
 sky130_fd_sc_hd__o211ai_1 _43022_ (.A1(_15894_),
    .A2(_15895_),
    .B1(_15860_),
    .C1(_15865_),
    .Y(_15902_));
 sky130_fd_sc_hd__a21bo_1 _43023_ (.A1(_15860_),
    .A2(_15864_),
    .B1_N(_15896_),
    .X(_15903_));
 sky130_fd_sc_hd__nand3_2 _43024_ (.A(_15901_),
    .B(_15902_),
    .C(_15903_),
    .Y(_15904_));
 sky130_fd_sc_hd__a21oi_2 _43025_ (.A1(_15323_),
    .A2(_15349_),
    .B1(_15347_),
    .Y(_15905_));
 sky130_fd_sc_hd__a21oi_1 _43026_ (.A1(_15325_),
    .A2(_15343_),
    .B1(_15346_),
    .Y(_15906_));
 sky130_fd_sc_hd__or4b_1 _43027_ (.A(_15260_),
    .B(_14062_),
    .C(_15869_),
    .D_N(_15259_),
    .X(_15907_));
 sky130_fd_sc_hd__and3_1 _43028_ (.A(_06432_),
    .B(_13050_),
    .C(_12029_),
    .X(_15908_));
 sky130_fd_sc_hd__a21oi_2 _43029_ (.A1(_13161_),
    .A2(_12029_),
    .B1(_13051_),
    .Y(_15909_));
 sky130_fd_sc_hd__or4_2 _43030_ (.A(_15266_),
    .B(_15269_),
    .C(_15908_),
    .D(_15909_),
    .X(_15911_));
 sky130_fd_sc_hd__o22ai_4 _43031_ (.A1(_15266_),
    .A2(_15269_),
    .B1(_15908_),
    .B2(_15909_),
    .Y(_15912_));
 sky130_fd_sc_hd__a21o_1 _43032_ (.A1(_15911_),
    .A2(_15912_),
    .B1(_15335_),
    .X(_15913_));
 sky130_fd_sc_hd__o2111ai_4 _43033_ (.A1(_15331_),
    .A2(_15333_),
    .B1(_15912_),
    .C1(_13060_),
    .D1(_15911_),
    .Y(_15914_));
 sky130_fd_sc_hd__nand2_1 _43034_ (.A(_15913_),
    .B(_15914_),
    .Y(_15915_));
 sky130_fd_sc_hd__a21oi_1 _43035_ (.A1(_15907_),
    .A2(_15272_),
    .B1(_15915_),
    .Y(_15916_));
 sky130_fd_sc_hd__o311a_1 _43036_ (.A1(_15261_),
    .A2(_15269_),
    .A3(_15270_),
    .B1(_15915_),
    .C1(_15907_),
    .X(_15917_));
 sky130_fd_sc_hd__nor2_1 _43037_ (.A(_15916_),
    .B(_15917_),
    .Y(_15918_));
 sky130_fd_sc_hd__o21a_1 _43038_ (.A1(_15337_),
    .A2(_15341_),
    .B1(_15918_),
    .X(_15919_));
 sky130_fd_sc_hd__or3_1 _43039_ (.A(_15337_),
    .B(_15341_),
    .C(_15918_),
    .X(_15920_));
 sky130_fd_sc_hd__inv_2 _43040_ (.A(_15920_),
    .Y(_15922_));
 sky130_fd_sc_hd__or3_2 _43041_ (.A(_15906_),
    .B(_15919_),
    .C(_15922_),
    .X(_15923_));
 sky130_fd_sc_hd__o21ai_2 _43042_ (.A1(_13113_),
    .A2(_15307_),
    .B1(_15305_),
    .Y(_15924_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43043_ (.A(_15302_),
    .X(_15925_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43044_ (.A(_11968_),
    .X(_15926_));
 sky130_fd_sc_hd__o21a_1 _43045_ (.A1(_12003_),
    .A2(_15302_),
    .B1(_12013_),
    .X(_15927_));
 sky130_fd_sc_hd__and3b_1 _43046_ (.A_N(_12003_),
    .B(_12015_),
    .C(_13134_),
    .X(_15928_));
 sky130_fd_sc_hd__or2_1 _43047_ (.A(_15927_),
    .B(_15928_),
    .X(_15929_));
 sky130_fd_sc_hd__nand2_1 _43048_ (.A(_13161_),
    .B(_12029_),
    .Y(_15930_));
 sky130_fd_sc_hd__o2bb2a_1 _43049_ (.A1_N(_11968_),
    .A2_N(_15930_),
    .B1(_15330_),
    .B2(_15908_),
    .X(_15931_));
 sky130_fd_sc_hd__and3_1 _43050_ (.A(_13135_),
    .B(_15311_),
    .C(_15931_),
    .X(_15933_));
 sky130_fd_sc_hd__nor2_2 _43051_ (.A(_15931_),
    .B(_15310_),
    .Y(_15934_));
 sky130_fd_sc_hd__a2111oi_2 _43052_ (.A1(_15925_),
    .A2(_15926_),
    .B1(_15929_),
    .C1(_15933_),
    .D1(_15934_),
    .Y(_15935_));
 sky130_fd_sc_hd__a2bb2o_1 _43053_ (.A1_N(_15931_),
    .A2_N(_15310_),
    .B1(_11968_),
    .B2(_15925_),
    .X(_15936_));
 sky130_fd_sc_hd__o22a_1 _43054_ (.A1(_15927_),
    .A2(_15928_),
    .B1(_15933_),
    .B2(_15936_),
    .X(_15937_));
 sky130_fd_sc_hd__a211o_1 _43055_ (.A1(_15312_),
    .A2(_15315_),
    .B1(_15935_),
    .C1(_15937_),
    .X(_15938_));
 sky130_fd_sc_hd__o211ai_1 _43056_ (.A1(_15935_),
    .A2(_15937_),
    .B1(_15312_),
    .C1(_15315_),
    .Y(_15939_));
 sky130_fd_sc_hd__nand2_1 _43057_ (.A(_15938_),
    .B(_15939_),
    .Y(_15940_));
 sky130_fd_sc_hd__or2_1 _43058_ (.A(_15924_),
    .B(_15940_),
    .X(_15941_));
 sky130_fd_sc_hd__nand2_1 _43059_ (.A(_15924_),
    .B(_15940_),
    .Y(_15942_));
 sky130_fd_sc_hd__and2_1 _43060_ (.A(_15941_),
    .B(_15942_),
    .X(_15944_));
 sky130_fd_sc_hd__o21ai_1 _43061_ (.A1(_15919_),
    .A2(_15922_),
    .B1(_15906_),
    .Y(_15945_));
 sky130_fd_sc_hd__nand3_2 _43062_ (.A(_15923_),
    .B(_15944_),
    .C(_15945_),
    .Y(_15946_));
 sky130_fd_sc_hd__inv_2 _43063_ (.A(_15946_),
    .Y(_15947_));
 sky130_fd_sc_hd__a21oi_1 _43064_ (.A1(_15945_),
    .A2(_15923_),
    .B1(_15944_),
    .Y(_15948_));
 sky130_fd_sc_hd__o221ai_1 _43065_ (.A1(_15278_),
    .A2(_15276_),
    .B1(_15947_),
    .B2(_15948_),
    .C1(_15277_),
    .Y(_15949_));
 sky130_fd_sc_hd__o21ai_1 _43066_ (.A1(_14071_),
    .A2(_14072_),
    .B1(_15280_),
    .Y(_15950_));
 sky130_fd_sc_hd__a211o_1 _43067_ (.A1(_15277_),
    .A2(_15950_),
    .B1(_15947_),
    .C1(_15948_),
    .X(_15951_));
 sky130_fd_sc_hd__nand2_1 _43068_ (.A(_15949_),
    .B(_15951_),
    .Y(_15952_));
 sky130_fd_sc_hd__xor2_2 _43069_ (.A(_15905_),
    .B(_15952_),
    .X(_15953_));
 sky130_fd_sc_hd__a21bo_2 _43070_ (.A1(_15900_),
    .A2(_15904_),
    .B1_N(_15953_),
    .X(_15955_));
 sky130_fd_sc_hd__nand3b_4 _43071_ (.A_N(_15953_),
    .B(_15900_),
    .C(_15904_),
    .Y(_15956_));
 sky130_fd_sc_hd__nand3_2 _43072_ (.A(_15825_),
    .B(_15955_),
    .C(_15956_),
    .Y(_15957_));
 sky130_fd_sc_hd__and2b_1 _43073_ (.A_N(_15378_),
    .B(_15368_),
    .X(_15958_));
 sky130_fd_sc_hd__inv_2 _43074_ (.A(_15958_),
    .Y(_15959_));
 sky130_fd_sc_hd__a21o_1 _43075_ (.A1(_15354_),
    .A2(_15356_),
    .B1(_15352_),
    .X(_15960_));
 sky130_fd_sc_hd__a21o_1 _43076_ (.A1(_14166_),
    .A2(_15377_),
    .B1(_15376_),
    .X(_15961_));
 sky130_fd_sc_hd__a2111oi_1 _43077_ (.A1(_15294_),
    .A2(_13125_),
    .B1(_15369_),
    .C1(_14167_),
    .D1(_15300_),
    .Y(_15962_));
 sky130_fd_sc_hd__a21o_1 _43078_ (.A1(_15294_),
    .A2(_13125_),
    .B1(_15300_),
    .X(_15963_));
 sky130_fd_sc_hd__o21a_1 _43079_ (.A1(_14167_),
    .A2(_15369_),
    .B1(_15963_),
    .X(_15964_));
 sky130_fd_sc_hd__o211a_1 _43080_ (.A1(net158),
    .A2(_15964_),
    .B1(_15319_),
    .C1(_15321_),
    .X(_15966_));
 sky130_fd_sc_hd__a211oi_1 _43081_ (.A1(_15319_),
    .A2(_15321_),
    .B1(net157),
    .C1(_15964_),
    .Y(_15967_));
 sky130_fd_sc_hd__or2_1 _43082_ (.A(_15966_),
    .B(_15967_),
    .X(_15968_));
 sky130_fd_sc_hd__a211o_1 _43083_ (.A1(_14098_),
    .A2(_15371_),
    .B1(_13209_),
    .C1(_15968_),
    .X(_15969_));
 sky130_fd_sc_hd__nand2_1 _43084_ (.A(_15373_),
    .B(_15968_),
    .Y(_15970_));
 sky130_fd_sc_hd__nand2_1 _43085_ (.A(_15969_),
    .B(_15970_),
    .Y(_15971_));
 sky130_fd_sc_hd__xnor2_1 _43086_ (.A(_15961_),
    .B(_15971_),
    .Y(_15972_));
 sky130_fd_sc_hd__xnor2_1 _43087_ (.A(_15960_),
    .B(_15972_),
    .Y(_15973_));
 sky130_fd_sc_hd__nor2_1 _43088_ (.A(_15959_),
    .B(_15973_),
    .Y(_15974_));
 sky130_fd_sc_hd__and2_1 _43089_ (.A(_15959_),
    .B(_15973_),
    .X(_15975_));
 sky130_fd_sc_hd__nor2_1 _43090_ (.A(_15974_),
    .B(_15975_),
    .Y(_15977_));
 sky130_fd_sc_hd__nand2_1 _43091_ (.A(_15957_),
    .B(_15977_),
    .Y(_15978_));
 sky130_fd_sc_hd__a21oi_2 _43092_ (.A1(_15955_),
    .A2(_15956_),
    .B1(_15825_),
    .Y(_15979_));
 sky130_fd_sc_hd__nand2_1 _43093_ (.A(_15366_),
    .B(_15385_),
    .Y(_15980_));
 sky130_fd_sc_hd__nand2_1 _43094_ (.A(_15389_),
    .B(_15980_),
    .Y(_15981_));
 sky130_fd_sc_hd__a21o_1 _43095_ (.A1(_15955_),
    .A2(_15956_),
    .B1(_15825_),
    .X(_15982_));
 sky130_fd_sc_hd__a21o_1 _43096_ (.A1(_15982_),
    .A2(_15957_),
    .B1(_15977_),
    .X(_15983_));
 sky130_fd_sc_hd__o211ai_4 _43097_ (.A1(_15978_),
    .A2(_15979_),
    .B1(_15981_),
    .C1(_15983_),
    .Y(_15984_));
 sky130_fd_sc_hd__a21bo_1 _43098_ (.A1(_15982_),
    .A2(_15957_),
    .B1_N(_15977_),
    .X(_15985_));
 sky130_fd_sc_hd__nand3b_1 _43099_ (.A_N(_15977_),
    .B(_15982_),
    .C(_15957_),
    .Y(_15986_));
 sky130_fd_sc_hd__nand4_4 _43100_ (.A(_15389_),
    .B(_15980_),
    .C(_15985_),
    .D(_15986_),
    .Y(_15988_));
 sky130_fd_sc_hd__o21ai_4 _43101_ (.A1(_15367_),
    .A2(_15384_),
    .B1(_15380_),
    .Y(_15989_));
 sky130_fd_sc_hd__a21bo_1 _43102_ (.A1(_15984_),
    .A2(_15988_),
    .B1_N(_15989_),
    .X(_15990_));
 sky130_fd_sc_hd__nand3b_2 _43103_ (.A_N(_15989_),
    .B(_15984_),
    .C(_15988_),
    .Y(_15991_));
 sky130_fd_sc_hd__a31o_1 _43104_ (.A1(_15387_),
    .A2(_15388_),
    .A3(_15390_),
    .B1(_15169_),
    .X(_15992_));
 sky130_fd_sc_hd__and2_1 _43105_ (.A(_15396_),
    .B(_15992_),
    .X(_15993_));
 sky130_fd_sc_hd__a21oi_2 _43106_ (.A1(_15990_),
    .A2(_15991_),
    .B1(_15993_),
    .Y(_15994_));
 sky130_fd_sc_hd__nand4_4 _43107_ (.A(_15396_),
    .B(_15992_),
    .C(_15990_),
    .D(_15991_),
    .Y(_15995_));
 sky130_fd_sc_hd__inv_2 _43108_ (.A(_15995_),
    .Y(_15996_));
 sky130_fd_sc_hd__nor2_1 _43109_ (.A(_15994_),
    .B(_15996_),
    .Y(_15997_));
 sky130_fd_sc_hd__o21ai_1 _43110_ (.A1(_13244_),
    .A2(_13254_),
    .B1(_14199_),
    .Y(_15999_));
 sky130_fd_sc_hd__nor3b_1 _43111_ (.A(_13250_),
    .B(_14195_),
    .C_N(_14198_),
    .Y(_16000_));
 sky130_fd_sc_hd__a22oi_4 _43112_ (.A1(_14206_),
    .A2(_15999_),
    .B1(_13264_),
    .B2(net61),
    .Y(_16001_));
 sky130_fd_sc_hd__o22ai_2 _43113_ (.A1(_15400_),
    .A2(_15398_),
    .B1(_15404_),
    .B2(_16001_),
    .Y(_16002_));
 sky130_fd_sc_hd__o22a_1 _43114_ (.A1(_15398_),
    .A2(_15400_),
    .B1(_15994_),
    .B2(_15996_),
    .X(_16003_));
 sky130_fd_sc_hd__o21ai_2 _43115_ (.A1(_15409_),
    .A2(_16001_),
    .B1(_16003_),
    .Y(_16004_));
 sky130_fd_sc_hd__o21ai_2 _43116_ (.A1(_15162_),
    .A2(_15164_),
    .B1(_16004_),
    .Y(_16005_));
 sky130_fd_sc_hd__a21oi_1 _43117_ (.A1(_15997_),
    .A2(_16002_),
    .B1(_16005_),
    .Y(_16006_));
 sky130_fd_sc_hd__clkbuf_2 _43118_ (.A(_12885_),
    .X(_16007_));
 sky130_fd_sc_hd__nand2_1 _43119_ (.A(_16002_),
    .B(_15997_),
    .Y(_16008_));
 sky130_fd_sc_hd__clkbuf_2 _43120_ (.A(_15429_),
    .X(_16010_));
 sky130_fd_sc_hd__a21oi_1 _43121_ (.A1(_16004_),
    .A2(_16008_),
    .B1(_16010_),
    .Y(_16011_));
 sky130_fd_sc_hd__nor3_1 _43122_ (.A(_16006_),
    .B(_16007_),
    .C(_16011_),
    .Y(_16012_));
 sky130_fd_sc_hd__a21o_1 _43123_ (.A1(_16004_),
    .A2(_16008_),
    .B1(_15429_),
    .X(_16013_));
 sky130_fd_sc_hd__inv_2 _43124_ (.A(_15994_),
    .Y(_16014_));
 sky130_fd_sc_hd__a31o_1 _43125_ (.A1(_16014_),
    .A2(_15995_),
    .A3(_16002_),
    .B1(_16005_),
    .X(_16015_));
 sky130_fd_sc_hd__a21oi_1 _43126_ (.A1(_16013_),
    .A2(_16015_),
    .B1(_12881_),
    .Y(_16016_));
 sky130_fd_sc_hd__a2111oi_1 _43127_ (.A1(_14857_),
    .A2(_14609_),
    .B1(net88),
    .C1(_14215_),
    .D1(_13802_),
    .Y(_16017_));
 sky130_fd_sc_hd__inv_2 _43128_ (.A(net84),
    .Y(_16018_));
 sky130_fd_sc_hd__o31a_1 _43129_ (.A1(_14857_),
    .A2(_14605_),
    .A3(_14607_),
    .B1(_16018_),
    .X(_16019_));
 sky130_fd_sc_hd__o21ai_1 _43130_ (.A1(_16012_),
    .A2(_16016_),
    .B1(_16019_),
    .Y(_16021_));
 sky130_fd_sc_hd__buf_2 _43131_ (.A(net88),
    .X(_16022_));
 sky130_fd_sc_hd__buf_2 _43132_ (.A(net86),
    .X(_16023_));
 sky130_fd_sc_hd__and3_1 _43133_ (.A(_16014_),
    .B(_15995_),
    .C(_16002_),
    .X(_16024_));
 sky130_fd_sc_hd__o211ai_4 _43134_ (.A1(_16005_),
    .A2(_16024_),
    .B1(_13294_),
    .C1(_16013_),
    .Y(_16025_));
 sky130_fd_sc_hd__o21bai_2 _43135_ (.A1(_16011_),
    .A2(_16006_),
    .B1_N(_13294_),
    .Y(_16026_));
 sky130_fd_sc_hd__o211ai_4 _43136_ (.A1(_16022_),
    .A2(_16023_),
    .B1(_16025_),
    .C1(_16026_),
    .Y(_16027_));
 sky130_fd_sc_hd__a31o_1 _43137_ (.A1(_16010_),
    .A2(_15408_),
    .A3(_15411_),
    .B1(_15423_),
    .X(_16028_));
 sky130_fd_sc_hd__a21oi_1 _43138_ (.A1(_16021_),
    .A2(_16027_),
    .B1(_16028_),
    .Y(_16029_));
 sky130_fd_sc_hd__o21a_1 _43139_ (.A1(_15161_),
    .A2(_15419_),
    .B1(_15421_),
    .X(_16030_));
 sky130_fd_sc_hd__a21o_1 _43140_ (.A1(_11580_),
    .A2(_14608_),
    .B1(_16023_),
    .X(_16032_));
 sky130_fd_sc_hd__a21oi_2 _43141_ (.A1(_16025_),
    .A2(_16026_),
    .B1(_16032_),
    .Y(_16033_));
 sky130_fd_sc_hd__o21ai_1 _43142_ (.A1(_15428_),
    .A2(_15423_),
    .B1(_16027_),
    .Y(_16034_));
 sky130_fd_sc_hd__o22ai_4 _43143_ (.A1(_15424_),
    .A2(_16030_),
    .B1(_16033_),
    .B2(_16034_),
    .Y(_16035_));
 sky130_fd_sc_hd__nor2_2 _43144_ (.A(_16029_),
    .B(_16035_),
    .Y(_16036_));
 sky130_fd_sc_hd__a31o_1 _43145_ (.A1(_15161_),
    .A2(_15426_),
    .A3(_15431_),
    .B1(_15421_),
    .X(_16037_));
 sky130_fd_sc_hd__o211a_1 _43146_ (.A1(_16022_),
    .A2(_16023_),
    .B1(_16025_),
    .C1(_16026_),
    .X(_16038_));
 sky130_fd_sc_hd__o21bai_1 _43147_ (.A1(_16033_),
    .A2(_16038_),
    .B1_N(_16028_),
    .Y(_16039_));
 sky130_fd_sc_hd__o211ai_1 _43148_ (.A1(_15428_),
    .A2(_15423_),
    .B1(_16021_),
    .C1(_16027_),
    .Y(_16040_));
 sky130_fd_sc_hd__a22oi_2 _43149_ (.A1(_15439_),
    .A2(_16037_),
    .B1(_16039_),
    .B2(_16040_),
    .Y(_16041_));
 sky130_fd_sc_hd__clkbuf_2 _43150_ (.A(_13296_),
    .X(_16043_));
 sky130_fd_sc_hd__clkbuf_2 _43151_ (.A(_03068_),
    .X(_16044_));
 sky130_fd_sc_hd__nand2_1 _43152_ (.A(_16044_),
    .B(_12151_),
    .Y(_16045_));
 sky130_fd_sc_hd__o21ai_2 _43153_ (.A1(_16044_),
    .A2(_05101_),
    .B1(_16045_),
    .Y(_16046_));
 sky130_fd_sc_hd__xor2_1 _43154_ (.A(_16043_),
    .B(_16046_),
    .X(_16047_));
 sky130_fd_sc_hd__o21bai_1 _43155_ (.A1(_16036_),
    .A2(_16041_),
    .B1_N(_16047_),
    .Y(_16048_));
 sky130_fd_sc_hd__or3_1 _43156_ (.A(_14863_),
    .B(_14864_),
    .C(_14862_),
    .X(_16049_));
 sky130_fd_sc_hd__a21oi_2 _43157_ (.A1(_16049_),
    .A2(_14869_),
    .B1(_14865_),
    .Y(_16050_));
 sky130_fd_sc_hd__clkbuf_2 _43158_ (.A(_16029_),
    .X(_16051_));
 sky130_fd_sc_hd__o211a_1 _43159_ (.A1(_15428_),
    .A2(_15423_),
    .B1(_16021_),
    .C1(_16027_),
    .X(_16052_));
 sky130_fd_sc_hd__o2bb2ai_2 _43160_ (.A1_N(_15439_),
    .A2_N(_16037_),
    .B1(_16051_),
    .B2(_16052_),
    .Y(_16054_));
 sky130_fd_sc_hd__o211ai_2 _43161_ (.A1(_16051_),
    .A2(_16035_),
    .B1(_16047_),
    .C1(_16054_),
    .Y(_16055_));
 sky130_fd_sc_hd__nand3_2 _43162_ (.A(_16048_),
    .B(_16050_),
    .C(_16055_),
    .Y(_16056_));
 sky130_fd_sc_hd__o31a_2 _43163_ (.A1(_14863_),
    .A2(_14864_),
    .A3(_14862_),
    .B1(_14869_),
    .X(_16057_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43164_ (.A(_12875_),
    .X(_16058_));
 sky130_fd_sc_hd__buf_2 _43165_ (.A(_16058_),
    .X(_16059_));
 sky130_fd_sc_hd__xor2_2 _43166_ (.A(_16059_),
    .B(_16046_),
    .X(_16060_));
 sky130_fd_sc_hd__o211ai_2 _43167_ (.A1(_16035_),
    .A2(_16051_),
    .B1(_16060_),
    .C1(_16054_),
    .Y(_16061_));
 sky130_fd_sc_hd__o21bai_2 _43168_ (.A1(_16036_),
    .A2(_16041_),
    .B1_N(_16060_),
    .Y(_16062_));
 sky130_fd_sc_hd__o211ai_4 _43169_ (.A1(_14865_),
    .A2(_16057_),
    .B1(_16061_),
    .C1(_16062_),
    .Y(_16063_));
 sky130_fd_sc_hd__o211a_1 _43170_ (.A1(_15824_),
    .A2(_15457_),
    .B1(_16056_),
    .C1(_16063_),
    .X(_16065_));
 sky130_fd_sc_hd__o2bb2a_1 _43171_ (.A1_N(_15455_),
    .A2_N(_15442_),
    .B1(_15452_),
    .B2(_15451_),
    .X(_16066_));
 sky130_fd_sc_hd__a21boi_4 _43172_ (.A1(_16056_),
    .A2(_16063_),
    .B1_N(_16066_),
    .Y(_16067_));
 sky130_fd_sc_hd__o22ai_4 _43173_ (.A1(_15821_),
    .A2(_15823_),
    .B1(_16065_),
    .B2(_16067_),
    .Y(_16068_));
 sky130_fd_sc_hd__clkbuf_2 _43174_ (.A(_16063_),
    .X(_16069_));
 sky130_fd_sc_hd__a21bo_1 _43175_ (.A1(_16056_),
    .A2(_16069_),
    .B1_N(_16066_),
    .X(_16070_));
 sky130_fd_sc_hd__nor2_1 _43176_ (.A(_15821_),
    .B(_15823_),
    .Y(_16071_));
 sky130_fd_sc_hd__o211ai_2 _43177_ (.A1(_15824_),
    .A2(_15457_),
    .B1(_16056_),
    .C1(_16069_),
    .Y(_16072_));
 sky130_fd_sc_hd__nand3_1 _43178_ (.A(_16070_),
    .B(_16071_),
    .C(_16072_),
    .Y(_16073_));
 sky130_fd_sc_hd__a22oi_2 _43179_ (.A1(_15155_),
    .A2(_15598_),
    .B1(_16068_),
    .B2(_16073_),
    .Y(_16074_));
 sky130_fd_sc_hd__nand2_1 _43180_ (.A(_16071_),
    .B(_16072_),
    .Y(_16076_));
 sky130_fd_sc_hd__inv_2 _43181_ (.A(_15156_),
    .Y(_16077_));
 sky130_fd_sc_hd__a31o_1 _43182_ (.A1(_15155_),
    .A2(_15462_),
    .A3(_15464_),
    .B1(_16077_),
    .X(_16078_));
 sky130_fd_sc_hd__o211a_1 _43183_ (.A1(_16067_),
    .A2(_16076_),
    .B1(_16078_),
    .C1(_16068_),
    .X(_16079_));
 sky130_fd_sc_hd__o22ai_1 _43184_ (.A1(_15596_),
    .A2(_15597_),
    .B1(_16074_),
    .B2(_16079_),
    .Y(_16080_));
 sky130_fd_sc_hd__nor2_1 _43185_ (.A(_15596_),
    .B(_15597_),
    .Y(_16081_));
 sky130_fd_sc_hd__a21o_1 _43186_ (.A1(_16068_),
    .A2(_16073_),
    .B1(_16078_),
    .X(_16082_));
 sky130_fd_sc_hd__o211ai_1 _43187_ (.A1(_16067_),
    .A2(_16076_),
    .B1(_16078_),
    .C1(_16068_),
    .Y(_16083_));
 sky130_fd_sc_hd__nand3_1 _43188_ (.A(_16081_),
    .B(_16082_),
    .C(_16083_),
    .Y(_16084_));
 sky130_fd_sc_hd__nand3_1 _43189_ (.A(_15564_),
    .B(_16080_),
    .C(_16084_),
    .Y(_16085_));
 sky130_fd_sc_hd__o21ai_1 _43190_ (.A1(_16074_),
    .A2(_16079_),
    .B1(_16081_),
    .Y(_16087_));
 sky130_fd_sc_hd__a32oi_2 _43191_ (.A1(_15470_),
    .A2(_15472_),
    .A3(_15473_),
    .B1(_15517_),
    .B2(_15521_),
    .Y(_16088_));
 sky130_fd_sc_hd__o22a_1 _43192_ (.A1(_15821_),
    .A2(_15823_),
    .B1(_16065_),
    .B2(_16067_),
    .X(_16089_));
 sky130_fd_sc_hd__o21ai_1 _43193_ (.A1(_16067_),
    .A2(_16076_),
    .B1(_16078_),
    .Y(_16090_));
 sky130_fd_sc_hd__o221ai_2 _43194_ (.A1(_15596_),
    .A2(_15597_),
    .B1(_16089_),
    .B2(_16090_),
    .C1(_16082_),
    .Y(_16091_));
 sky130_fd_sc_hd__nand3_2 _43195_ (.A(_16087_),
    .B(_16088_),
    .C(_16091_),
    .Y(_16092_));
 sky130_fd_sc_hd__o21ai_1 _43196_ (.A1(_15509_),
    .A2(_15476_),
    .B1(_15513_),
    .Y(_16093_));
 sky130_fd_sc_hd__a21oi_4 _43197_ (.A1(_14808_),
    .A2(_14791_),
    .B1(_14807_),
    .Y(_16094_));
 sky130_fd_sc_hd__and3_1 _43198_ (.A(_15495_),
    .B(_15496_),
    .C(_15502_),
    .X(_16095_));
 sky130_fd_sc_hd__and2_1 _43199_ (.A(_15488_),
    .B(_15503_),
    .X(_16096_));
 sky130_fd_sc_hd__o221a_1 _43200_ (.A1(_03002_),
    .A2(_14796_),
    .B1(_04551_),
    .B2(_08969_),
    .C1(_08967_),
    .X(_16098_));
 sky130_fd_sc_hd__a211oi_1 _43201_ (.A1(_03005_),
    .A2(_10297_),
    .B1(_08969_),
    .C1(_04551_),
    .Y(_16099_));
 sky130_fd_sc_hd__o21ai_2 _43202_ (.A1(_07508_),
    .A2(_08961_),
    .B1(_14796_),
    .Y(_16100_));
 sky130_fd_sc_hd__o31a_2 _43203_ (.A1(_14796_),
    .A2(_16098_),
    .A3(_16099_),
    .B1(_16100_),
    .X(_16101_));
 sky130_fd_sc_hd__a21oi_2 _43204_ (.A1(_15487_),
    .A2(_14706_),
    .B1(_16101_),
    .Y(_16102_));
 sky130_fd_sc_hd__nor2_1 _43205_ (.A(_01420_),
    .B(_04582_),
    .Y(_16103_));
 sky130_fd_sc_hd__a31o_2 _43206_ (.A1(_15487_),
    .A2(_16103_),
    .A3(_03005_),
    .B1(_14801_),
    .X(_16104_));
 sky130_fd_sc_hd__and3_1 _43207_ (.A(_15487_),
    .B(_14706_),
    .C(_16101_),
    .X(_16105_));
 sky130_fd_sc_hd__or3_1 _43208_ (.A(_16102_),
    .B(_16104_),
    .C(_16105_),
    .X(_16106_));
 sky130_fd_sc_hd__o21ai_1 _43209_ (.A1(_16105_),
    .A2(_16102_),
    .B1(_16104_),
    .Y(_16107_));
 sky130_fd_sc_hd__and4bb_1 _43210_ (.A_N(_16095_),
    .B_N(_16096_),
    .C(_16106_),
    .D(_16107_),
    .X(_16109_));
 sky130_fd_sc_hd__a2bb2oi_2 _43211_ (.A1_N(_16095_),
    .A2_N(_16096_),
    .B1(_16106_),
    .B2(_16107_),
    .Y(_16110_));
 sky130_fd_sc_hd__a21oi_4 _43212_ (.A1(_14804_),
    .A2(_14795_),
    .B1(_14802_),
    .Y(_16111_));
 sky130_fd_sc_hd__o21a_1 _43213_ (.A1(_16109_),
    .A2(_16110_),
    .B1(_16111_),
    .X(_16112_));
 sky130_fd_sc_hd__nor3_1 _43214_ (.A(_16111_),
    .B(_16109_),
    .C(_16110_),
    .Y(_16113_));
 sky130_fd_sc_hd__or2_2 _43215_ (.A(_16112_),
    .B(_16113_),
    .X(_16114_));
 sky130_fd_sc_hd__xnor2_1 _43216_ (.A(_16094_),
    .B(_16114_),
    .Y(_16115_));
 sky130_fd_sc_hd__a21o_1 _43217_ (.A1(_15511_),
    .A2(_16093_),
    .B1(_16115_),
    .X(_16116_));
 sky130_fd_sc_hd__nand3_1 _43218_ (.A(_15511_),
    .B(_16093_),
    .C(_16115_),
    .Y(_16117_));
 sky130_fd_sc_hd__and3_1 _43219_ (.A(_16116_),
    .B(_16117_),
    .C(_14812_),
    .X(_16118_));
 sky130_fd_sc_hd__a21oi_1 _43220_ (.A1(_16116_),
    .A2(_16117_),
    .B1(_14812_),
    .Y(_16120_));
 sky130_fd_sc_hd__nor2_1 _43221_ (.A(_16118_),
    .B(_16120_),
    .Y(_16121_));
 sky130_fd_sc_hd__a21oi_1 _43222_ (.A1(_16085_),
    .A2(_16092_),
    .B1(_16121_),
    .Y(_16122_));
 sky130_fd_sc_hd__and3_1 _43223_ (.A(_16085_),
    .B(_16092_),
    .C(_16121_),
    .X(_16123_));
 sky130_fd_sc_hd__a21bo_1 _43224_ (.A1(_15542_),
    .A2(_15523_),
    .B1_N(_15530_),
    .X(_16124_));
 sky130_fd_sc_hd__o21bai_1 _43225_ (.A1(_16122_),
    .A2(_16123_),
    .B1_N(_16124_),
    .Y(_16125_));
 sky130_fd_sc_hd__o2bb2ai_1 _43226_ (.A1_N(_16085_),
    .A2_N(_16092_),
    .B1(_16118_),
    .B2(_16120_),
    .Y(_16126_));
 sky130_fd_sc_hd__nand3_1 _43227_ (.A(_16085_),
    .B(_16092_),
    .C(_16121_),
    .Y(_16127_));
 sky130_fd_sc_hd__nand3_1 _43228_ (.A(_16124_),
    .B(_16126_),
    .C(_16127_),
    .Y(_16128_));
 sky130_fd_sc_hd__nand3b_2 _43229_ (.A_N(_15541_),
    .B(_16125_),
    .C(_16128_),
    .Y(_16129_));
 sky130_fd_sc_hd__nand2_1 _43230_ (.A(_15545_),
    .B(_15540_),
    .Y(_16131_));
 sky130_fd_sc_hd__nand2_1 _43231_ (.A(_16124_),
    .B(_16127_),
    .Y(_16132_));
 sky130_fd_sc_hd__o21ai_1 _43232_ (.A1(_16122_),
    .A2(_16132_),
    .B1(_16125_),
    .Y(_16133_));
 sky130_fd_sc_hd__a22oi_2 _43233_ (.A1(_15549_),
    .A2(_16131_),
    .B1(_16133_),
    .B2(_15541_),
    .Y(_16134_));
 sky130_fd_sc_hd__a21oi_1 _43234_ (.A1(_16126_),
    .A2(_16127_),
    .B1(_16124_),
    .Y(_16135_));
 sky130_fd_sc_hd__nor2_1 _43235_ (.A(_16122_),
    .B(_16132_),
    .Y(_16136_));
 sky130_fd_sc_hd__o22ai_2 _43236_ (.A1(_14819_),
    .A2(_14816_),
    .B1(_16135_),
    .B2(_16136_),
    .Y(_16137_));
 sky130_fd_sc_hd__a2bb2o_1 _43237_ (.A1_N(_15531_),
    .A2_N(_15538_),
    .B1(_15540_),
    .B2(_15544_),
    .X(_16138_));
 sky130_fd_sc_hd__a21oi_2 _43238_ (.A1(_16137_),
    .A2(_16129_),
    .B1(_16138_),
    .Y(_16139_));
 sky130_fd_sc_hd__a21oi_4 _43239_ (.A1(_16129_),
    .A2(_16134_),
    .B1(_16139_),
    .Y(_16140_));
 sky130_fd_sc_hd__xor2_1 _43240_ (.A(_15563_),
    .B(_16140_),
    .X(_00017_));
 sky130_fd_sc_hd__clkbuf_2 _43241_ (.A(_15593_),
    .X(_16142_));
 sky130_fd_sc_hd__nand3_1 _43242_ (.A(_15595_),
    .B(_16142_),
    .C(_15594_),
    .Y(_16143_));
 sky130_fd_sc_hd__a21oi_2 _43243_ (.A1(_04553_),
    .A2(_08962_),
    .B1(_15579_),
    .Y(_16144_));
 sky130_fd_sc_hd__and4b_2 _43244_ (.A_N(_07498_),
    .B(_12764_),
    .C(_10429_),
    .D(_15576_),
    .X(_16145_));
 sky130_fd_sc_hd__or4b_2 _43245_ (.A(_03002_),
    .B(_14796_),
    .C(_04553_),
    .D_N(_15576_),
    .X(_16146_));
 sky130_fd_sc_hd__o211ai_4 _43246_ (.A1(_16144_),
    .A2(_16145_),
    .B1(_16100_),
    .C1(_16146_),
    .Y(_16147_));
 sky130_fd_sc_hd__a21o_1 _43247_ (.A1(_16100_),
    .A2(_16146_),
    .B1(_16144_),
    .X(_16148_));
 sky130_fd_sc_hd__a211oi_2 _43248_ (.A1(_16147_),
    .A2(_16148_),
    .B1(_15586_),
    .C1(_15587_),
    .Y(_16149_));
 sky130_fd_sc_hd__o211a_1 _43249_ (.A1(_15586_),
    .A2(_15587_),
    .B1(_16147_),
    .C1(_16148_),
    .X(_16150_));
 sky130_fd_sc_hd__inv_2 _43250_ (.A(_16102_),
    .Y(_16152_));
 sky130_fd_sc_hd__a21oi_1 _43251_ (.A1(_16104_),
    .A2(_16152_),
    .B1(_16105_),
    .Y(_16153_));
 sky130_fd_sc_hd__o21bai_2 _43252_ (.A1(_16149_),
    .A2(_16150_),
    .B1_N(_16153_),
    .Y(_16154_));
 sky130_fd_sc_hd__a2111o_1 _43253_ (.A1(_16104_),
    .A2(_16152_),
    .B1(_16149_),
    .C1(_16150_),
    .D1(_16105_),
    .X(_16155_));
 sky130_fd_sc_hd__nand2_1 _43254_ (.A(_16154_),
    .B(_16155_),
    .Y(_16156_));
 sky130_fd_sc_hd__or3_1 _43255_ (.A(_16110_),
    .B(_16156_),
    .C(_16113_),
    .X(_16157_));
 sky130_fd_sc_hd__a2bb2o_2 _43256_ (.A1_N(_16110_),
    .A2_N(_16113_),
    .B1(_16154_),
    .B2(_16155_),
    .X(_16158_));
 sky130_fd_sc_hd__nand2_1 _43257_ (.A(_16157_),
    .B(_16158_),
    .Y(_16159_));
 sky130_fd_sc_hd__a21o_2 _43258_ (.A1(_16142_),
    .A2(_16143_),
    .B1(_16159_),
    .X(_16160_));
 sky130_fd_sc_hd__a311oi_1 _43259_ (.A1(_16142_),
    .A2(_16143_),
    .A3(_16159_),
    .B1(_16114_),
    .C1(_16094_),
    .Y(_16161_));
 sky130_fd_sc_hd__nand3_1 _43260_ (.A(_16142_),
    .B(_16143_),
    .C(_16159_),
    .Y(_16163_));
 sky130_fd_sc_hd__a2bb2oi_1 _43261_ (.A1_N(_16114_),
    .A2_N(_16094_),
    .B1(_16163_),
    .B2(_16160_),
    .Y(_16164_));
 sky130_fd_sc_hd__a21o_1 _43262_ (.A1(_16160_),
    .A2(_16161_),
    .B1(_16164_),
    .X(_16165_));
 sky130_fd_sc_hd__o31a_1 _43263_ (.A1(_15596_),
    .A2(_15597_),
    .A3(_16074_),
    .B1(_16083_),
    .X(_16166_));
 sky130_fd_sc_hd__nor2_2 _43264_ (.A(_15603_),
    .B(_15627_),
    .Y(_16167_));
 sky130_fd_sc_hd__a21oi_2 _43265_ (.A1(_14854_),
    .A2(_15600_),
    .B1(_15628_),
    .Y(_16168_));
 sky130_fd_sc_hd__inv_2 _43266_ (.A(_16028_),
    .Y(_16169_));
 sky130_fd_sc_hd__o21ai_1 _43267_ (.A1(_16169_),
    .A2(_16033_),
    .B1(_16027_),
    .Y(_16170_));
 sky130_fd_sc_hd__clkbuf_2 _43268_ (.A(_16010_),
    .X(_16171_));
 sky130_fd_sc_hd__a21oi_1 _43269_ (.A1(_15408_),
    .A2(_16003_),
    .B1(_16024_),
    .Y(_16172_));
 sky130_fd_sc_hd__a31o_1 _43270_ (.A1(_16010_),
    .A2(_16004_),
    .A3(_16008_),
    .B1(_12881_),
    .X(_16174_));
 sky130_fd_sc_hd__and2_2 _43271_ (.A(_15401_),
    .B(_15402_),
    .X(_16175_));
 sky130_fd_sc_hd__o21ai_2 _43272_ (.A1(_14186_),
    .A2(_14191_),
    .B1(_16175_),
    .Y(_16176_));
 sky130_fd_sc_hd__o2111ai_4 _43273_ (.A1(_15403_),
    .A2(_16175_),
    .B1(_16176_),
    .C1(_16014_),
    .D1(_15995_),
    .Y(_16177_));
 sky130_fd_sc_hd__a21boi_2 _43274_ (.A1(_15900_),
    .A2(_15953_),
    .B1_N(_15904_),
    .Y(_16178_));
 sky130_fd_sc_hd__a31oi_2 _43275_ (.A1(_15209_),
    .A2(_15836_),
    .A3(_15838_),
    .B1(_15853_),
    .Y(_16179_));
 sky130_fd_sc_hd__a31o_1 _43276_ (.A1(_13970_),
    .A2(_13972_),
    .A3(_15186_),
    .B1(_13980_),
    .X(_16180_));
 sky130_fd_sc_hd__a31o_1 _43277_ (.A1(_13968_),
    .A2(_13951_),
    .A3(_13945_),
    .B1(_13980_),
    .X(_16181_));
 sky130_fd_sc_hd__a21oi_1 _43278_ (.A1(_15828_),
    .A2(_15831_),
    .B1(_15834_),
    .Y(_16182_));
 sky130_fd_sc_hd__o22ai_4 _43279_ (.A1(_16181_),
    .A2(_15832_),
    .B1(_13982_),
    .B2(_16182_),
    .Y(_16183_));
 sky130_fd_sc_hd__a21o_1 _43280_ (.A1(_15193_),
    .A2(_16180_),
    .B1(_16183_),
    .X(_16185_));
 sky130_fd_sc_hd__nand2_1 _43281_ (.A(_16183_),
    .B(_15835_),
    .Y(_16186_));
 sky130_fd_sc_hd__and2_1 _43282_ (.A(_15878_),
    .B(_15216_),
    .X(_16187_));
 sky130_fd_sc_hd__and4b_1 _43283_ (.A_N(_14010_),
    .B(_15881_),
    .C(_15217_),
    .D(_10500_),
    .X(_16188_));
 sky130_fd_sc_hd__o21ba_1 _43284_ (.A1(_16187_),
    .A2(_15847_),
    .B1_N(_16188_),
    .X(_16189_));
 sky130_fd_sc_hd__a21o_1 _43285_ (.A1(_16185_),
    .A2(_16186_),
    .B1(_16189_),
    .X(_16190_));
 sky130_fd_sc_hd__nand3_1 _43286_ (.A(_16185_),
    .B(_16186_),
    .C(_16189_),
    .Y(_16191_));
 sky130_fd_sc_hd__nand2_1 _43287_ (.A(_16190_),
    .B(_16191_),
    .Y(_16192_));
 sky130_fd_sc_hd__o21bai_2 _43288_ (.A1(_15839_),
    .A2(_16179_),
    .B1_N(_16192_),
    .Y(_16193_));
 sky130_fd_sc_hd__o211ai_4 _43289_ (.A1(_15853_),
    .A2(_15837_),
    .B1(_15856_),
    .C1(_16192_),
    .Y(_16194_));
 sky130_fd_sc_hd__o21ai_2 _43290_ (.A1(_15224_),
    .A2(_15841_),
    .B1(_14019_),
    .Y(_16196_));
 sky130_fd_sc_hd__or3_2 _43291_ (.A(_13006_),
    .B(_16187_),
    .C(_15845_),
    .X(_16197_));
 sky130_fd_sc_hd__o21ai_4 _43292_ (.A1(_15217_),
    .A2(_15842_),
    .B1(_16197_),
    .Y(_16198_));
 sky130_fd_sc_hd__and3_1 _43293_ (.A(_15878_),
    .B(_07691_),
    .C(_14060_),
    .X(_16199_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43294_ (.A(_15868_),
    .X(_16200_));
 sky130_fd_sc_hd__nor2_1 _43295_ (.A(_16200_),
    .B(_15881_),
    .Y(_16201_));
 sky130_fd_sc_hd__a21oi_1 _43296_ (.A1(_16200_),
    .A2(_16199_),
    .B1(_16201_),
    .Y(_16202_));
 sky130_fd_sc_hd__nand2_1 _43297_ (.A(_15867_),
    .B(_07665_),
    .Y(_16203_));
 sky130_fd_sc_hd__mux2_1 _43298_ (.A0(_16199_),
    .A1(_16202_),
    .S(_16203_),
    .X(_16204_));
 sky130_fd_sc_hd__or3_1 _43299_ (.A(_16196_),
    .B(_16198_),
    .C(_16204_),
    .X(_16205_));
 sky130_fd_sc_hd__o21ai_1 _43300_ (.A1(_16196_),
    .A2(_16198_),
    .B1(_16204_),
    .Y(_16207_));
 sky130_fd_sc_hd__and2_1 _43301_ (.A(_16205_),
    .B(_16207_),
    .X(_16208_));
 sky130_fd_sc_hd__xnor2_1 _43302_ (.A(_15851_),
    .B(_16208_),
    .Y(_16209_));
 sky130_fd_sc_hd__and3_1 _43303_ (.A(_15886_),
    .B(_15887_),
    .C(_16209_),
    .X(_16210_));
 sky130_fd_sc_hd__a21oi_1 _43304_ (.A1(_15886_),
    .A2(_15887_),
    .B1(_16209_),
    .Y(_16211_));
 sky130_fd_sc_hd__nor2_2 _43305_ (.A(_16210_),
    .B(_16211_),
    .Y(_16212_));
 sky130_fd_sc_hd__a21oi_2 _43306_ (.A1(_16193_),
    .A2(_16194_),
    .B1(_16212_),
    .Y(_16213_));
 sky130_fd_sc_hd__and3_1 _43307_ (.A(_16193_),
    .B(_16194_),
    .C(_16212_),
    .X(_16214_));
 sky130_fd_sc_hd__nor2_1 _43308_ (.A(_16213_),
    .B(_16214_),
    .Y(_16215_));
 sky130_fd_sc_hd__a21oi_2 _43309_ (.A1(_15854_),
    .A2(_15857_),
    .B1(_15863_),
    .Y(_16216_));
 sky130_fd_sc_hd__o21ai_1 _43310_ (.A1(_15896_),
    .A2(_16216_),
    .B1(_15865_),
    .Y(_16218_));
 sky130_fd_sc_hd__nand2_2 _43311_ (.A(_16215_),
    .B(_16218_),
    .Y(_16219_));
 sky130_fd_sc_hd__o221ai_4 _43312_ (.A1(_16216_),
    .A2(_15896_),
    .B1(_16213_),
    .B2(_16214_),
    .C1(_15865_),
    .Y(_16220_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43313_ (.A(_15925_),
    .X(_16221_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43314_ (.A(_13105_),
    .X(_16222_));
 sky130_fd_sc_hd__o21ai_1 _43315_ (.A1(_15294_),
    .A2(_16221_),
    .B1(_16222_),
    .Y(_16223_));
 sky130_fd_sc_hd__and2_1 _43316_ (.A(_15926_),
    .B(_15329_),
    .X(_16224_));
 sky130_fd_sc_hd__or2_1 _43317_ (.A(_10803_),
    .B(_10804_),
    .X(_16225_));
 sky130_fd_sc_hd__o221a_1 _43318_ (.A1(_15927_),
    .A2(_15928_),
    .B1(_16224_),
    .B2(_16225_),
    .C1(_13140_),
    .X(_16226_));
 sky130_fd_sc_hd__or3_1 _43319_ (.A(_10803_),
    .B(_10804_),
    .C(_16224_),
    .X(_16227_));
 sky130_fd_sc_hd__a21oi_1 _43320_ (.A1(_16227_),
    .A2(_13140_),
    .B1(_15929_),
    .Y(_16229_));
 sky130_fd_sc_hd__or4_2 _43321_ (.A(_15934_),
    .B(net159),
    .C(_16226_),
    .D(_16229_),
    .X(_16230_));
 sky130_fd_sc_hd__o22ai_4 _43322_ (.A1(_15934_),
    .A2(net159),
    .B1(_16226_),
    .B2(_16229_),
    .Y(_16231_));
 sky130_fd_sc_hd__and3_1 _43323_ (.A(_16223_),
    .B(_16230_),
    .C(_16231_),
    .X(_16232_));
 sky130_fd_sc_hd__a21oi_1 _43324_ (.A1(_16230_),
    .A2(_16231_),
    .B1(_16223_),
    .Y(_16233_));
 sky130_fd_sc_hd__o21ai_1 _43325_ (.A1(_15925_),
    .A2(_15926_),
    .B1(_16203_),
    .Y(_16234_));
 sky130_fd_sc_hd__or3_1 _43326_ (.A(_15925_),
    .B(_07668_),
    .C(_15926_),
    .X(_16235_));
 sky130_fd_sc_hd__and4bb_1 _43327_ (.A_N(_15874_),
    .B_N(_15875_),
    .C(_16234_),
    .D(_16235_),
    .X(_16236_));
 sky130_fd_sc_hd__a2bb2oi_1 _43328_ (.A1_N(_15874_),
    .A2_N(_15875_),
    .B1(_16234_),
    .B2(_16235_),
    .Y(_16237_));
 sky130_fd_sc_hd__a211o_1 _43329_ (.A1(_15912_),
    .A2(_15914_),
    .B1(_16236_),
    .C1(_16237_),
    .X(_16238_));
 sky130_fd_sc_hd__o211ai_1 _43330_ (.A1(_16236_),
    .A2(_16237_),
    .B1(_15912_),
    .C1(_15914_),
    .Y(_16240_));
 sky130_fd_sc_hd__o211a_1 _43331_ (.A1(_15916_),
    .A2(_15919_),
    .B1(_16238_),
    .C1(_16240_),
    .X(_16241_));
 sky130_fd_sc_hd__a211oi_1 _43332_ (.A1(_16238_),
    .A2(_16240_),
    .B1(_15916_),
    .C1(_15919_),
    .Y(_16242_));
 sky130_fd_sc_hd__or4_1 _43333_ (.A(_16232_),
    .B(_16233_),
    .C(_16241_),
    .D(_16242_),
    .X(_16243_));
 sky130_fd_sc_hd__o22ai_1 _43334_ (.A1(_16232_),
    .A2(_16233_),
    .B1(_16241_),
    .B2(_16242_),
    .Y(_16244_));
 sky130_fd_sc_hd__a21boi_1 _43335_ (.A1(_15893_),
    .A2(_15892_),
    .B1_N(_15891_),
    .Y(_16245_));
 sky130_fd_sc_hd__a21boi_1 _43336_ (.A1(_16243_),
    .A2(_16244_),
    .B1_N(_16245_),
    .Y(_16246_));
 sky130_fd_sc_hd__and3b_1 _43337_ (.A_N(_16245_),
    .B(_16243_),
    .C(_16244_),
    .X(_16247_));
 sky130_fd_sc_hd__o211a_1 _43338_ (.A1(_16246_),
    .A2(_16247_),
    .B1(_15923_),
    .C1(_15946_),
    .X(_16248_));
 sky130_fd_sc_hd__a211oi_2 _43339_ (.A1(_15923_),
    .A2(_15946_),
    .B1(_16246_),
    .C1(_16247_),
    .Y(_16249_));
 sky130_fd_sc_hd__nor2_1 _43340_ (.A(_16248_),
    .B(_16249_),
    .Y(_16251_));
 sky130_fd_sc_hd__a21o_1 _43341_ (.A1(_16219_),
    .A2(_16220_),
    .B1(_16251_),
    .X(_16252_));
 sky130_fd_sc_hd__nand3_2 _43342_ (.A(_16219_),
    .B(_16220_),
    .C(_16251_),
    .Y(_16253_));
 sky130_fd_sc_hd__nand2_1 _43343_ (.A(_16252_),
    .B(_16253_),
    .Y(_16254_));
 sky130_fd_sc_hd__nor2_1 _43344_ (.A(_16178_),
    .B(_16254_),
    .Y(_16255_));
 sky130_fd_sc_hd__or2b_1 _43345_ (.A(_15971_),
    .B_N(_15961_),
    .X(_16256_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43346_ (.A(_13205_),
    .X(_16257_));
 sky130_fd_sc_hd__or3_1 _43347_ (.A(_16257_),
    .B(_15369_),
    .C(_15924_),
    .X(_16258_));
 sky130_fd_sc_hd__o21ai_1 _43348_ (.A1(_16257_),
    .A2(_15370_),
    .B1(_15924_),
    .Y(_16259_));
 sky130_fd_sc_hd__nand2_1 _43349_ (.A(_16258_),
    .B(_16259_),
    .Y(_16260_));
 sky130_fd_sc_hd__a21o_1 _43350_ (.A1(_15938_),
    .A2(_15941_),
    .B1(_16260_),
    .X(_16262_));
 sky130_fd_sc_hd__o211ai_1 _43351_ (.A1(_15924_),
    .A2(_15940_),
    .B1(_16260_),
    .C1(_15938_),
    .Y(_16263_));
 sky130_fd_sc_hd__o2111ai_1 _43352_ (.A1(_16257_),
    .A2(_15370_),
    .B1(_15963_),
    .C1(_16262_),
    .D1(_16263_),
    .Y(_16264_));
 sky130_fd_sc_hd__a21o_1 _43353_ (.A1(_16262_),
    .A2(_16263_),
    .B1(_15964_),
    .X(_16265_));
 sky130_fd_sc_hd__nand2_1 _43354_ (.A(_16264_),
    .B(_16265_),
    .Y(_16266_));
 sky130_fd_sc_hd__inv_2 _43355_ (.A(_15967_),
    .Y(_16267_));
 sky130_fd_sc_hd__o211ai_1 _43356_ (.A1(_15373_),
    .A2(_15968_),
    .B1(_16266_),
    .C1(_16267_),
    .Y(_16268_));
 sky130_fd_sc_hd__a21o_1 _43357_ (.A1(_16267_),
    .A2(_15969_),
    .B1(_16266_),
    .X(_16269_));
 sky130_fd_sc_hd__o21ai_2 _43358_ (.A1(_15905_),
    .A2(_15952_),
    .B1(_15951_),
    .Y(_16270_));
 sky130_fd_sc_hd__a21oi_1 _43359_ (.A1(_16268_),
    .A2(_16269_),
    .B1(_16270_),
    .Y(_16271_));
 sky130_fd_sc_hd__and3_1 _43360_ (.A(_16268_),
    .B(_16269_),
    .C(_16270_),
    .X(_16273_));
 sky130_fd_sc_hd__or2_1 _43361_ (.A(_16271_),
    .B(_16273_),
    .X(_16274_));
 sky130_fd_sc_hd__xnor2_1 _43362_ (.A(_16256_),
    .B(_16274_),
    .Y(_16275_));
 sky130_fd_sc_hd__a21o_1 _43363_ (.A1(_16254_),
    .A2(_16178_),
    .B1(_16275_),
    .X(_16276_));
 sky130_fd_sc_hd__nand2_1 _43364_ (.A(_15901_),
    .B(_15903_),
    .Y(_16277_));
 sky130_fd_sc_hd__o211a_1 _43365_ (.A1(_15894_),
    .A2(_15895_),
    .B1(_15860_),
    .C1(_15865_),
    .X(_16278_));
 sky130_fd_sc_hd__o2bb2ai_1 _43366_ (.A1_N(_15953_),
    .A2_N(_15900_),
    .B1(_16277_),
    .B2(_16278_),
    .Y(_16279_));
 sky130_fd_sc_hd__a21oi_1 _43367_ (.A1(_16252_),
    .A2(_16253_),
    .B1(_16279_),
    .Y(_16280_));
 sky130_fd_sc_hd__o21ai_1 _43368_ (.A1(_16280_),
    .A2(_16255_),
    .B1(_16275_),
    .Y(_16281_));
 sky130_fd_sc_hd__o21ai_4 _43369_ (.A1(_16255_),
    .A2(_16276_),
    .B1(_16281_),
    .Y(_16282_));
 sky130_fd_sc_hd__a21oi_1 _43370_ (.A1(_15982_),
    .A2(_15978_),
    .B1(_16282_),
    .Y(_16284_));
 sky130_fd_sc_hd__a21oi_1 _43371_ (.A1(_15957_),
    .A2(_15977_),
    .B1(_15979_),
    .Y(_16285_));
 sky130_fd_sc_hd__a21o_1 _43372_ (.A1(_15960_),
    .A2(_15972_),
    .B1(_15974_),
    .X(_16286_));
 sky130_fd_sc_hd__a21bo_1 _43373_ (.A1(_16282_),
    .A2(_16285_),
    .B1_N(_16286_),
    .X(_16287_));
 sky130_fd_sc_hd__xor2_1 _43374_ (.A(_16285_),
    .B(_16282_),
    .X(_16288_));
 sky130_fd_sc_hd__o22ai_4 _43375_ (.A1(_16284_),
    .A2(_16287_),
    .B1(_16286_),
    .B2(_16288_),
    .Y(_16289_));
 sky130_fd_sc_hd__a21boi_4 _43376_ (.A1(_15989_),
    .A2(_15988_),
    .B1_N(_15984_),
    .Y(_16290_));
 sky130_fd_sc_hd__nand2_1 _43377_ (.A(_16289_),
    .B(_16290_),
    .Y(_16291_));
 sky130_fd_sc_hd__or2_1 _43378_ (.A(_16290_),
    .B(_16289_),
    .X(_16292_));
 sky130_fd_sc_hd__nand2_4 _43379_ (.A(_16291_),
    .B(_16292_),
    .Y(_16293_));
 sky130_fd_sc_hd__a21oi_2 _43380_ (.A1(_16175_),
    .A2(_15403_),
    .B1(_15994_),
    .Y(_16295_));
 sky130_fd_sc_hd__a31o_1 _43381_ (.A1(_15993_),
    .A2(_15990_),
    .A3(_15991_),
    .B1(_16295_),
    .X(_16296_));
 sky130_fd_sc_hd__o211ai_4 _43382_ (.A1(_16177_),
    .A2(_16001_),
    .B1(_16293_),
    .C1(_16296_),
    .Y(_16297_));
 sky130_fd_sc_hd__o22ai_4 _43383_ (.A1(_15996_),
    .A2(_16295_),
    .B1(_16177_),
    .B2(_16001_),
    .Y(_16298_));
 sky130_fd_sc_hd__inv_2 _43384_ (.A(_16293_),
    .Y(_16299_));
 sky130_fd_sc_hd__nand2_2 _43385_ (.A(_16298_),
    .B(_16299_),
    .Y(_16300_));
 sky130_fd_sc_hd__buf_6 _43386_ (.A(_16300_),
    .X(_16301_));
 sky130_fd_sc_hd__o211a_2 _43387_ (.A1(_15162_),
    .A2(_15164_),
    .B1(_16297_),
    .C1(_16301_),
    .X(_16302_));
 sky130_fd_sc_hd__a21oi_2 _43388_ (.A1(_16297_),
    .A2(_16301_),
    .B1(_15429_),
    .Y(_16303_));
 sky130_fd_sc_hd__o21ai_1 _43389_ (.A1(_16302_),
    .A2(_16303_),
    .B1(_12881_),
    .Y(_16304_));
 sky130_fd_sc_hd__o211ai_2 _43390_ (.A1(_15162_),
    .A2(_15164_),
    .B1(_16297_),
    .C1(_16301_),
    .Y(_16306_));
 sky130_fd_sc_hd__a21o_1 _43391_ (.A1(_16297_),
    .A2(_16301_),
    .B1(_15429_),
    .X(_16307_));
 sky130_fd_sc_hd__nand3_1 _43392_ (.A(_16007_),
    .B(_16306_),
    .C(_16307_),
    .Y(_16308_));
 sky130_fd_sc_hd__nand3_2 _43393_ (.A(_16304_),
    .B(_16308_),
    .C(_16019_),
    .Y(_16309_));
 sky130_fd_sc_hd__nand2_1 _43394_ (.A(_16307_),
    .B(_13294_),
    .Y(_16310_));
 sky130_fd_sc_hd__o21ai_1 _43395_ (.A1(_16302_),
    .A2(_16303_),
    .B1(_16007_),
    .Y(_16311_));
 sky130_fd_sc_hd__o221ai_4 _43396_ (.A1(_16022_),
    .A2(_16023_),
    .B1(_16302_),
    .B2(_16310_),
    .C1(_16311_),
    .Y(_16312_));
 sky130_fd_sc_hd__o2111ai_2 _43397_ (.A1(_16171_),
    .A2(_16172_),
    .B1(_16174_),
    .C1(_16309_),
    .D1(_16312_),
    .Y(_16313_));
 sky130_fd_sc_hd__a22o_1 _43398_ (.A1(_16013_),
    .A2(_16174_),
    .B1(_16309_),
    .B2(_16312_),
    .X(_16314_));
 sky130_fd_sc_hd__nand3_1 _43399_ (.A(_16170_),
    .B(_16313_),
    .C(_16314_),
    .Y(_16315_));
 sky130_fd_sc_hd__inv_2 _43400_ (.A(_16315_),
    .Y(_16317_));
 sky130_fd_sc_hd__o2111a_1 _43401_ (.A1(_16171_),
    .A2(_16172_),
    .B1(_16174_),
    .C1(_16309_),
    .D1(_16312_),
    .X(_16318_));
 sky130_fd_sc_hd__a22oi_1 _43402_ (.A1(_16013_),
    .A2(_16174_),
    .B1(_16309_),
    .B2(_16312_),
    .Y(_16319_));
 sky130_fd_sc_hd__o21bai_2 _43403_ (.A1(_16318_),
    .A2(_16319_),
    .B1_N(_16170_),
    .Y(_16320_));
 sky130_fd_sc_hd__buf_1 _43404_ (.A(_12153_),
    .X(_16321_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43405_ (.A(_16321_),
    .X(_16322_));
 sky130_fd_sc_hd__buf_1 _43406_ (.A(_12151_),
    .X(_16323_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43407_ (.A(_16323_),
    .X(_16324_));
 sky130_fd_sc_hd__nor2_1 _43408_ (.A(_16322_),
    .B(_16324_),
    .Y(_16325_));
 sky130_fd_sc_hd__nand2_1 _43409_ (.A(_16320_),
    .B(_16325_),
    .Y(_16326_));
 sky130_fd_sc_hd__o2bb2ai_1 _43410_ (.A1_N(_16315_),
    .A2_N(_16320_),
    .B1(_16322_),
    .B2(_16324_),
    .Y(_16328_));
 sky130_fd_sc_hd__o221ai_2 _43411_ (.A1(_16167_),
    .A2(_16168_),
    .B1(_16317_),
    .B2(_16326_),
    .C1(_16328_),
    .Y(_16329_));
 sky130_fd_sc_hd__o21ai_1 _43412_ (.A1(_16322_),
    .A2(_16324_),
    .B1(_16320_),
    .Y(_16330_));
 sky130_fd_sc_hd__nor2_1 _43413_ (.A(_16167_),
    .B(_16168_),
    .Y(_16331_));
 sky130_fd_sc_hd__or2_1 _43414_ (.A(_16321_),
    .B(_16323_),
    .X(_16332_));
 sky130_fd_sc_hd__a21o_1 _43415_ (.A1(_16315_),
    .A2(_16320_),
    .B1(_16332_),
    .X(_16333_));
 sky130_fd_sc_hd__o211ai_4 _43416_ (.A1(_16317_),
    .A2(_16330_),
    .B1(_16331_),
    .C1(_16333_),
    .Y(_16334_));
 sky130_fd_sc_hd__a2bb2o_1 _43417_ (.A1_N(_16035_),
    .A2_N(_16051_),
    .B1(_16060_),
    .B2(_16054_),
    .X(_16335_));
 sky130_fd_sc_hd__a21o_1 _43418_ (.A1(_16329_),
    .A2(_16334_),
    .B1(_16335_),
    .X(_16336_));
 sky130_fd_sc_hd__and3_1 _43419_ (.A(_14854_),
    .B(_15600_),
    .C(_15628_),
    .X(_16337_));
 sky130_fd_sc_hd__o31ai_1 _43420_ (.A1(_15816_),
    .A2(_16168_),
    .A3(_16337_),
    .B1(_15817_),
    .Y(_16339_));
 sky130_fd_sc_hd__o21a_1 _43421_ (.A1(_15753_),
    .A2(_15727_),
    .B1(_15754_),
    .X(_16340_));
 sky130_fd_sc_hd__a21boi_1 _43422_ (.A1(_15713_),
    .A2(_15696_),
    .B1_N(_15697_),
    .Y(_16341_));
 sky130_fd_sc_hd__o31a_1 _43423_ (.A1(_15071_),
    .A2(_11209_),
    .A3(_15073_),
    .B1(_11206_),
    .X(_16342_));
 sky130_fd_sc_hd__buf_1 _43424_ (.A(_14296_),
    .X(_16343_));
 sky130_fd_sc_hd__buf_1 _43425_ (.A(_14294_),
    .X(_16344_));
 sky130_fd_sc_hd__a2bb2o_1 _43426_ (.A1_N(_16343_),
    .A2_N(_16344_),
    .B1(_12421_),
    .B2(_15087_),
    .X(_16345_));
 sky130_fd_sc_hd__a21oi_1 _43427_ (.A1(_16343_),
    .A2(_16344_),
    .B1(_16345_),
    .Y(_16346_));
 sky130_fd_sc_hd__a21oi_1 _43428_ (.A1(_15087_),
    .A2(_16343_),
    .B1(_16346_),
    .Y(_16347_));
 sky130_fd_sc_hd__a21o_1 _43429_ (.A1(_15730_),
    .A2(_15733_),
    .B1(_16347_),
    .X(_16348_));
 sky130_fd_sc_hd__nand3_1 _43430_ (.A(_15730_),
    .B(_15733_),
    .C(_16347_),
    .Y(_16350_));
 sky130_fd_sc_hd__a31o_1 _43431_ (.A1(_15113_),
    .A2(_15114_),
    .A3(_07119_),
    .B1(_15737_),
    .X(_16351_));
 sky130_fd_sc_hd__a31o_1 _43432_ (.A1(_15736_),
    .A2(_15109_),
    .A3(_15110_),
    .B1(_16351_),
    .X(_16352_));
 sky130_fd_sc_hd__a21bo_1 _43433_ (.A1(_15742_),
    .A2(_15744_),
    .B1_N(_15743_),
    .X(_16353_));
 sky130_fd_sc_hd__xnor2_1 _43434_ (.A(_16352_),
    .B(_16353_),
    .Y(_16354_));
 sky130_fd_sc_hd__o21bai_1 _43435_ (.A1(_15749_),
    .A2(_15751_),
    .B1_N(_15748_),
    .Y(_16355_));
 sky130_fd_sc_hd__and2b_1 _43436_ (.A_N(_16354_),
    .B(_16355_),
    .X(_16356_));
 sky130_fd_sc_hd__and2b_1 _43437_ (.A_N(_16355_),
    .B(_16354_),
    .X(_16357_));
 sky130_fd_sc_hd__nor2_1 _43438_ (.A(_16356_),
    .B(_16357_),
    .Y(_16358_));
 sky130_fd_sc_hd__nand3_1 _43439_ (.A(_16348_),
    .B(_16350_),
    .C(_16358_),
    .Y(_16359_));
 sky130_fd_sc_hd__a21o_1 _43440_ (.A1(_16348_),
    .A2(_16350_),
    .B1(_16358_),
    .X(_16361_));
 sky130_fd_sc_hd__o211a_1 _43441_ (.A1(_15725_),
    .A2(_16342_),
    .B1(_16359_),
    .C1(_16361_),
    .X(_16362_));
 sky130_fd_sc_hd__a211oi_1 _43442_ (.A1(_16359_),
    .A2(_16361_),
    .B1(_15725_),
    .C1(_16342_),
    .Y(_16363_));
 sky130_fd_sc_hd__or3_1 _43443_ (.A(net74),
    .B(_16362_),
    .C(_16363_),
    .X(_16364_));
 sky130_fd_sc_hd__o21ai_1 _43444_ (.A1(_16362_),
    .A2(_16363_),
    .B1(net74),
    .Y(_16365_));
 sky130_fd_sc_hd__nand2_1 _43445_ (.A(_16364_),
    .B(_16365_),
    .Y(_16366_));
 sky130_fd_sc_hd__xnor2_1 _43446_ (.A(_16340_),
    .B(_16366_),
    .Y(_16367_));
 sky130_fd_sc_hd__a31o_1 _43447_ (.A1(_14967_),
    .A2(_14986_),
    .A3(_15658_),
    .B1(_15716_),
    .X(_16368_));
 sky130_fd_sc_hd__inv_2 _43448_ (.A(net79),
    .Y(_16369_));
 sky130_fd_sc_hd__buf_1 _43449_ (.A(_14391_),
    .X(_16370_));
 sky130_fd_sc_hd__a2bb2o_1 _43450_ (.A1_N(_15648_),
    .A2_N(_16370_),
    .B1(_13573_),
    .B2(_14970_),
    .X(_16372_));
 sky130_fd_sc_hd__a21oi_1 _43451_ (.A1(_15648_),
    .A2(_16370_),
    .B1(_16372_),
    .Y(_16373_));
 sky130_fd_sc_hd__a21oi_2 _43452_ (.A1(_14970_),
    .A2(_15648_),
    .B1(_16373_),
    .Y(_16374_));
 sky130_fd_sc_hd__a21o_1 _43453_ (.A1(_15650_),
    .A2(_15651_),
    .B1(_16374_),
    .X(_16375_));
 sky130_fd_sc_hd__nand3_1 _43454_ (.A(_15650_),
    .B(_15651_),
    .C(_16374_),
    .Y(_16376_));
 sky130_fd_sc_hd__nand2_2 _43455_ (.A(_16375_),
    .B(_16376_),
    .Y(_16377_));
 sky130_fd_sc_hd__o21a_1 _43456_ (.A1(_14958_),
    .A2(_14369_),
    .B1(_13552_),
    .X(_16378_));
 sky130_fd_sc_hd__or2_1 _43457_ (.A(_15630_),
    .B(_16378_),
    .X(_16379_));
 sky130_fd_sc_hd__o31a_1 _43458_ (.A1(_13521_),
    .A2(_14945_),
    .A3(_14947_),
    .B1(_14353_),
    .X(_16380_));
 sky130_fd_sc_hd__nor4_1 _43459_ (.A(_16379_),
    .B(_16380_),
    .C(_15637_),
    .D(_15642_),
    .Y(_16381_));
 sky130_fd_sc_hd__o32a_1 _43460_ (.A1(_15630_),
    .A2(_15637_),
    .A3(_16378_),
    .B1(_16380_),
    .B2(_15642_),
    .X(_16383_));
 sky130_fd_sc_hd__nor2_1 _43461_ (.A(_16381_),
    .B(_16383_),
    .Y(_16384_));
 sky130_fd_sc_hd__xor2_4 _43462_ (.A(_16377_),
    .B(_16384_),
    .X(_16385_));
 sky130_fd_sc_hd__o211ai_4 _43463_ (.A1(_15653_),
    .A2(_15654_),
    .B1(_16369_),
    .C1(_16385_),
    .Y(_16386_));
 sky130_fd_sc_hd__a21oi_4 _43464_ (.A1(_16369_),
    .A2(_15655_),
    .B1(_16385_),
    .Y(_16387_));
 sky130_fd_sc_hd__inv_2 _43465_ (.A(_16387_),
    .Y(_16388_));
 sky130_fd_sc_hd__a21bo_1 _43466_ (.A1(_15669_),
    .A2(_13634_),
    .B1_N(_08741_),
    .X(_16389_));
 sky130_fd_sc_hd__nor3b_2 _43467_ (.A(_16389_),
    .B(_15670_),
    .C_N(_15666_),
    .Y(_16390_));
 sky130_fd_sc_hd__buf_2 _43468_ (.A(_12179_),
    .X(_16391_));
 sky130_fd_sc_hd__and4b_1 _43469_ (.A_N(_15664_),
    .B(_07425_),
    .C(_15669_),
    .D(_16391_),
    .X(_16392_));
 sky130_fd_sc_hd__o211a_1 _43470_ (.A1(_16390_),
    .A2(_16392_),
    .B1(_15673_),
    .C1(_15677_),
    .X(_16394_));
 sky130_fd_sc_hd__a21oi_4 _43471_ (.A1(_15673_),
    .A2(_15677_),
    .B1(_16390_),
    .Y(_16395_));
 sky130_fd_sc_hd__a31o_1 _43472_ (.A1(_15013_),
    .A2(_15014_),
    .A3(_12236_),
    .B1(_15680_),
    .X(_16396_));
 sky130_fd_sc_hd__a31o_1 _43473_ (.A1(_15678_),
    .A2(_15016_),
    .A3(_15017_),
    .B1(_16396_),
    .X(_16397_));
 sky130_fd_sc_hd__a21bo_1 _43474_ (.A1(_15685_),
    .A2(_15687_),
    .B1_N(_15686_),
    .X(_16398_));
 sky130_fd_sc_hd__xnor2_2 _43475_ (.A(_16397_),
    .B(_16398_),
    .Y(_16399_));
 sky130_fd_sc_hd__o21ba_1 _43476_ (.A1(_15691_),
    .A2(_15694_),
    .B1_N(_15692_),
    .X(_16400_));
 sky130_fd_sc_hd__xnor2_2 _43477_ (.A(_16399_),
    .B(_16400_),
    .Y(_16401_));
 sky130_fd_sc_hd__nor3_4 _43478_ (.A(_16394_),
    .B(_16395_),
    .C(_16401_),
    .Y(_16402_));
 sky130_fd_sc_hd__o21ai_2 _43479_ (.A1(_16394_),
    .A2(_16395_),
    .B1(_16401_),
    .Y(_16403_));
 sky130_fd_sc_hd__and2b_1 _43480_ (.A_N(_16402_),
    .B(_16403_),
    .X(_16405_));
 sky130_fd_sc_hd__o21a_1 _43481_ (.A1(_15705_),
    .A2(_15706_),
    .B1(_15707_),
    .X(_16406_));
 sky130_fd_sc_hd__a21oi_1 _43482_ (.A1(_15705_),
    .A2(_15706_),
    .B1(_15707_),
    .Y(_16407_));
 sky130_fd_sc_hd__o21ai_1 _43483_ (.A1(_07330_),
    .A2(_07331_),
    .B1(_05603_),
    .Y(_16408_));
 sky130_fd_sc_hd__o211a_1 _43484_ (.A1(_16406_),
    .A2(_16407_),
    .B1(_16408_),
    .C1(_15700_),
    .X(_16409_));
 sky130_fd_sc_hd__and4bb_1 _43485_ (.A_N(_15705_),
    .B_N(_15706_),
    .C(_15707_),
    .D(_14469_),
    .X(_16410_));
 sky130_fd_sc_hd__a211o_1 _43486_ (.A1(_15708_),
    .A2(_15711_),
    .B1(_16409_),
    .C1(_16410_),
    .X(_16411_));
 sky130_fd_sc_hd__a31o_1 _43487_ (.A1(_15705_),
    .A2(_15706_),
    .A3(_15707_),
    .B1(_15702_),
    .X(_16412_));
 sky130_fd_sc_hd__o221ai_2 _43488_ (.A1(_16412_),
    .A2(_15703_),
    .B1(_16409_),
    .B2(_16410_),
    .C1(_15711_),
    .Y(_16413_));
 sky130_fd_sc_hd__nand2_1 _43489_ (.A(_16411_),
    .B(_16413_),
    .Y(_16414_));
 sky130_fd_sc_hd__xor2_2 _43490_ (.A(_16405_),
    .B(_16414_),
    .X(_16416_));
 sky130_fd_sc_hd__a21boi_2 _43491_ (.A1(_16386_),
    .A2(_16388_),
    .B1_N(_16416_),
    .Y(_16417_));
 sky130_fd_sc_hd__nor3b_4 _43492_ (.A(_16416_),
    .B(_16387_),
    .C_N(_16386_),
    .Y(_16418_));
 sky130_fd_sc_hd__a211o_4 _43493_ (.A1(_15659_),
    .A2(_16368_),
    .B1(_16417_),
    .C1(_16418_),
    .X(_16419_));
 sky130_fd_sc_hd__o221ai_4 _43494_ (.A1(_15661_),
    .A2(_15658_),
    .B1(_16417_),
    .B2(_16418_),
    .C1(_16368_),
    .Y(_16420_));
 sky130_fd_sc_hd__nand2_1 _43495_ (.A(_16419_),
    .B(net64),
    .Y(_16421_));
 sky130_fd_sc_hd__and2b_1 _43496_ (.A_N(_16367_),
    .B(net64),
    .X(_16422_));
 sky130_fd_sc_hd__a21oi_2 _43497_ (.A1(_15759_),
    .A2(_15760_),
    .B1(net65),
    .Y(_16423_));
 sky130_fd_sc_hd__a221o_1 _43498_ (.A1(_16367_),
    .A2(_16421_),
    .B1(_16422_),
    .B2(_16419_),
    .C1(_16423_),
    .X(_16424_));
 sky130_fd_sc_hd__a22o_1 _43499_ (.A1(_16367_),
    .A2(_16421_),
    .B1(_16422_),
    .B2(_16419_),
    .X(_16425_));
 sky130_fd_sc_hd__nand2_1 _43500_ (.A(_16425_),
    .B(_16423_),
    .Y(_16427_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43501_ (.A(_15803_),
    .X(_16428_));
 sky130_fd_sc_hd__or3_1 _43502_ (.A(_15770_),
    .B(_15791_),
    .C(_15792_),
    .X(_16429_));
 sky130_fd_sc_hd__o21a_1 _43503_ (.A1(_15794_),
    .A2(_16428_),
    .B1(_16429_),
    .X(_16430_));
 sky130_fd_sc_hd__a2bb2o_1 _43504_ (.A1_N(_14878_),
    .A2_N(_15780_),
    .B1(_15776_),
    .B2(_12588_),
    .X(_16431_));
 sky130_fd_sc_hd__o31ai_2 _43505_ (.A1(_15781_),
    .A2(_15783_),
    .A3(_15780_),
    .B1(_16431_),
    .Y(_16432_));
 sky130_fd_sc_hd__and2_1 _43506_ (.A(_15785_),
    .B(_15786_),
    .X(_16433_));
 sky130_fd_sc_hd__o21ai_2 _43507_ (.A1(_16432_),
    .A2(_16433_),
    .B1(_15771_),
    .Y(_16434_));
 sky130_fd_sc_hd__or3_1 _43508_ (.A(_15771_),
    .B(_16432_),
    .C(_16433_),
    .X(_16435_));
 sky130_fd_sc_hd__a21o_1 _43509_ (.A1(_16434_),
    .A2(_16435_),
    .B1(_15769_),
    .X(_16436_));
 sky130_fd_sc_hd__nand3_1 _43510_ (.A(_16435_),
    .B(_15769_),
    .C(_16434_),
    .Y(_16438_));
 sky130_fd_sc_hd__nand2_1 _43511_ (.A(_16436_),
    .B(_16438_),
    .Y(_16439_));
 sky130_fd_sc_hd__a21boi_1 _43512_ (.A1(_15790_),
    .A2(_15769_),
    .B1_N(_15788_),
    .Y(_16440_));
 sky130_fd_sc_hd__xnor2_1 _43513_ (.A(_16439_),
    .B(_16440_),
    .Y(_16441_));
 sky130_fd_sc_hd__nand2_1 _43514_ (.A(_16428_),
    .B(_16441_),
    .Y(_16442_));
 sky130_fd_sc_hd__or2_1 _43515_ (.A(_15803_),
    .B(_16441_),
    .X(_16443_));
 sky130_fd_sc_hd__o21a_1 _43516_ (.A1(net78),
    .A2(_15757_),
    .B1(_15720_),
    .X(_16444_));
 sky130_fd_sc_hd__a21o_1 _43517_ (.A1(net78),
    .A2(_15757_),
    .B1(_16444_),
    .X(_16445_));
 sky130_fd_sc_hd__a21oi_1 _43518_ (.A1(_16442_),
    .A2(_16443_),
    .B1(_16445_),
    .Y(_16446_));
 sky130_fd_sc_hd__nand3_1 _43519_ (.A(_16445_),
    .B(_16442_),
    .C(_16443_),
    .Y(_16447_));
 sky130_fd_sc_hd__or2b_1 _43520_ (.A(_16446_),
    .B_N(_16447_),
    .X(_16449_));
 sky130_fd_sc_hd__xnor2_1 _43521_ (.A(_16430_),
    .B(_16449_),
    .Y(_16450_));
 sky130_fd_sc_hd__a21boi_1 _43522_ (.A1(_16424_),
    .A2(_16427_),
    .B1_N(_16450_),
    .Y(_16451_));
 sky130_fd_sc_hd__and3b_1 _43523_ (.A_N(_16450_),
    .B(_16424_),
    .C(_16427_),
    .X(_16452_));
 sky130_fd_sc_hd__o221ai_1 _43524_ (.A1(_15765_),
    .A2(_15808_),
    .B1(_16451_),
    .B2(_16452_),
    .C1(_15810_),
    .Y(_16453_));
 sky130_fd_sc_hd__a211o_1 _43525_ (.A1(_15810_),
    .A2(_15809_),
    .B1(_16451_),
    .C1(_16452_),
    .X(_16454_));
 sky130_fd_sc_hd__nand2_1 _43526_ (.A(_16453_),
    .B(_16454_),
    .Y(_16455_));
 sky130_fd_sc_hd__a2bb2o_4 _43527_ (.A1_N(_15797_),
    .A2_N(_15801_),
    .B1(_15798_),
    .B2(_15799_),
    .X(_16456_));
 sky130_fd_sc_hd__and3_1 _43528_ (.A(_14839_),
    .B(_15611_),
    .C(_15612_),
    .X(_16457_));
 sky130_fd_sc_hd__o211a_1 _43529_ (.A1(_15607_),
    .A2(_14827_),
    .B1(_15615_),
    .C1(_15609_),
    .X(_16458_));
 sky130_fd_sc_hd__a21o_1 _43530_ (.A1(_14842_),
    .A2(_16457_),
    .B1(_16458_),
    .X(_16460_));
 sky130_fd_sc_hd__xnor2_4 _43531_ (.A(_16456_),
    .B(_16460_),
    .Y(_16461_));
 sky130_fd_sc_hd__inv_2 _43532_ (.A(_15621_),
    .Y(_16462_));
 sky130_fd_sc_hd__a21o_2 _43533_ (.A1(_16462_),
    .A2(_15619_),
    .B1(_15618_),
    .X(_16463_));
 sky130_fd_sc_hd__nor2_1 _43534_ (.A(_16461_),
    .B(_16463_),
    .Y(_16464_));
 sky130_fd_sc_hd__nand2_1 _43535_ (.A(_16463_),
    .B(_16461_),
    .Y(_16465_));
 sky130_fd_sc_hd__or2b_1 _43536_ (.A(_16464_),
    .B_N(_16465_),
    .X(_16466_));
 sky130_fd_sc_hd__xor2_2 _43537_ (.A(_14861_),
    .B(_16466_),
    .X(_16467_));
 sky130_fd_sc_hd__a31o_1 _43538_ (.A1(_15136_),
    .A2(_15768_),
    .A3(_15804_),
    .B1(_15766_),
    .X(_16468_));
 sky130_fd_sc_hd__nand2_1 _43539_ (.A(_15805_),
    .B(_16468_),
    .Y(_16469_));
 sky130_fd_sc_hd__nand2_1 _43540_ (.A(_16467_),
    .B(_16469_),
    .Y(_16471_));
 sky130_fd_sc_hd__or2_1 _43541_ (.A(_16469_),
    .B(_16467_),
    .X(_16472_));
 sky130_fd_sc_hd__o2bb2a_1 _43542_ (.A1_N(_15625_),
    .A2_N(_15606_),
    .B1(_14861_),
    .B2(_15626_),
    .X(_16473_));
 sky130_fd_sc_hd__o21bai_2 _43543_ (.A1(_16469_),
    .A2(_16467_),
    .B1_N(_16473_),
    .Y(_16474_));
 sky130_fd_sc_hd__a21oi_1 _43544_ (.A1(_16471_),
    .A2(_16472_),
    .B1(_16473_),
    .Y(_16475_));
 sky130_fd_sc_hd__a31oi_2 _43545_ (.A1(_16471_),
    .A2(_16472_),
    .A3(_16474_),
    .B1(_16475_),
    .Y(_16476_));
 sky130_fd_sc_hd__xor2_1 _43546_ (.A(_16455_),
    .B(_16476_),
    .X(_16477_));
 sky130_fd_sc_hd__nand2_1 _43547_ (.A(_16339_),
    .B(_16477_),
    .Y(_16478_));
 sky130_fd_sc_hd__inv_2 _43548_ (.A(_16478_),
    .Y(_16479_));
 sky130_fd_sc_hd__nor2_1 _43549_ (.A(_16477_),
    .B(_16339_),
    .Y(_16480_));
 sky130_fd_sc_hd__nor2_1 _43550_ (.A(_16479_),
    .B(_16480_),
    .Y(_16482_));
 sky130_fd_sc_hd__o211a_1 _43551_ (.A1(_16035_),
    .A2(_16051_),
    .B1(_16060_),
    .C1(_16054_),
    .X(_16483_));
 sky130_fd_sc_hd__clkbuf_2 _43552_ (.A(_16329_),
    .X(_16484_));
 sky130_fd_sc_hd__o211ai_1 _43553_ (.A1(_16036_),
    .A2(_16483_),
    .B1(_16484_),
    .C1(_16334_),
    .Y(_16485_));
 sky130_fd_sc_hd__nand3_1 _43554_ (.A(_16336_),
    .B(_16482_),
    .C(_16485_),
    .Y(_16486_));
 sky130_fd_sc_hd__o211a_1 _43555_ (.A1(_16036_),
    .A2(_16483_),
    .B1(_16484_),
    .C1(_16334_),
    .X(_16487_));
 sky130_fd_sc_hd__a21oi_1 _43556_ (.A1(_16484_),
    .A2(_16334_),
    .B1(_16335_),
    .Y(_16488_));
 sky130_fd_sc_hd__o22ai_2 _43557_ (.A1(_16479_),
    .A2(_16480_),
    .B1(_16487_),
    .B2(_16488_),
    .Y(_16489_));
 sky130_fd_sc_hd__a31o_1 _43558_ (.A1(_16070_),
    .A2(_16071_),
    .A3(_16072_),
    .B1(_15823_),
    .X(_16490_));
 sky130_fd_sc_hd__a21o_1 _43559_ (.A1(_16486_),
    .A2(_16489_),
    .B1(_16490_),
    .X(_16491_));
 sky130_fd_sc_hd__a31o_1 _43560_ (.A1(_16048_),
    .A2(_16050_),
    .A3(_16055_),
    .B1(_16066_),
    .X(_16493_));
 sky130_fd_sc_hd__o21a_1 _43561_ (.A1(_10321_),
    .A2(_09004_),
    .B1(_10435_),
    .X(_16494_));
 sky130_fd_sc_hd__nand2_1 _43562_ (.A(_15577_),
    .B(_16494_),
    .Y(_16495_));
 sky130_fd_sc_hd__or2_1 _43563_ (.A(_15576_),
    .B(_16494_),
    .X(_16496_));
 sky130_fd_sc_hd__a21oi_1 _43564_ (.A1(_16495_),
    .A2(_16496_),
    .B1(_15501_),
    .Y(_16497_));
 sky130_fd_sc_hd__and3_1 _43565_ (.A(_16496_),
    .B(_15501_),
    .C(_16495_),
    .X(_16498_));
 sky130_fd_sc_hd__or2_2 _43566_ (.A(_16497_),
    .B(_16498_),
    .X(_16499_));
 sky130_fd_sc_hd__clkbuf_2 _43567_ (.A(_15566_),
    .X(_16500_));
 sky130_fd_sc_hd__clkbuf_2 _43568_ (.A(_13296_),
    .X(_16501_));
 sky130_fd_sc_hd__o21a_1 _43569_ (.A1(_16044_),
    .A2(_05101_),
    .B1(_16501_),
    .X(_16502_));
 sky130_fd_sc_hd__a221oi_1 _43570_ (.A1(_16323_),
    .A2(_16044_),
    .B1(_15443_),
    .B2(_16500_),
    .C1(_16502_),
    .Y(_16504_));
 sky130_fd_sc_hd__and3_1 _43571_ (.A(_16323_),
    .B(_16321_),
    .C(_14259_),
    .X(_16505_));
 sky130_fd_sc_hd__o221a_1 _43572_ (.A1(_16321_),
    .A2(_03566_),
    .B1(_16505_),
    .B2(_16502_),
    .C1(_16500_),
    .X(_16506_));
 sky130_fd_sc_hd__clkbuf_2 _43573_ (.A(_16059_),
    .X(_16507_));
 sky130_fd_sc_hd__o21ai_1 _43574_ (.A1(_16507_),
    .A2(_15445_),
    .B1(_15565_),
    .Y(_16508_));
 sky130_fd_sc_hd__clkbuf_2 _43575_ (.A(_15570_),
    .X(_16509_));
 sky130_fd_sc_hd__and4bb_1 _43576_ (.A_N(_16504_),
    .B_N(_16506_),
    .C(_16508_),
    .D(_16509_),
    .X(_16510_));
 sky130_fd_sc_hd__o2bb2a_1 _43577_ (.A1_N(_16508_),
    .A2_N(_16509_),
    .B1(_16504_),
    .B2(_16506_),
    .X(_16511_));
 sky130_fd_sc_hd__or2_1 _43578_ (.A(_16510_),
    .B(_16511_),
    .X(_16512_));
 sky130_fd_sc_hd__xnor2_1 _43579_ (.A(_16499_),
    .B(_16512_),
    .Y(_16513_));
 sky130_fd_sc_hd__a21o_1 _43580_ (.A1(_16069_),
    .A2(_16493_),
    .B1(_16513_),
    .X(_16515_));
 sky130_fd_sc_hd__nand3_2 _43581_ (.A(_16069_),
    .B(_16493_),
    .C(_16513_),
    .Y(_16516_));
 sky130_fd_sc_hd__o21a_1 _43582_ (.A1(_15573_),
    .A2(net144),
    .B1(_16516_),
    .X(_16517_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43583_ (.A(_15574_),
    .X(_16518_));
 sky130_fd_sc_hd__buf_2 _43584_ (.A(_16518_),
    .X(_16519_));
 sky130_fd_sc_hd__a41o_1 _43585_ (.A1(_16519_),
    .A2(_15568_),
    .A3(_15571_),
    .A4(_15572_),
    .B1(net144),
    .X(_16520_));
 sky130_fd_sc_hd__a21oi_1 _43586_ (.A1(_16515_),
    .A2(_16516_),
    .B1(_16520_),
    .Y(_16521_));
 sky130_fd_sc_hd__a21oi_1 _43587_ (.A1(_16515_),
    .A2(_16517_),
    .B1(_16521_),
    .Y(_16522_));
 sky130_fd_sc_hd__nand3_1 _43588_ (.A(_16490_),
    .B(_16486_),
    .C(_16489_),
    .Y(_16523_));
 sky130_fd_sc_hd__nand3_1 _43589_ (.A(_16491_),
    .B(_16522_),
    .C(_16523_),
    .Y(_16524_));
 sky130_fd_sc_hd__and3_1 _43590_ (.A(_16520_),
    .B(_16515_),
    .C(_16516_),
    .X(_16526_));
 sky130_fd_sc_hd__and3_1 _43591_ (.A(_16490_),
    .B(_16486_),
    .C(_16489_),
    .X(_16527_));
 sky130_fd_sc_hd__a21oi_1 _43592_ (.A1(_16486_),
    .A2(_16489_),
    .B1(_16490_),
    .Y(_16528_));
 sky130_fd_sc_hd__o22ai_1 _43593_ (.A1(_16521_),
    .A2(_16526_),
    .B1(_16527_),
    .B2(_16528_),
    .Y(_16529_));
 sky130_fd_sc_hd__nand3b_1 _43594_ (.A_N(_16166_),
    .B(_16524_),
    .C(_16529_),
    .Y(_16530_));
 sky130_fd_sc_hd__o21ai_1 _43595_ (.A1(_16527_),
    .A2(_16528_),
    .B1(_16522_),
    .Y(_16531_));
 sky130_fd_sc_hd__o211ai_1 _43596_ (.A1(_16521_),
    .A2(_16526_),
    .B1(_16523_),
    .C1(_16491_),
    .Y(_16532_));
 sky130_fd_sc_hd__nand3_1 _43597_ (.A(_16531_),
    .B(_16532_),
    .C(_16166_),
    .Y(_16533_));
 sky130_fd_sc_hd__nand2_1 _43598_ (.A(_16530_),
    .B(_16533_),
    .Y(_16534_));
 sky130_fd_sc_hd__nand2_1 _43599_ (.A(_16165_),
    .B(_16534_),
    .Y(_16535_));
 sky130_fd_sc_hd__nand3b_1 _43600_ (.A_N(_16165_),
    .B(_16530_),
    .C(_16533_),
    .Y(_16537_));
 sky130_fd_sc_hd__a32o_1 _43601_ (.A1(_15564_),
    .A2(_16080_),
    .A3(_16084_),
    .B1(_16092_),
    .B2(_16121_),
    .X(_16538_));
 sky130_fd_sc_hd__a21o_1 _43602_ (.A1(_16535_),
    .A2(_16537_),
    .B1(_16538_),
    .X(_16539_));
 sky130_fd_sc_hd__nand3_1 _43603_ (.A(_16538_),
    .B(_16535_),
    .C(_16537_),
    .Y(_16540_));
 sky130_fd_sc_hd__a21boi_2 _43604_ (.A1(_14812_),
    .A2(_16117_),
    .B1_N(_16116_),
    .Y(_16541_));
 sky130_fd_sc_hd__a21bo_1 _43605_ (.A1(_16539_),
    .A2(_16540_),
    .B1_N(_16541_),
    .X(_16542_));
 sky130_fd_sc_hd__nand3b_1 _43606_ (.A_N(_16541_),
    .B(_16539_),
    .C(_16540_),
    .Y(_16543_));
 sky130_fd_sc_hd__o21ai_1 _43607_ (.A1(_15541_),
    .A2(_16135_),
    .B1(_16128_),
    .Y(_16544_));
 sky130_fd_sc_hd__a21oi_1 _43608_ (.A1(_16542_),
    .A2(_16543_),
    .B1(_16544_),
    .Y(_16545_));
 sky130_fd_sc_hd__and3_1 _43609_ (.A(_16544_),
    .B(_16542_),
    .C(_16543_),
    .X(_16546_));
 sky130_fd_sc_hd__nor2_1 _43610_ (.A(_16545_),
    .B(_16546_),
    .Y(_16548_));
 sky130_fd_sc_hd__nand4_2 _43611_ (.A(_15556_),
    .B(_15561_),
    .C(_16140_),
    .D(_13924_),
    .Y(_16549_));
 sky130_fd_sc_hd__inv_2 _43612_ (.A(_16139_),
    .Y(_16550_));
 sky130_fd_sc_hd__nand3_1 _43613_ (.A(_16138_),
    .B(_16137_),
    .C(_16129_),
    .Y(_16551_));
 sky130_fd_sc_hd__nand2_1 _43614_ (.A(_15555_),
    .B(_16551_),
    .Y(_16552_));
 sky130_fd_sc_hd__nor2_1 _43615_ (.A(_14776_),
    .B(_14778_),
    .Y(_16553_));
 sky130_fd_sc_hd__clkinvlp_2 _43616_ (.A(_14780_),
    .Y(_16554_));
 sky130_fd_sc_hd__o2111a_1 _43617_ (.A1(_16553_),
    .A2(_16554_),
    .B1(_15555_),
    .C1(_15552_),
    .D1(_15560_),
    .X(_16555_));
 sky130_fd_sc_hd__a22oi_2 _43618_ (.A1(_16550_),
    .A2(_16552_),
    .B1(_16555_),
    .B2(_16140_),
    .Y(_16556_));
 sky130_fd_sc_hd__nand3_1 _43619_ (.A(_09107_),
    .B(_10415_),
    .C(_10420_),
    .Y(_16557_));
 sky130_fd_sc_hd__nand4b_1 _43620_ (.A_N(_16557_),
    .B(_09106_),
    .C(_11690_),
    .D(_12871_),
    .Y(_16559_));
 sky130_fd_sc_hd__a21oi_2 _43621_ (.A1(_07632_),
    .A2(_07638_),
    .B1(_16559_),
    .Y(_16560_));
 sky130_fd_sc_hd__nand4_2 _43622_ (.A(_16560_),
    .B(_15556_),
    .C(_15561_),
    .D(_16140_),
    .Y(_16561_));
 sky130_fd_sc_hd__and4b_1 _43623_ (.A_N(_16548_),
    .B(_16549_),
    .C(_16556_),
    .D(_16561_),
    .X(_16562_));
 sky130_fd_sc_hd__a311oi_2 _43624_ (.A1(_16556_),
    .A2(_16561_),
    .A3(_16549_),
    .B1(_16546_),
    .C1(_16545_),
    .Y(_16563_));
 sky130_fd_sc_hd__nor2_1 _43625_ (.A(_16562_),
    .B(_16563_),
    .Y(_00018_));
 sky130_fd_sc_hd__nand3_1 _43626_ (.A(_16556_),
    .B(_16561_),
    .C(_16549_),
    .Y(_16564_));
 sky130_fd_sc_hd__a21oi_1 _43627_ (.A1(_16564_),
    .A2(_16548_),
    .B1(_16546_),
    .Y(_16565_));
 sky130_fd_sc_hd__a21oi_1 _43628_ (.A1(_16535_),
    .A2(_16537_),
    .B1(_16538_),
    .Y(_16566_));
 sky130_fd_sc_hd__a311o_2 _43629_ (.A1(_16142_),
    .A2(_16143_),
    .A3(_16159_),
    .B1(_16114_),
    .C1(_16094_),
    .X(_16567_));
 sky130_fd_sc_hd__a21o_1 _43630_ (.A1(_16491_),
    .A2(_16522_),
    .B1(_16527_),
    .X(_16569_));
 sky130_fd_sc_hd__nand2_1 _43631_ (.A(_16312_),
    .B(_16313_),
    .Y(_16570_));
 sky130_fd_sc_hd__nor2_1 _43632_ (.A(_12876_),
    .B(_16303_),
    .Y(_16571_));
 sky130_fd_sc_hd__clkbuf_2 _43633_ (.A(_16292_),
    .X(_16572_));
 sky130_fd_sc_hd__o21ba_1 _43634_ (.A1(_16256_),
    .A2(_16274_),
    .B1_N(_16273_),
    .X(_16573_));
 sky130_fd_sc_hd__o21a_1 _43635_ (.A1(_15299_),
    .A2(_15304_),
    .B1(_13209_),
    .X(_16574_));
 sky130_fd_sc_hd__buf_1 _43636_ (.A(_15294_),
    .X(_16575_));
 sky130_fd_sc_hd__o221a_1 _43637_ (.A1(_16257_),
    .A2(_15370_),
    .B1(_16575_),
    .B2(_16221_),
    .C1(_16222_),
    .X(_16576_));
 sky130_fd_sc_hd__o211ai_2 _43638_ (.A1(_15299_),
    .A2(_15304_),
    .B1(_16230_),
    .C1(_16231_),
    .Y(_16577_));
 sky130_fd_sc_hd__o211a_1 _43639_ (.A1(_16574_),
    .A2(_16576_),
    .B1(_16231_),
    .C1(_16577_),
    .X(_16578_));
 sky130_fd_sc_hd__a211oi_2 _43640_ (.A1(_16231_),
    .A2(_16577_),
    .B1(_16574_),
    .C1(_16576_),
    .Y(_16580_));
 sky130_fd_sc_hd__nor3_1 _43641_ (.A(_16259_),
    .B(_16578_),
    .C(_16580_),
    .Y(_16581_));
 sky130_fd_sc_hd__o21a_1 _43642_ (.A1(_16578_),
    .A2(_16580_),
    .B1(_16259_),
    .X(_16582_));
 sky130_fd_sc_hd__and2_1 _43643_ (.A(_16262_),
    .B(_16264_),
    .X(_16583_));
 sky130_fd_sc_hd__o21ai_1 _43644_ (.A1(net124),
    .A2(_16582_),
    .B1(_16583_),
    .Y(_16584_));
 sky130_fd_sc_hd__or3_1 _43645_ (.A(net124),
    .B(_16582_),
    .C(_16583_),
    .X(_16585_));
 sky130_fd_sc_hd__a211oi_2 _43646_ (.A1(_16584_),
    .A2(_16585_),
    .B1(_16247_),
    .C1(_16249_),
    .Y(_16586_));
 sky130_fd_sc_hd__o211a_1 _43647_ (.A1(_16247_),
    .A2(_16249_),
    .B1(_16584_),
    .C1(_16585_),
    .X(_16587_));
 sky130_fd_sc_hd__or3_1 _43648_ (.A(_16269_),
    .B(_16586_),
    .C(_16587_),
    .X(_16588_));
 sky130_fd_sc_hd__o21ai_1 _43649_ (.A1(_16586_),
    .A2(_16587_),
    .B1(_16269_),
    .Y(_16589_));
 sky130_fd_sc_hd__and2b_1 _43650_ (.A_N(_16241_),
    .B(_16243_),
    .X(_16591_));
 sky130_fd_sc_hd__a2bb2o_1 _43651_ (.A1_N(_15874_),
    .A2_N(_15875_),
    .B1(_16234_),
    .B2(_16235_),
    .X(_16592_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43652_ (.A(_15867_),
    .X(_16593_));
 sky130_fd_sc_hd__nand2_2 _43653_ (.A(_16200_),
    .B(_15867_),
    .Y(_16594_));
 sky130_fd_sc_hd__o21a_1 _43654_ (.A1(_13045_),
    .A2(_16594_),
    .B1(_16202_),
    .X(_16595_));
 sky130_fd_sc_hd__a31o_1 _43655_ (.A1(_16200_),
    .A2(_16593_),
    .A3(_16199_),
    .B1(_16595_),
    .X(_16596_));
 sky130_fd_sc_hd__nor2b_2 _43656_ (.A(_16596_),
    .B_N(_16234_),
    .Y(_16597_));
 sky130_fd_sc_hd__o211a_1 _43657_ (.A1(_16221_),
    .A2(_15926_),
    .B1(_16203_),
    .C1(_16596_),
    .X(_16598_));
 sky130_fd_sc_hd__a211o_1 _43658_ (.A1(_16592_),
    .A2(_16238_),
    .B1(_16597_),
    .C1(_16598_),
    .X(_16599_));
 sky130_fd_sc_hd__or3b_1 _43659_ (.A(_15332_),
    .B(_16593_),
    .C_N(_13161_),
    .X(_16600_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43660_ (.A(_13140_),
    .X(_16602_));
 sky130_fd_sc_hd__o311a_1 _43661_ (.A1(_16225_),
    .A2(_16224_),
    .A3(_15929_),
    .B1(_16600_),
    .C1(_16602_),
    .X(_16603_));
 sky130_fd_sc_hd__a21oi_1 _43662_ (.A1(_16600_),
    .A2(_16602_),
    .B1(_15928_),
    .Y(_16604_));
 sky130_fd_sc_hd__a21oi_1 _43663_ (.A1(_16603_),
    .A2(_16223_),
    .B1(_16604_),
    .Y(_16605_));
 sky130_fd_sc_hd__o211ai_2 _43664_ (.A1(_16597_),
    .A2(_16598_),
    .B1(_16592_),
    .C1(_16238_),
    .Y(_16606_));
 sky130_fd_sc_hd__and3_1 _43665_ (.A(_16599_),
    .B(_16605_),
    .C(_16606_),
    .X(_16607_));
 sky130_fd_sc_hd__a21oi_1 _43666_ (.A1(_16606_),
    .A2(_16599_),
    .B1(_16605_),
    .Y(_16608_));
 sky130_fd_sc_hd__or2_1 _43667_ (.A(_16607_),
    .B(_16608_),
    .X(_16609_));
 sky130_fd_sc_hd__a21oi_2 _43668_ (.A1(_15851_),
    .A2(_16208_),
    .B1(_16211_),
    .Y(_16610_));
 sky130_fd_sc_hd__xnor2_1 _43669_ (.A(_16609_),
    .B(_16610_),
    .Y(_16611_));
 sky130_fd_sc_hd__nand2_1 _43670_ (.A(_16591_),
    .B(_16611_),
    .Y(_16613_));
 sky130_fd_sc_hd__or2_1 _43671_ (.A(_16611_),
    .B(_16591_),
    .X(_16614_));
 sky130_fd_sc_hd__and2_1 _43672_ (.A(_16613_),
    .B(_16614_),
    .X(_16615_));
 sky130_fd_sc_hd__clkbuf_2 _43673_ (.A(_16200_),
    .X(_16616_));
 sky130_fd_sc_hd__or2_1 _43674_ (.A(_16616_),
    .B(_15881_),
    .X(_16617_));
 sky130_fd_sc_hd__a21o_1 _43675_ (.A1(_16594_),
    .A2(_16617_),
    .B1(_16198_),
    .X(_16618_));
 sky130_fd_sc_hd__o211ai_4 _43676_ (.A1(_15881_),
    .A2(_16616_),
    .B1(_16594_),
    .C1(_16198_),
    .Y(_16619_));
 sky130_fd_sc_hd__and3_1 _43677_ (.A(_16618_),
    .B(_16188_),
    .C(_16619_),
    .X(_16620_));
 sky130_fd_sc_hd__a21oi_1 _43678_ (.A1(_16619_),
    .A2(_16618_),
    .B1(_16188_),
    .Y(_16621_));
 sky130_fd_sc_hd__o21ba_1 _43679_ (.A1(_16198_),
    .A2(_16204_),
    .B1_N(_16196_),
    .X(_16622_));
 sky130_fd_sc_hd__o21ai_2 _43680_ (.A1(_16620_),
    .A2(_16621_),
    .B1(_16622_),
    .Y(_16624_));
 sky130_fd_sc_hd__or3_2 _43681_ (.A(_16622_),
    .B(_16620_),
    .C(_16621_),
    .X(_16625_));
 sky130_fd_sc_hd__nand2_1 _43682_ (.A(_16624_),
    .B(_16625_),
    .Y(_16626_));
 sky130_fd_sc_hd__a21oi_4 _43683_ (.A1(_15193_),
    .A2(_16180_),
    .B1(_16183_),
    .Y(_16627_));
 sky130_fd_sc_hd__a2bb2o_2 _43684_ (.A1_N(_11804_),
    .A2_N(_13945_),
    .B1(_15829_),
    .B2(_13980_),
    .X(_16628_));
 sky130_fd_sc_hd__o2bb2a_1 _43685_ (.A1_N(_15828_),
    .A2_N(_15831_),
    .B1(_13980_),
    .B2(_15834_),
    .X(_16629_));
 sky130_fd_sc_hd__xnor2_1 _43686_ (.A(_16628_),
    .B(_16629_),
    .Y(_16630_));
 sky130_fd_sc_hd__nand2_2 _43687_ (.A(_16191_),
    .B(_16630_),
    .Y(_16631_));
 sky130_fd_sc_hd__a21o_1 _43688_ (.A1(_16189_),
    .A2(_16186_),
    .B1(_16627_),
    .X(_16632_));
 sky130_fd_sc_hd__xor2_2 _43689_ (.A(_16628_),
    .B(_16629_),
    .X(_16633_));
 sky130_fd_sc_hd__nand2_2 _43690_ (.A(_16632_),
    .B(_16633_),
    .Y(_16635_));
 sky130_fd_sc_hd__o21ai_1 _43691_ (.A1(_16627_),
    .A2(_16631_),
    .B1(_16635_),
    .Y(_16636_));
 sky130_fd_sc_hd__nand2_1 _43692_ (.A(_16626_),
    .B(_16636_),
    .Y(_16637_));
 sky130_fd_sc_hd__o2111ai_4 _43693_ (.A1(_16627_),
    .A2(_16631_),
    .B1(_16635_),
    .C1(_16625_),
    .D1(_16624_),
    .Y(_16638_));
 sky130_fd_sc_hd__o21ba_1 _43694_ (.A1(_15839_),
    .A2(_16179_),
    .B1_N(_16192_),
    .X(_16639_));
 sky130_fd_sc_hd__a221oi_2 _43695_ (.A1(_16212_),
    .A2(_16194_),
    .B1(_16637_),
    .B2(_16638_),
    .C1(_16639_),
    .Y(_16640_));
 sky130_fd_sc_hd__nand2_1 _43696_ (.A(_16194_),
    .B(_16212_),
    .Y(_16641_));
 sky130_fd_sc_hd__nand2_1 _43697_ (.A(_16637_),
    .B(_16638_),
    .Y(_16642_));
 sky130_fd_sc_hd__a21oi_2 _43698_ (.A1(_16193_),
    .A2(_16641_),
    .B1(_16642_),
    .Y(_16643_));
 sky130_fd_sc_hd__nor3_1 _43699_ (.A(_16615_),
    .B(_16640_),
    .C(_16643_),
    .Y(_16644_));
 sky130_fd_sc_hd__o21a_1 _43700_ (.A1(_16640_),
    .A2(_16643_),
    .B1(_16615_),
    .X(_16646_));
 sky130_fd_sc_hd__nor2_1 _43701_ (.A(_16644_),
    .B(_16646_),
    .Y(_16647_));
 sky130_fd_sc_hd__a21o_1 _43702_ (.A1(_16219_),
    .A2(_16253_),
    .B1(_16647_),
    .X(_16648_));
 sky130_fd_sc_hd__nand3_1 _43703_ (.A(_16219_),
    .B(_16253_),
    .C(_16647_),
    .Y(_16649_));
 sky130_fd_sc_hd__a22oi_2 _43704_ (.A1(_16588_),
    .A2(_16589_),
    .B1(_16648_),
    .B2(_16649_),
    .Y(_16650_));
 sky130_fd_sc_hd__and4_1 _43705_ (.A(_16588_),
    .B(_16589_),
    .C(_16648_),
    .D(_16649_),
    .X(_16651_));
 sky130_fd_sc_hd__o21a_1 _43706_ (.A1(_16178_),
    .A2(_16254_),
    .B1(_16276_),
    .X(_16652_));
 sky130_fd_sc_hd__o21a_1 _43707_ (.A1(_16650_),
    .A2(_16651_),
    .B1(_16652_),
    .X(_16653_));
 sky130_fd_sc_hd__or2_1 _43708_ (.A(_16178_),
    .B(_16254_),
    .X(_16654_));
 sky130_fd_sc_hd__a211oi_2 _43709_ (.A1(_16654_),
    .A2(_16276_),
    .B1(_16650_),
    .C1(_16651_),
    .Y(_16655_));
 sky130_fd_sc_hd__or3_2 _43710_ (.A(_16573_),
    .B(_16653_),
    .C(_16655_),
    .X(_16657_));
 sky130_fd_sc_hd__o21ai_2 _43711_ (.A1(_16653_),
    .A2(_16655_),
    .B1(_16573_),
    .Y(_16658_));
 sky130_fd_sc_hd__o21a_1 _43712_ (.A1(_16285_),
    .A2(_16282_),
    .B1(_16287_),
    .X(_16659_));
 sky130_fd_sc_hd__a21bo_2 _43713_ (.A1(_16657_),
    .A2(_16658_),
    .B1_N(_16659_),
    .X(_16660_));
 sky130_fd_sc_hd__inv_2 _43714_ (.A(_16660_),
    .Y(_16661_));
 sky130_fd_sc_hd__nand3b_4 _43715_ (.A_N(_16659_),
    .B(_16657_),
    .C(_16658_),
    .Y(_16662_));
 sky130_fd_sc_hd__inv_2 _43716_ (.A(_16662_),
    .Y(_16663_));
 sky130_fd_sc_hd__o2bb2ai_2 _43717_ (.A1_N(_16572_),
    .A2_N(_16300_),
    .B1(_16661_),
    .B2(_16663_),
    .Y(_16664_));
 sky130_fd_sc_hd__nor2_1 _43718_ (.A(_16661_),
    .B(_16663_),
    .Y(_16665_));
 sky130_fd_sc_hd__o211ai_4 _43719_ (.A1(_16290_),
    .A2(_16289_),
    .B1(_16665_),
    .C1(_16300_),
    .Y(_16666_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43720_ (.A(_15414_),
    .X(_16668_));
 sky130_fd_sc_hd__buf_2 _43721_ (.A(_16668_),
    .X(_16669_));
 sky130_fd_sc_hd__a31oi_4 _43722_ (.A1(_16664_),
    .A2(_16666_),
    .A3(_16669_),
    .B1(_16007_),
    .Y(_16670_));
 sky130_fd_sc_hd__buf_2 _43723_ (.A(_15162_),
    .X(_16671_));
 sky130_fd_sc_hd__buf_2 _43724_ (.A(_15164_),
    .X(_16672_));
 sky130_fd_sc_hd__nor2_1 _43725_ (.A(_15404_),
    .B(_15994_),
    .Y(_16673_));
 sky130_fd_sc_hd__and3_1 _43726_ (.A(_16673_),
    .B(_15995_),
    .C(_16176_),
    .X(_16674_));
 sky130_fd_sc_hd__a2bb2oi_2 _43727_ (.A1_N(_15996_),
    .A2_N(_16295_),
    .B1(_16674_),
    .B2(_15168_),
    .Y(_16675_));
 sky130_fd_sc_hd__o221ai_4 _43728_ (.A1(_16661_),
    .A2(_16663_),
    .B1(_16293_),
    .B2(_16675_),
    .C1(_16572_),
    .Y(_16676_));
 sky130_fd_sc_hd__o21ai_1 _43729_ (.A1(_16293_),
    .A2(_16675_),
    .B1(_16572_),
    .Y(_16677_));
 sky130_fd_sc_hd__nand2_1 _43730_ (.A(_16677_),
    .B(_16665_),
    .Y(_16679_));
 sky130_fd_sc_hd__o211ai_4 _43731_ (.A1(_16671_),
    .A2(_16672_),
    .B1(_16676_),
    .C1(_16679_),
    .Y(_16680_));
 sky130_fd_sc_hd__buf_2 _43732_ (.A(_16019_),
    .X(_16681_));
 sky130_fd_sc_hd__nand3_1 _43733_ (.A(_16664_),
    .B(_16666_),
    .C(_16668_),
    .Y(_16682_));
 sky130_fd_sc_hd__a21oi_1 _43734_ (.A1(_16680_),
    .A2(_16682_),
    .B1(_13296_),
    .Y(_16683_));
 sky130_fd_sc_hd__a211oi_1 _43735_ (.A1(_16670_),
    .A2(_16680_),
    .B1(_16681_),
    .C1(_16683_),
    .Y(_16684_));
 sky130_fd_sc_hd__nand2_1 _43736_ (.A(_16670_),
    .B(_16680_),
    .Y(_16685_));
 sky130_fd_sc_hd__a21o_1 _43737_ (.A1(_16680_),
    .A2(_16682_),
    .B1(_13296_),
    .X(_16686_));
 sky130_fd_sc_hd__a21oi_1 _43738_ (.A1(_16685_),
    .A2(_16686_),
    .B1(_16032_),
    .Y(_16687_));
 sky130_fd_sc_hd__o22ai_1 _43739_ (.A1(_16302_),
    .A2(_16571_),
    .B1(_16684_),
    .B2(_16687_),
    .Y(_16688_));
 sky130_fd_sc_hd__o211a_1 _43740_ (.A1(_16671_),
    .A2(_16672_),
    .B1(_16676_),
    .C1(_16679_),
    .X(_16690_));
 sky130_fd_sc_hd__a31o_1 _43741_ (.A1(_16664_),
    .A2(_16666_),
    .A3(_16669_),
    .B1(_16007_),
    .X(_16691_));
 sky130_fd_sc_hd__inv_2 _43742_ (.A(_16022_),
    .Y(_16692_));
 sky130_fd_sc_hd__nand2_1 _43743_ (.A(_16680_),
    .B(_16682_),
    .Y(_16693_));
 sky130_fd_sc_hd__a22oi_1 _43744_ (.A1(_16692_),
    .A2(_16018_),
    .B1(_16693_),
    .B2(_16058_),
    .Y(_16694_));
 sky130_fd_sc_hd__o21ai_1 _43745_ (.A1(_16690_),
    .A2(_16691_),
    .B1(_16694_),
    .Y(_16695_));
 sky130_fd_sc_hd__o2bb2ai_1 _43746_ (.A1_N(_16058_),
    .A2_N(_16693_),
    .B1(_16690_),
    .B2(_16691_),
    .Y(_16696_));
 sky130_fd_sc_hd__nand2_1 _43747_ (.A(_16696_),
    .B(_16681_),
    .Y(_16697_));
 sky130_fd_sc_hd__o2111ai_2 _43748_ (.A1(_16303_),
    .A2(_16059_),
    .B1(_16306_),
    .C1(_16695_),
    .D1(_16697_),
    .Y(_16698_));
 sky130_fd_sc_hd__nand3b_2 _43749_ (.A_N(_16570_),
    .B(_16688_),
    .C(_16698_),
    .Y(_16699_));
 sky130_fd_sc_hd__clkbuf_2 _43750_ (.A(_16699_),
    .X(_16701_));
 sky130_fd_sc_hd__a31o_1 _43751_ (.A1(_16171_),
    .A2(_16297_),
    .A3(_16301_),
    .B1(_16571_),
    .X(_16702_));
 sky130_fd_sc_hd__o21bai_1 _43752_ (.A1(_16684_),
    .A2(_16687_),
    .B1_N(_16702_),
    .Y(_16703_));
 sky130_fd_sc_hd__o211ai_1 _43753_ (.A1(_16302_),
    .A2(_16571_),
    .B1(_16695_),
    .C1(_16697_),
    .Y(_16704_));
 sky130_fd_sc_hd__nand3_1 _43754_ (.A(_16703_),
    .B(_16570_),
    .C(_16704_),
    .Y(_16705_));
 sky130_fd_sc_hd__clkbuf_2 _43755_ (.A(_16705_),
    .X(_16706_));
 sky130_fd_sc_hd__buf_2 _43756_ (.A(_16507_),
    .X(_16707_));
 sky130_fd_sc_hd__nor2_2 _43757_ (.A(_13293_),
    .B(_16707_),
    .Y(_16708_));
 sky130_fd_sc_hd__a21oi_2 _43758_ (.A1(_16701_),
    .A2(_16706_),
    .B1(_16708_),
    .Y(_16709_));
 sky130_fd_sc_hd__inv_2 _43759_ (.A(_16471_),
    .Y(_16710_));
 sky130_fd_sc_hd__inv_2 _43760_ (.A(_16474_),
    .Y(_16712_));
 sky130_fd_sc_hd__nand3_1 _43761_ (.A(_16699_),
    .B(_16706_),
    .C(_16708_),
    .Y(_16713_));
 sky130_fd_sc_hd__o21ai_1 _43762_ (.A1(_16710_),
    .A2(_16712_),
    .B1(_16713_),
    .Y(_16714_));
 sky130_fd_sc_hd__nor2_1 _43763_ (.A(_16709_),
    .B(_16714_),
    .Y(_16715_));
 sky130_fd_sc_hd__clkbuf_2 _43764_ (.A(_16707_),
    .X(_16716_));
 sky130_fd_sc_hd__o2bb2ai_2 _43765_ (.A1_N(_16699_),
    .A2_N(_16706_),
    .B1(_13293_),
    .B2(_16716_),
    .Y(_16717_));
 sky130_fd_sc_hd__a21o_1 _43766_ (.A1(_16469_),
    .A2(_16467_),
    .B1(_16712_),
    .X(_16718_));
 sky130_fd_sc_hd__a21oi_2 _43767_ (.A1(_16717_),
    .A2(_16713_),
    .B1(_16718_),
    .Y(_16719_));
 sky130_fd_sc_hd__a21oi_1 _43768_ (.A1(_16325_),
    .A2(_16320_),
    .B1(_16317_),
    .Y(_16720_));
 sky130_fd_sc_hd__buf_1 _43769_ (.A(_16720_),
    .X(_16721_));
 sky130_fd_sc_hd__o21ai_2 _43770_ (.A1(_16715_),
    .A2(_16719_),
    .B1(_16721_),
    .Y(_16723_));
 sky130_fd_sc_hd__inv_2 _43771_ (.A(_16718_),
    .Y(_16724_));
 sky130_fd_sc_hd__a31oi_2 _43772_ (.A1(_16701_),
    .A2(_16706_),
    .A3(_16708_),
    .B1(_16724_),
    .Y(_16725_));
 sky130_fd_sc_hd__a21oi_1 _43773_ (.A1(_16725_),
    .A2(_16717_),
    .B1(_16720_),
    .Y(_16726_));
 sky130_fd_sc_hd__and3_1 _43774_ (.A(_16701_),
    .B(_16706_),
    .C(_16708_),
    .X(_16727_));
 sky130_fd_sc_hd__o21ai_2 _43775_ (.A1(_16709_),
    .A2(_16727_),
    .B1(_16724_),
    .Y(_16728_));
 sky130_fd_sc_hd__nand2_1 _43776_ (.A(_16726_),
    .B(_16728_),
    .Y(_16729_));
 sky130_fd_sc_hd__o21ai_2 _43777_ (.A1(_16455_),
    .A2(_16476_),
    .B1(_16454_),
    .Y(_16730_));
 sky130_fd_sc_hd__a21o_1 _43778_ (.A1(_16423_),
    .A2(_16425_),
    .B1(_16450_),
    .X(_16731_));
 sky130_fd_sc_hd__or2b_1 _43779_ (.A(_16340_),
    .B_N(_16365_),
    .X(_16732_));
 sky130_fd_sc_hd__xnor2_1 _43780_ (.A(_15771_),
    .B(_15776_),
    .Y(_16734_));
 sky130_fd_sc_hd__xor2_1 _43781_ (.A(_15769_),
    .B(_16734_),
    .X(_16735_));
 sky130_fd_sc_hd__a21oi_1 _43782_ (.A1(_16434_),
    .A2(_16438_),
    .B1(_16735_),
    .Y(_16736_));
 sky130_fd_sc_hd__and3_1 _43783_ (.A(_16434_),
    .B(_16438_),
    .C(_16735_),
    .X(_16737_));
 sky130_fd_sc_hd__or3_1 _43784_ (.A(_16736_),
    .B(_16737_),
    .C(_15803_),
    .X(_16738_));
 sky130_fd_sc_hd__o21ai_1 _43785_ (.A1(_16736_),
    .A2(_16737_),
    .B1(_16428_),
    .Y(_16739_));
 sky130_fd_sc_hd__nand2_1 _43786_ (.A(_16738_),
    .B(_16739_),
    .Y(_16740_));
 sky130_fd_sc_hd__a21oi_2 _43787_ (.A1(_16364_),
    .A2(_16732_),
    .B1(_16740_),
    .Y(_16741_));
 sky130_fd_sc_hd__o311a_1 _43788_ (.A1(net74),
    .A2(_16362_),
    .A3(_16363_),
    .B1(_16732_),
    .C1(_16740_),
    .X(_16742_));
 sky130_fd_sc_hd__o21a_1 _43789_ (.A1(_16439_),
    .A2(_16440_),
    .B1(_16443_),
    .X(_16743_));
 sky130_fd_sc_hd__o21ai_1 _43790_ (.A1(_16741_),
    .A2(_16742_),
    .B1(_16743_),
    .Y(_16745_));
 sky130_fd_sc_hd__or3_1 _43791_ (.A(_16743_),
    .B(_16741_),
    .C(_16742_),
    .X(_16746_));
 sky130_fd_sc_hd__nand2_1 _43792_ (.A(_16745_),
    .B(_16746_),
    .Y(_16747_));
 sky130_fd_sc_hd__o31a_1 _43793_ (.A1(_15664_),
    .A2(_12182_),
    .A3(_16391_),
    .B1(_15669_),
    .X(_16748_));
 sky130_fd_sc_hd__o31a_1 _43794_ (.A1(_15013_),
    .A2(_15014_),
    .A3(_15678_),
    .B1(_14439_),
    .X(_16749_));
 sky130_fd_sc_hd__nor2_1 _43795_ (.A(_16399_),
    .B(_16400_),
    .Y(_16750_));
 sky130_fd_sc_hd__o22ai_4 _43796_ (.A1(_16395_),
    .A2(_16748_),
    .B1(_16749_),
    .B2(_16750_),
    .Y(_16751_));
 sky130_fd_sc_hd__inv_2 _43797_ (.A(net76),
    .Y(_16752_));
 sky130_fd_sc_hd__nor2_1 _43798_ (.A(_16406_),
    .B(_16410_),
    .Y(_16753_));
 sky130_fd_sc_hd__nand2_1 _43799_ (.A(_16411_),
    .B(_16753_),
    .Y(_16754_));
 sky130_fd_sc_hd__or3_1 _43800_ (.A(_15664_),
    .B(_12182_),
    .C(_16391_),
    .X(_16756_));
 sky130_fd_sc_hd__a2111o_2 _43801_ (.A1(_15669_),
    .A2(_16756_),
    .B1(_16749_),
    .C1(_16750_),
    .D1(_16395_),
    .X(_16757_));
 sky130_fd_sc_hd__nand2_4 _43802_ (.A(_16754_),
    .B(_16757_),
    .Y(_16758_));
 sky130_fd_sc_hd__and2_1 _43803_ (.A(net76),
    .B(_16757_),
    .X(_16759_));
 sky130_fd_sc_hd__o22a_1 _43804_ (.A1(_16752_),
    .A2(_16758_),
    .B1(_16754_),
    .B2(_16759_),
    .X(_16760_));
 sky130_fd_sc_hd__clkbuf_2 _43805_ (.A(_14947_),
    .X(_16761_));
 sky130_fd_sc_hd__clkbuf_2 _43806_ (.A(_13552_),
    .X(_16762_));
 sky130_fd_sc_hd__nor2_2 _43807_ (.A(_16761_),
    .B(_16762_),
    .Y(_16763_));
 sky130_fd_sc_hd__and2_2 _43808_ (.A(_16761_),
    .B(_16762_),
    .X(_16764_));
 sky130_fd_sc_hd__o21a_1 _43809_ (.A1(_15648_),
    .A2(_09961_),
    .B1(_16370_),
    .X(_16765_));
 sky130_fd_sc_hd__a21oi_2 _43810_ (.A1(_15650_),
    .A2(_15651_),
    .B1(_16374_),
    .Y(_16767_));
 sky130_fd_sc_hd__o22ai_4 _43811_ (.A1(_16763_),
    .A2(_16764_),
    .B1(_16765_),
    .B2(_16767_),
    .Y(_16768_));
 sky130_fd_sc_hd__nor2_1 _43812_ (.A(_16763_),
    .B(_16764_),
    .Y(_16769_));
 sky130_fd_sc_hd__or3b_2 _43813_ (.A(_16767_),
    .B(_16765_),
    .C_N(_16769_),
    .X(_16770_));
 sky130_fd_sc_hd__o21ba_2 _43814_ (.A1(_16381_),
    .A2(_16377_),
    .B1_N(_16383_),
    .X(_16771_));
 sky130_fd_sc_hd__a21oi_4 _43815_ (.A1(_16768_),
    .A2(_16770_),
    .B1(_16771_),
    .Y(_16772_));
 sky130_fd_sc_hd__nand3_4 _43816_ (.A(_16771_),
    .B(_16768_),
    .C(_16770_),
    .Y(_16773_));
 sky130_fd_sc_hd__and2b_1 _43817_ (.A_N(_16772_),
    .B(_16773_),
    .X(_16774_));
 sky130_fd_sc_hd__xnor2_1 _43818_ (.A(_16760_),
    .B(_16774_),
    .Y(_16775_));
 sky130_fd_sc_hd__o21ba_4 _43819_ (.A1(_16387_),
    .A2(_16418_),
    .B1_N(_16775_),
    .X(_16776_));
 sky130_fd_sc_hd__nor3b_2 _43820_ (.A(_16387_),
    .B(_16418_),
    .C_N(_16775_),
    .Y(_16778_));
 sky130_fd_sc_hd__nor2_1 _43821_ (.A(_16776_),
    .B(net66),
    .Y(_16779_));
 sky130_fd_sc_hd__o21ai_1 _43822_ (.A1(_15725_),
    .A2(_16342_),
    .B1(_16361_),
    .Y(_16780_));
 sky130_fd_sc_hd__and2_1 _43823_ (.A(_16359_),
    .B(_16780_),
    .X(_16781_));
 sky130_fd_sc_hd__and3_4 _43824_ (.A(_16403_),
    .B(_16411_),
    .C(_16413_),
    .X(_16782_));
 sky130_fd_sc_hd__o2bb2a_1 _43825_ (.A1_N(_15730_),
    .A2_N(_15733_),
    .B1(_16346_),
    .B2(_11275_),
    .X(_16783_));
 sky130_fd_sc_hd__o21a_1 _43826_ (.A1(_16343_),
    .A2(_10077_),
    .B1(_16344_),
    .X(_16784_));
 sky130_fd_sc_hd__or3_1 _43827_ (.A(_15113_),
    .B(_15114_),
    .C(_15736_),
    .X(_16785_));
 sky130_fd_sc_hd__a21o_1 _43828_ (.A1(_14319_),
    .A2(_16785_),
    .B1(_16356_),
    .X(_16786_));
 sky130_fd_sc_hd__o21a_1 _43829_ (.A1(_16783_),
    .A2(_16784_),
    .B1(_16786_),
    .X(_16787_));
 sky130_fd_sc_hd__inv_2 _43830_ (.A(_16787_),
    .Y(_16789_));
 sky130_fd_sc_hd__a21o_1 _43831_ (.A1(_12421_),
    .A2(_15087_),
    .B1(_16343_),
    .X(_16790_));
 sky130_fd_sc_hd__a211o_1 _43832_ (.A1(_16344_),
    .A2(_16790_),
    .B1(_16783_),
    .C1(_16786_),
    .X(_16791_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _43833_ (.A(_15073_),
    .X(_16792_));
 sky130_fd_sc_hd__a21o_1 _43834_ (.A1(_16789_),
    .A2(_16791_),
    .B1(_16792_),
    .X(_16793_));
 sky130_fd_sc_hd__nand3_1 _43835_ (.A(_16789_),
    .B(_16791_),
    .C(_16792_),
    .Y(_16794_));
 sky130_fd_sc_hd__o211a_1 _43836_ (.A1(net77),
    .A2(_16782_),
    .B1(_16793_),
    .C1(_16794_),
    .X(_16795_));
 sky130_fd_sc_hd__a211oi_2 _43837_ (.A1(_16793_),
    .A2(_16794_),
    .B1(net77),
    .C1(_16782_),
    .Y(_16796_));
 sky130_fd_sc_hd__nor2_1 _43838_ (.A(_16795_),
    .B(_16796_),
    .Y(_16797_));
 sky130_fd_sc_hd__xnor2_1 _43839_ (.A(_16781_),
    .B(_16797_),
    .Y(_16798_));
 sky130_fd_sc_hd__nand2_1 _43840_ (.A(_16779_),
    .B(_16798_),
    .Y(_16800_));
 sky130_fd_sc_hd__or2_1 _43841_ (.A(_16798_),
    .B(_16779_),
    .X(_16801_));
 sky130_fd_sc_hd__inv_2 _43842_ (.A(_16422_),
    .Y(_16802_));
 sky130_fd_sc_hd__nand2_1 _43843_ (.A(_16419_),
    .B(_16802_),
    .Y(_16803_));
 sky130_fd_sc_hd__a21oi_1 _43844_ (.A1(_16800_),
    .A2(_16801_),
    .B1(_16803_),
    .Y(_16804_));
 sky130_fd_sc_hd__nand3_1 _43845_ (.A(_16803_),
    .B(_16800_),
    .C(_16801_),
    .Y(_16805_));
 sky130_fd_sc_hd__or2b_1 _43846_ (.A(_16804_),
    .B_N(_16805_),
    .X(_16806_));
 sky130_fd_sc_hd__xnor2_1 _43847_ (.A(_16747_),
    .B(_16806_),
    .Y(_16807_));
 sky130_fd_sc_hd__o211ai_2 _43848_ (.A1(_16423_),
    .A2(_16425_),
    .B1(_16731_),
    .C1(_16807_),
    .Y(_16808_));
 sky130_fd_sc_hd__a21o_1 _43849_ (.A1(_16424_),
    .A2(_16731_),
    .B1(_16807_),
    .X(_16809_));
 sky130_fd_sc_hd__o21ai_2 _43850_ (.A1(_15599_),
    .A2(_16464_),
    .B1(_16465_),
    .Y(_16811_));
 sky130_fd_sc_hd__or2_1 _43851_ (.A(_16430_),
    .B(_16446_),
    .X(_16812_));
 sky130_fd_sc_hd__a2111oi_1 _43852_ (.A1(_14839_),
    .A2(_15612_),
    .B1(_15611_),
    .C1(_14842_),
    .D1(_16456_),
    .Y(_16813_));
 sky130_fd_sc_hd__a31o_2 _43853_ (.A1(_14842_),
    .A2(_16457_),
    .A3(_16456_),
    .B1(_16813_),
    .X(_16814_));
 sky130_fd_sc_hd__xnor2_2 _43854_ (.A(_14860_),
    .B(_16814_),
    .Y(_16815_));
 sky130_fd_sc_hd__clkbuf_2 _43855_ (.A(_16815_),
    .X(_16816_));
 sky130_fd_sc_hd__a21oi_1 _43856_ (.A1(_16447_),
    .A2(_16812_),
    .B1(_16816_),
    .Y(_16817_));
 sky130_fd_sc_hd__o211ai_2 _43857_ (.A1(_16430_),
    .A2(_16446_),
    .B1(_16447_),
    .C1(_16816_),
    .Y(_16818_));
 sky130_fd_sc_hd__or2b_1 _43858_ (.A(_16817_),
    .B_N(_16818_),
    .X(_16819_));
 sky130_fd_sc_hd__xor2_1 _43859_ (.A(_16811_),
    .B(_16819_),
    .X(_16820_));
 sky130_fd_sc_hd__inv_2 _43860_ (.A(_16820_),
    .Y(_16822_));
 sky130_fd_sc_hd__nand3_1 _43861_ (.A(_16808_),
    .B(_16809_),
    .C(_16822_),
    .Y(_16823_));
 sky130_fd_sc_hd__a21o_1 _43862_ (.A1(_16808_),
    .A2(_16809_),
    .B1(_16822_),
    .X(_16824_));
 sky130_fd_sc_hd__nand2_1 _43863_ (.A(_16823_),
    .B(_16824_),
    .Y(_16825_));
 sky130_fd_sc_hd__xor2_1 _43864_ (.A(_16730_),
    .B(_16825_),
    .X(_16826_));
 sky130_fd_sc_hd__a21boi_1 _43865_ (.A1(_16723_),
    .A2(_16729_),
    .B1_N(_16826_),
    .Y(_16827_));
 sky130_fd_sc_hd__inv_2 _43866_ (.A(_16730_),
    .Y(_16828_));
 sky130_fd_sc_hd__a21oi_1 _43867_ (.A1(_16823_),
    .A2(_16824_),
    .B1(_16828_),
    .Y(_16829_));
 sky130_fd_sc_hd__and3_1 _43868_ (.A(_16828_),
    .B(_16823_),
    .C(_16824_),
    .X(_16830_));
 sky130_fd_sc_hd__o21bai_1 _43869_ (.A1(_16709_),
    .A2(_16714_),
    .B1_N(_16721_),
    .Y(_16831_));
 sky130_fd_sc_hd__o22ai_2 _43870_ (.A1(_16829_),
    .A2(_16830_),
    .B1(_16719_),
    .B2(_16831_),
    .Y(_16833_));
 sky130_fd_sc_hd__nand2_1 _43871_ (.A(_16725_),
    .B(_16717_),
    .Y(_16834_));
 sky130_fd_sc_hd__a21boi_2 _43872_ (.A1(_16834_),
    .A2(_16728_),
    .B1_N(_16721_),
    .Y(_16835_));
 sky130_fd_sc_hd__nor2_1 _43873_ (.A(_16833_),
    .B(_16835_),
    .Y(_16836_));
 sky130_fd_sc_hd__a31o_1 _43874_ (.A1(_16336_),
    .A2(_16482_),
    .A3(_16485_),
    .B1(_16479_),
    .X(_16837_));
 sky130_fd_sc_hd__o21bai_2 _43875_ (.A1(_16827_),
    .A2(_16836_),
    .B1_N(_16837_),
    .Y(_16838_));
 sky130_fd_sc_hd__a21bo_1 _43876_ (.A1(_16723_),
    .A2(_16729_),
    .B1_N(_16826_),
    .X(_16839_));
 sky130_fd_sc_hd__o211ai_1 _43877_ (.A1(_16833_),
    .A2(_16835_),
    .B1(_16837_),
    .C1(_16839_),
    .Y(_16840_));
 sky130_fd_sc_hd__clkbuf_2 _43878_ (.A(_16840_),
    .X(_16841_));
 sky130_fd_sc_hd__nand2_1 _43879_ (.A(_16838_),
    .B(_16841_),
    .Y(_16842_));
 sky130_fd_sc_hd__o21ai_1 _43880_ (.A1(_16036_),
    .A2(_16483_),
    .B1(_16334_),
    .Y(_16844_));
 sky130_fd_sc_hd__clkbuf_2 _43881_ (.A(_15577_),
    .X(_16845_));
 sky130_fd_sc_hd__nor2_1 _43882_ (.A(_16500_),
    .B(_16845_),
    .Y(_16846_));
 sky130_fd_sc_hd__and2_1 _43883_ (.A(_16500_),
    .B(_15577_),
    .X(_16847_));
 sky130_fd_sc_hd__o211a_1 _43884_ (.A1(_16846_),
    .A2(_16847_),
    .B1(_10304_),
    .C1(_10324_),
    .X(_16848_));
 sky130_fd_sc_hd__nor2_1 _43885_ (.A(_16846_),
    .B(_16847_),
    .Y(_16849_));
 sky130_fd_sc_hd__o211a_1 _43886_ (.A1(_15499_),
    .A2(_16518_),
    .B1(_16849_),
    .C1(_15491_),
    .X(_16850_));
 sky130_fd_sc_hd__nor2_1 _43887_ (.A(_16848_),
    .B(_16850_),
    .Y(_16851_));
 sky130_fd_sc_hd__o2111ai_1 _43888_ (.A1(_16322_),
    .A2(_16324_),
    .B1(_16509_),
    .C1(_12155_),
    .D1(_16045_),
    .Y(_16852_));
 sky130_fd_sc_hd__a22o_1 _43889_ (.A1(_15574_),
    .A2(_16045_),
    .B1(_16332_),
    .B2(_12155_),
    .X(_16853_));
 sky130_fd_sc_hd__a2bb2o_1 _43890_ (.A1_N(_16321_),
    .A2_N(_03566_),
    .B1(_16045_),
    .B2(_16502_),
    .X(_16855_));
 sky130_fd_sc_hd__and4_1 _43891_ (.A(_16852_),
    .B(_16853_),
    .C(_16855_),
    .D(_16509_),
    .X(_16856_));
 sky130_fd_sc_hd__a22oi_1 _43892_ (.A1(_16852_),
    .A2(_16853_),
    .B1(_16855_),
    .B2(_16518_),
    .Y(_16857_));
 sky130_fd_sc_hd__nor2_1 _43893_ (.A(_16856_),
    .B(_16857_),
    .Y(_16858_));
 sky130_fd_sc_hd__xnor2_1 _43894_ (.A(_16851_),
    .B(_16858_),
    .Y(_16859_));
 sky130_fd_sc_hd__a21o_1 _43895_ (.A1(_16484_),
    .A2(_16844_),
    .B1(_16859_),
    .X(_16860_));
 sky130_fd_sc_hd__nand3_1 _43896_ (.A(_16484_),
    .B(_16844_),
    .C(_16859_),
    .Y(_16861_));
 sky130_fd_sc_hd__o21bai_2 _43897_ (.A1(_16511_),
    .A2(_16499_),
    .B1_N(_16510_),
    .Y(_16862_));
 sky130_fd_sc_hd__a21o_1 _43898_ (.A1(_16860_),
    .A2(_16861_),
    .B1(_16862_),
    .X(_16863_));
 sky130_fd_sc_hd__nand3_2 _43899_ (.A(_16862_),
    .B(_16860_),
    .C(_16861_),
    .Y(_16864_));
 sky130_fd_sc_hd__nand2_2 _43900_ (.A(_16863_),
    .B(_16864_),
    .Y(_16866_));
 sky130_fd_sc_hd__nand2_1 _43901_ (.A(_16842_),
    .B(_16866_),
    .Y(_16867_));
 sky130_fd_sc_hd__nand4_2 _43902_ (.A(_16838_),
    .B(_16841_),
    .C(_16863_),
    .D(_16864_),
    .Y(_16868_));
 sky130_fd_sc_hd__nand3_1 _43903_ (.A(_16569_),
    .B(_16867_),
    .C(_16868_),
    .Y(_16869_));
 sky130_fd_sc_hd__a21o_1 _43904_ (.A1(_16838_),
    .A2(_16840_),
    .B1(_16866_),
    .X(_16870_));
 sky130_fd_sc_hd__nand3_1 _43905_ (.A(_16838_),
    .B(_16841_),
    .C(_16866_),
    .Y(_16871_));
 sky130_fd_sc_hd__a21oi_1 _43906_ (.A1(_16491_),
    .A2(_16522_),
    .B1(_16527_),
    .Y(_16872_));
 sky130_fd_sc_hd__nand3_2 _43907_ (.A(_16870_),
    .B(_16871_),
    .C(_16872_),
    .Y(_16873_));
 sky130_fd_sc_hd__or2b_2 _43908_ (.A(_16145_),
    .B_N(_16148_),
    .X(_16874_));
 sky130_fd_sc_hd__nand2_2 _43909_ (.A(_08961_),
    .B(_16494_),
    .Y(_16875_));
 sky130_fd_sc_hd__a211o_1 _43910_ (.A1(_15577_),
    .A2(_16494_),
    .B1(_08961_),
    .C1(_08969_),
    .X(_16877_));
 sky130_fd_sc_hd__a32o_1 _43911_ (.A1(_16496_),
    .A2(_15501_),
    .A3(_16495_),
    .B1(_07548_),
    .B2(_15499_),
    .X(_16878_));
 sky130_fd_sc_hd__and3_1 _43912_ (.A(_16875_),
    .B(_16877_),
    .C(_16878_),
    .X(_16879_));
 sky130_fd_sc_hd__a221o_1 _43913_ (.A1(_15499_),
    .A2(_07548_),
    .B1(_16875_),
    .B2(_16877_),
    .C1(_16498_),
    .X(_16880_));
 sky130_fd_sc_hd__and2b_1 _43914_ (.A_N(_16879_),
    .B(_16880_),
    .X(_16881_));
 sky130_fd_sc_hd__xor2_2 _43915_ (.A(_16874_),
    .B(_16881_),
    .X(_16882_));
 sky130_fd_sc_hd__o21bai_2 _43916_ (.A1(_16153_),
    .A2(_16149_),
    .B1_N(_16150_),
    .Y(_16883_));
 sky130_fd_sc_hd__and2_2 _43917_ (.A(_16882_),
    .B(_16883_),
    .X(_16884_));
 sky130_fd_sc_hd__nor2_1 _43918_ (.A(_16882_),
    .B(_16883_),
    .Y(_16885_));
 sky130_fd_sc_hd__nor2_1 _43919_ (.A(_16884_),
    .B(_16885_),
    .Y(_16886_));
 sky130_fd_sc_hd__a21oi_1 _43920_ (.A1(_16069_),
    .A2(_16493_),
    .B1(_16513_),
    .Y(_16888_));
 sky130_fd_sc_hd__a211o_1 _43921_ (.A1(_16520_),
    .A2(_16516_),
    .B1(_16886_),
    .C1(_16888_),
    .X(_16889_));
 sky130_fd_sc_hd__o21ai_1 _43922_ (.A1(_16888_),
    .A2(_16517_),
    .B1(_16886_),
    .Y(_16890_));
 sky130_fd_sc_hd__nand2_2 _43923_ (.A(_16889_),
    .B(_16890_),
    .Y(_16891_));
 sky130_fd_sc_hd__xor2_4 _43924_ (.A(_16158_),
    .B(_16891_),
    .X(_16892_));
 sky130_fd_sc_hd__a21o_1 _43925_ (.A1(_16869_),
    .A2(_16873_),
    .B1(_16892_),
    .X(_16893_));
 sky130_fd_sc_hd__nand3_1 _43926_ (.A(_16869_),
    .B(_16873_),
    .C(_16892_),
    .Y(_16894_));
 sky130_fd_sc_hd__a21boi_1 _43927_ (.A1(_16165_),
    .A2(_16530_),
    .B1_N(_16533_),
    .Y(_16895_));
 sky130_fd_sc_hd__and3_1 _43928_ (.A(_16893_),
    .B(_16894_),
    .C(_16895_),
    .X(_16896_));
 sky130_fd_sc_hd__a21oi_2 _43929_ (.A1(_16893_),
    .A2(_16894_),
    .B1(_16895_),
    .Y(_16897_));
 sky130_fd_sc_hd__a211o_1 _43930_ (.A1(_16160_),
    .A2(_16567_),
    .B1(_16896_),
    .C1(_16897_),
    .X(_16899_));
 sky130_fd_sc_hd__o211ai_1 _43931_ (.A1(_16896_),
    .A2(_16897_),
    .B1(_16160_),
    .C1(_16567_),
    .Y(_16900_));
 sky130_fd_sc_hd__nand2_1 _43932_ (.A(_16899_),
    .B(_16900_),
    .Y(_16901_));
 sky130_fd_sc_hd__o211a_1 _43933_ (.A1(_16541_),
    .A2(_16566_),
    .B1(_16540_),
    .C1(_16901_),
    .X(_16902_));
 sky130_fd_sc_hd__o21a_1 _43934_ (.A1(_16541_),
    .A2(_16566_),
    .B1(_16540_),
    .X(_16903_));
 sky130_fd_sc_hd__nor2_1 _43935_ (.A(_16903_),
    .B(_16901_),
    .Y(_16904_));
 sky130_fd_sc_hd__nor2_1 _43936_ (.A(_16902_),
    .B(_16904_),
    .Y(_16905_));
 sky130_fd_sc_hd__xnor2_1 _43937_ (.A(_16565_),
    .B(_16905_),
    .Y(_00019_));
 sky130_fd_sc_hd__nand3_1 _43938_ (.A(_16893_),
    .B(_16894_),
    .C(_16895_),
    .Y(_16906_));
 sky130_fd_sc_hd__a31oi_4 _43939_ (.A1(_16160_),
    .A2(_16567_),
    .A3(_16906_),
    .B1(_16897_),
    .Y(_16907_));
 sky130_fd_sc_hd__inv_2 _43940_ (.A(_16890_),
    .Y(_16909_));
 sky130_fd_sc_hd__or2_1 _43941_ (.A(_16110_),
    .B(_16113_),
    .X(_16910_));
 sky130_fd_sc_hd__o311a_1 _43942_ (.A1(_16888_),
    .A2(_16517_),
    .A3(_16886_),
    .B1(_16156_),
    .C1(_16910_),
    .X(_16911_));
 sky130_fd_sc_hd__a32oi_4 _43943_ (.A1(_16569_),
    .A2(_16867_),
    .A3(_16868_),
    .B1(_16873_),
    .B2(_16892_),
    .Y(_16912_));
 sky130_fd_sc_hd__o21ai_1 _43944_ (.A1(_16721_),
    .A2(_16719_),
    .B1(_16834_),
    .Y(_16913_));
 sky130_fd_sc_hd__clkbuf_2 _43945_ (.A(_16845_),
    .X(_16914_));
 sky130_fd_sc_hd__clkbuf_2 _43946_ (.A(_05099_),
    .X(_16915_));
 sky130_fd_sc_hd__a22o_1 _43947_ (.A1(_16323_),
    .A2(_16044_),
    .B1(_16332_),
    .B2(_16043_),
    .X(_16916_));
 sky130_fd_sc_hd__nor2_1 _43948_ (.A(_15570_),
    .B(_16507_),
    .Y(_16917_));
 sky130_fd_sc_hd__and3_1 _43949_ (.A(_16915_),
    .B(_12882_),
    .C(_15570_),
    .X(_16918_));
 sky130_fd_sc_hd__a221o_1 _43950_ (.A1(_13293_),
    .A2(_16917_),
    .B1(_16916_),
    .B2(_15574_),
    .C1(_16918_),
    .X(_16920_));
 sky130_fd_sc_hd__nand2_1 _43951_ (.A(_16920_),
    .B(_16914_),
    .Y(_16921_));
 sky130_fd_sc_hd__a31o_1 _43952_ (.A1(_16518_),
    .A2(_16915_),
    .A3(_16916_),
    .B1(_16921_),
    .X(_16922_));
 sky130_fd_sc_hd__a32o_1 _43953_ (.A1(_16518_),
    .A2(_16915_),
    .A3(_16916_),
    .B1(_16920_),
    .B2(_16845_),
    .X(_16923_));
 sky130_fd_sc_hd__inv_2 _43954_ (.A(_16923_),
    .Y(_16924_));
 sky130_fd_sc_hd__a22o_1 _43955_ (.A1(_16914_),
    .A2(_16922_),
    .B1(_16924_),
    .B2(_16920_),
    .X(_16925_));
 sky130_fd_sc_hd__nand2_2 _43956_ (.A(_16913_),
    .B(_16925_),
    .Y(_16926_));
 sky130_fd_sc_hd__a21oi_1 _43957_ (.A1(_16725_),
    .A2(_16717_),
    .B1(_16925_),
    .Y(_16927_));
 sky130_fd_sc_hd__o21ai_1 _43958_ (.A1(_16721_),
    .A2(_16719_),
    .B1(_16927_),
    .Y(_16928_));
 sky130_fd_sc_hd__a21o_1 _43959_ (.A1(_16851_),
    .A2(_16858_),
    .B1(_16856_),
    .X(_16929_));
 sky130_fd_sc_hd__a21o_1 _43960_ (.A1(_16926_),
    .A2(_16928_),
    .B1(_16929_),
    .X(_16931_));
 sky130_fd_sc_hd__nand3_2 _43961_ (.A(_16929_),
    .B(_16926_),
    .C(_16928_),
    .Y(_16932_));
 sky130_fd_sc_hd__inv_2 _43962_ (.A(_16705_),
    .Y(_16933_));
 sky130_fd_sc_hd__clkbuf_2 _43963_ (.A(_16043_),
    .X(_16934_));
 sky130_fd_sc_hd__and3_1 _43964_ (.A(_16324_),
    .B(_16701_),
    .C(_16934_),
    .X(_16935_));
 sky130_fd_sc_hd__a21o_1 _43965_ (.A1(_16811_),
    .A2(_16818_),
    .B1(_16817_),
    .X(_16936_));
 sky130_fd_sc_hd__o21ba_4 _43966_ (.A1(_16573_),
    .A2(_16653_),
    .B1_N(_16655_),
    .X(_16937_));
 sky130_fd_sc_hd__o21bai_4 _43967_ (.A1(_16269_),
    .A2(_16586_),
    .B1_N(_16587_),
    .Y(_16938_));
 sky130_fd_sc_hd__o2bb2a_1 _43968_ (.A1_N(_16219_),
    .A2_N(_16253_),
    .B1(_16644_),
    .B2(_16646_),
    .X(_16939_));
 sky130_fd_sc_hd__nor2_1 _43969_ (.A(_16610_),
    .B(_16609_),
    .Y(_16940_));
 sky130_fd_sc_hd__inv_2 _43970_ (.A(_16940_),
    .Y(_16942_));
 sky130_fd_sc_hd__nor2_1 _43971_ (.A(_16580_),
    .B(_16581_),
    .Y(_16943_));
 sky130_fd_sc_hd__nor2_1 _43972_ (.A(_16604_),
    .B(_16603_),
    .Y(_16944_));
 sky130_fd_sc_hd__o32a_1 _43973_ (.A1(_15332_),
    .A2(_16221_),
    .A3(_15329_),
    .B1(_15927_),
    .B2(_16944_),
    .X(_16945_));
 sky130_fd_sc_hd__xnor2_2 _43974_ (.A(_16574_),
    .B(_16945_),
    .Y(_16946_));
 sky130_fd_sc_hd__xnor2_1 _43975_ (.A(_16943_),
    .B(_16946_),
    .Y(_16947_));
 sky130_fd_sc_hd__a21oi_1 _43976_ (.A1(_16942_),
    .A2(_16614_),
    .B1(_16947_),
    .Y(_16948_));
 sky130_fd_sc_hd__and3_1 _43977_ (.A(_16942_),
    .B(_16614_),
    .C(_16947_),
    .X(_16949_));
 sky130_fd_sc_hd__nor3_1 _43978_ (.A(_16585_),
    .B(_16948_),
    .C(_16949_),
    .Y(_16950_));
 sky130_fd_sc_hd__o32a_1 _43979_ (.A1(net124),
    .A2(_16582_),
    .A3(_16583_),
    .B1(_16948_),
    .B2(_16949_),
    .X(_16951_));
 sky130_fd_sc_hd__or2_1 _43980_ (.A(_16950_),
    .B(_16951_),
    .X(_16953_));
 sky130_fd_sc_hd__o21ai_2 _43981_ (.A1(_16626_),
    .A2(_16636_),
    .B1(_16619_),
    .Y(_16954_));
 sky130_fd_sc_hd__nand3_1 _43982_ (.A(_16618_),
    .B(_16188_),
    .C(_16619_),
    .Y(_16955_));
 sky130_fd_sc_hd__and3b_1 _43983_ (.A_N(_16593_),
    .B(_16199_),
    .C(_16616_),
    .X(_16956_));
 sky130_fd_sc_hd__a311oi_1 _43984_ (.A1(_16602_),
    .A2(_16222_),
    .A3(_16575_),
    .B1(_16956_),
    .C1(_16597_),
    .Y(_16957_));
 sky130_fd_sc_hd__o2111a_1 _43985_ (.A1(_16597_),
    .A2(_16956_),
    .B1(_16602_),
    .C1(_16575_),
    .D1(_16222_),
    .X(_16958_));
 sky130_fd_sc_hd__nor2_1 _43986_ (.A(_16957_),
    .B(_16958_),
    .Y(_16959_));
 sky130_fd_sc_hd__and3_1 _43987_ (.A(_16955_),
    .B(_16625_),
    .C(_16959_),
    .X(_16960_));
 sky130_fd_sc_hd__o2bb2a_1 _43988_ (.A1_N(_16955_),
    .A2_N(_16625_),
    .B1(_16957_),
    .B2(_16958_),
    .X(_16961_));
 sky130_fd_sc_hd__nor2_1 _43989_ (.A(_16960_),
    .B(_16961_),
    .Y(_16962_));
 sky130_fd_sc_hd__a21bo_1 _43990_ (.A1(_16605_),
    .A2(_16606_),
    .B1_N(_16599_),
    .X(_16964_));
 sky130_fd_sc_hd__xor2_2 _43991_ (.A(_16962_),
    .B(_16964_),
    .X(_16965_));
 sky130_fd_sc_hd__nand2_2 _43992_ (.A(_16954_),
    .B(_16965_),
    .Y(_16966_));
 sky130_fd_sc_hd__or2_1 _43993_ (.A(_16965_),
    .B(_16954_),
    .X(_16967_));
 sky130_fd_sc_hd__a221o_1 _43994_ (.A1(_16212_),
    .A2(_16194_),
    .B1(_16637_),
    .B2(_16638_),
    .C1(_16639_),
    .X(_16968_));
 sky130_fd_sc_hd__a221o_1 _43995_ (.A1(_16966_),
    .A2(_16967_),
    .B1(_16968_),
    .B2(_16615_),
    .C1(_16643_),
    .X(_16969_));
 sky130_fd_sc_hd__a21oi_1 _43996_ (.A1(_16968_),
    .A2(_16615_),
    .B1(_16643_),
    .Y(_16970_));
 sky130_fd_sc_hd__nand3b_1 _43997_ (.A_N(_16970_),
    .B(_16966_),
    .C(_16967_),
    .Y(_16971_));
 sky130_fd_sc_hd__nand2_1 _43998_ (.A(_16969_),
    .B(_16971_),
    .Y(_16972_));
 sky130_fd_sc_hd__xor2_1 _43999_ (.A(_16953_),
    .B(_16972_),
    .X(_16973_));
 sky130_fd_sc_hd__o21a_2 _44000_ (.A1(_16939_),
    .A2(_16651_),
    .B1(_16973_),
    .X(_16975_));
 sky130_fd_sc_hd__a311oi_1 _44001_ (.A1(_16588_),
    .A2(_16589_),
    .A3(_16649_),
    .B1(_16973_),
    .C1(_16939_),
    .Y(_16976_));
 sky130_fd_sc_hd__or3_1 _44002_ (.A(_16938_),
    .B(_16975_),
    .C(net63),
    .X(_16977_));
 sky130_fd_sc_hd__o21ai_1 _44003_ (.A1(_16975_),
    .A2(net63),
    .B1(_16938_),
    .Y(_16978_));
 sky130_fd_sc_hd__nand2_2 _44004_ (.A(_16977_),
    .B(_16978_),
    .Y(_16979_));
 sky130_fd_sc_hd__xor2_4 _44005_ (.A(_16937_),
    .B(_16979_),
    .X(_16980_));
 sky130_fd_sc_hd__o21ai_4 _44006_ (.A1(_16290_),
    .A2(_16289_),
    .B1(_16662_),
    .Y(_16981_));
 sky130_fd_sc_hd__and4_2 _44007_ (.A(_16291_),
    .B(_16572_),
    .C(_16660_),
    .D(_16662_),
    .X(_16982_));
 sky130_fd_sc_hd__a22oi_4 _44008_ (.A1(_16660_),
    .A2(_16981_),
    .B1(_16298_),
    .B2(_16982_),
    .Y(_16983_));
 sky130_fd_sc_hd__nand2_2 _44009_ (.A(_16980_),
    .B(_16983_),
    .Y(_16984_));
 sky130_fd_sc_hd__inv_2 _44010_ (.A(_16980_),
    .Y(_16986_));
 sky130_fd_sc_hd__inv_2 _44011_ (.A(_16981_),
    .Y(_16987_));
 sky130_fd_sc_hd__inv_2 _44012_ (.A(_16982_),
    .Y(_16988_));
 sky130_fd_sc_hd__o22ai_1 _44013_ (.A1(_16661_),
    .A2(_16987_),
    .B1(_16988_),
    .B2(_16675_),
    .Y(_16989_));
 sky130_fd_sc_hd__nand2_2 _44014_ (.A(_16986_),
    .B(_16989_),
    .Y(_16990_));
 sky130_fd_sc_hd__nand2_1 _44015_ (.A(_16984_),
    .B(_16990_),
    .Y(_16991_));
 sky130_fd_sc_hd__a21oi_4 _44016_ (.A1(_16991_),
    .A2(_16669_),
    .B1(_12876_),
    .Y(_16992_));
 sky130_fd_sc_hd__o211ai_4 _44017_ (.A1(_16671_),
    .A2(_16672_),
    .B1(_16984_),
    .C1(_16990_),
    .Y(_16993_));
 sky130_fd_sc_hd__a221oi_2 _44018_ (.A1(_16660_),
    .A2(_16981_),
    .B1(_16298_),
    .B2(_16982_),
    .C1(_16986_),
    .Y(_16994_));
 sky130_fd_sc_hd__a21o_1 _44019_ (.A1(_16572_),
    .A2(_16662_),
    .B1(_16661_),
    .X(_16995_));
 sky130_fd_sc_hd__nand2_1 _44020_ (.A(_16298_),
    .B(_16982_),
    .Y(_16997_));
 sky130_fd_sc_hd__a21oi_1 _44021_ (.A1(_16995_),
    .A2(_16997_),
    .B1(_16980_),
    .Y(_16998_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44022_ (.A(_16668_),
    .X(_16999_));
 sky130_fd_sc_hd__o21ai_2 _44023_ (.A1(_16994_),
    .A2(_16998_),
    .B1(_16999_),
    .Y(_17000_));
 sky130_fd_sc_hd__a21oi_1 _44024_ (.A1(_17000_),
    .A2(_16993_),
    .B1(_16501_),
    .Y(_17001_));
 sky130_fd_sc_hd__a221oi_2 _44025_ (.A1(_16692_),
    .A2(_16018_),
    .B1(_16992_),
    .B2(_16993_),
    .C1(_17001_),
    .Y(_17002_));
 sky130_fd_sc_hd__o21ai_1 _44026_ (.A1(_16999_),
    .A2(_16991_),
    .B1(_16992_),
    .Y(_17003_));
 sky130_fd_sc_hd__a21o_1 _44027_ (.A1(_17000_),
    .A2(_16993_),
    .B1(_16501_),
    .X(_17004_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44028_ (.A(_16032_),
    .X(_17005_));
 sky130_fd_sc_hd__a21oi_1 _44029_ (.A1(_17003_),
    .A2(_17004_),
    .B1(_17005_),
    .Y(_17006_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44030_ (.A(_16171_),
    .X(_17008_));
 sky130_fd_sc_hd__a31o_1 _44031_ (.A1(_17008_),
    .A2(_16676_),
    .A3(_16679_),
    .B1(_16670_),
    .X(_17009_));
 sky130_fd_sc_hd__o21bai_2 _44032_ (.A1(_17002_),
    .A2(_17006_),
    .B1_N(_17009_),
    .Y(_17010_));
 sky130_fd_sc_hd__clkbuf_2 _44033_ (.A(_16022_),
    .X(_17011_));
 sky130_fd_sc_hd__clkbuf_2 _44034_ (.A(_16023_),
    .X(_17012_));
 sky130_fd_sc_hd__inv_2 _44035_ (.A(_16993_),
    .Y(_17013_));
 sky130_fd_sc_hd__nand2_1 _44036_ (.A(_17000_),
    .B(_16501_),
    .Y(_17014_));
 sky130_fd_sc_hd__o221ai_1 _44037_ (.A1(_17011_),
    .A2(_17012_),
    .B1(_17013_),
    .B2(_17014_),
    .C1(_17004_),
    .Y(_17015_));
 sky130_fd_sc_hd__a21o_1 _44038_ (.A1(_17003_),
    .A2(_17004_),
    .B1(_17005_),
    .X(_17016_));
 sky130_fd_sc_hd__o211ai_1 _44039_ (.A1(_16690_),
    .A2(_16670_),
    .B1(_17015_),
    .C1(_17016_),
    .Y(_17017_));
 sky130_fd_sc_hd__a22o_2 _44040_ (.A1(_16685_),
    .A2(_16694_),
    .B1(_16697_),
    .B2(_16702_),
    .X(_17019_));
 sky130_fd_sc_hd__a21o_1 _44041_ (.A1(_17010_),
    .A2(_17017_),
    .B1(_17019_),
    .X(_17020_));
 sky130_fd_sc_hd__clkbuf_2 _44042_ (.A(_17002_),
    .X(_17021_));
 sky130_fd_sc_hd__clkbuf_2 _44043_ (.A(_16681_),
    .X(_17022_));
 sky130_fd_sc_hd__o21ai_1 _44044_ (.A1(_17014_),
    .A2(_17013_),
    .B1(_17004_),
    .Y(_17023_));
 sky130_fd_sc_hd__o2bb2ai_2 _44045_ (.A1_N(_17022_),
    .A2_N(_17023_),
    .B1(_16670_),
    .B2(_16690_),
    .Y(_17024_));
 sky130_fd_sc_hd__o211ai_2 _44046_ (.A1(_17021_),
    .A2(_17024_),
    .B1(_17010_),
    .C1(_17019_),
    .Y(_17025_));
 sky130_fd_sc_hd__nand3_2 _44047_ (.A(_16936_),
    .B(_17020_),
    .C(_17025_),
    .Y(_17026_));
 sky130_fd_sc_hd__a21oi_1 _44048_ (.A1(_17010_),
    .A2(_17017_),
    .B1(_17019_),
    .Y(_17027_));
 sky130_fd_sc_hd__o211a_1 _44049_ (.A1(_17024_),
    .A2(_17021_),
    .B1(_17019_),
    .C1(_17010_),
    .X(_17028_));
 sky130_fd_sc_hd__a21oi_2 _44050_ (.A1(_16811_),
    .A2(_16818_),
    .B1(_16817_),
    .Y(_17030_));
 sky130_fd_sc_hd__o21ai_2 _44051_ (.A1(_17027_),
    .A2(_17028_),
    .B1(_17030_),
    .Y(_17031_));
 sky130_fd_sc_hd__a2bb2oi_1 _44052_ (.A1_N(_16933_),
    .A2_N(_16935_),
    .B1(_17026_),
    .B2(_17031_),
    .Y(_17032_));
 sky130_fd_sc_hd__a21oi_4 _44053_ (.A1(_16708_),
    .A2(_16701_),
    .B1(_16933_),
    .Y(_17033_));
 sky130_fd_sc_hd__o311a_1 _44054_ (.A1(_17030_),
    .A2(_17027_),
    .A3(_17028_),
    .B1(_17033_),
    .C1(_17031_),
    .X(_17034_));
 sky130_fd_sc_hd__a21bo_1 _44055_ (.A1(_16808_),
    .A2(_16822_),
    .B1_N(_16809_),
    .X(_17035_));
 sky130_fd_sc_hd__nor2_1 _44056_ (.A(_16776_),
    .B(_16798_),
    .Y(_17036_));
 sky130_fd_sc_hd__or3_2 _44057_ (.A(_14386_),
    .B(_16763_),
    .C(_16764_),
    .X(_17037_));
 sky130_fd_sc_hd__o21ai_2 _44058_ (.A1(_16763_),
    .A2(_16764_),
    .B1(_14386_),
    .Y(_17038_));
 sky130_fd_sc_hd__o21a_1 _44059_ (.A1(_16767_),
    .A2(_16765_),
    .B1(_16769_),
    .X(_17039_));
 sky130_fd_sc_hd__a221oi_4 _44060_ (.A1(_16761_),
    .A2(_16762_),
    .B1(_17037_),
    .B2(_17038_),
    .C1(_17039_),
    .Y(_17041_));
 sky130_fd_sc_hd__or2_1 _44061_ (.A(_15678_),
    .B(_16391_),
    .X(_17042_));
 sky130_fd_sc_hd__nand2_4 _44062_ (.A(_15678_),
    .B(_16391_),
    .Y(_17043_));
 sky130_fd_sc_hd__nand3_4 _44063_ (.A(_17042_),
    .B(_17043_),
    .C(_14469_),
    .Y(_17044_));
 sky130_fd_sc_hd__a21o_2 _44064_ (.A1(_17042_),
    .A2(_17043_),
    .B1(_14469_),
    .X(_17045_));
 sky130_fd_sc_hd__nand2_1 _44065_ (.A(_17044_),
    .B(_17045_),
    .Y(_17046_));
 sky130_fd_sc_hd__o211a_4 _44066_ (.A1(_16764_),
    .A2(_17039_),
    .B1(_17037_),
    .C1(_17038_),
    .X(_17047_));
 sky130_fd_sc_hd__or3_2 _44067_ (.A(_17041_),
    .B(_17046_),
    .C(_17047_),
    .X(_17048_));
 sky130_fd_sc_hd__buf_4 _44068_ (.A(_17046_),
    .X(_17049_));
 sky130_fd_sc_hd__o21ai_2 _44069_ (.A1(_17041_),
    .A2(_17047_),
    .B1(_17049_),
    .Y(_17050_));
 sky130_fd_sc_hd__a221o_4 _44070_ (.A1(_16760_),
    .A2(_16773_),
    .B1(_17048_),
    .B2(_17050_),
    .C1(_16772_),
    .X(_17052_));
 sky130_fd_sc_hd__a21oi_1 _44071_ (.A1(_16760_),
    .A2(_16773_),
    .B1(_16772_),
    .Y(_17053_));
 sky130_fd_sc_hd__nand3b_4 _44072_ (.A_N(_17053_),
    .B(_17048_),
    .C(_17050_),
    .Y(_17054_));
 sky130_fd_sc_hd__nand2_1 _44073_ (.A(_10045_),
    .B(_14290_),
    .Y(_17055_));
 sky130_fd_sc_hd__nand2_1 _44074_ (.A(_15736_),
    .B(_16344_),
    .Y(_17056_));
 sky130_fd_sc_hd__nand3_1 _44075_ (.A(_17055_),
    .B(_17056_),
    .C(_16792_),
    .Y(_17057_));
 sky130_fd_sc_hd__a21o_1 _44076_ (.A1(_17055_),
    .A2(_17056_),
    .B1(_15073_),
    .X(_17058_));
 sky130_fd_sc_hd__nand2_1 _44077_ (.A(_17057_),
    .B(_17058_),
    .Y(_17059_));
 sky130_fd_sc_hd__a21oi_1 _44078_ (.A1(net76),
    .A2(_16758_),
    .B1(_17059_),
    .Y(_17060_));
 sky130_fd_sc_hd__and3_1 _44079_ (.A(net76),
    .B(_16758_),
    .C(_17059_),
    .X(_17061_));
 sky130_fd_sc_hd__a21oi_1 _44080_ (.A1(_16791_),
    .A2(_16792_),
    .B1(_16787_),
    .Y(_17063_));
 sky130_fd_sc_hd__o21bai_1 _44081_ (.A1(_17060_),
    .A2(_17061_),
    .B1_N(_17063_),
    .Y(_17064_));
 sky130_fd_sc_hd__a2111o_1 _44082_ (.A1(_16791_),
    .A2(_16792_),
    .B1(_16787_),
    .C1(_17060_),
    .D1(_17061_),
    .X(_17065_));
 sky130_fd_sc_hd__and2_1 _44083_ (.A(_17064_),
    .B(_17065_),
    .X(_17066_));
 sky130_fd_sc_hd__a21bo_1 _44084_ (.A1(_17052_),
    .A2(_17054_),
    .B1_N(_17066_),
    .X(_17067_));
 sky130_fd_sc_hd__nand3b_2 _44085_ (.A_N(_17066_),
    .B(_17052_),
    .C(_17054_),
    .Y(_17068_));
 sky130_fd_sc_hd__a2bb2oi_1 _44086_ (.A1_N(net66),
    .A2_N(_17036_),
    .B1(_17067_),
    .B2(_17068_),
    .Y(_17069_));
 sky130_fd_sc_hd__and4bb_1 _44087_ (.A_N(net66),
    .B_N(_17036_),
    .C(_17067_),
    .D(_17068_),
    .X(_17070_));
 sky130_fd_sc_hd__a21o_1 _44088_ (.A1(_16434_),
    .A2(_16438_),
    .B1(_16735_),
    .X(_17071_));
 sky130_fd_sc_hd__and3_1 _44089_ (.A(_15771_),
    .B(_14903_),
    .C(_15776_),
    .X(_17072_));
 sky130_fd_sc_hd__and3_1 _44090_ (.A(_07040_),
    .B(_06992_),
    .C(_14572_),
    .X(_17074_));
 sky130_fd_sc_hd__or2_1 _44091_ (.A(_17072_),
    .B(_17074_),
    .X(_17075_));
 sky130_fd_sc_hd__xnor2_2 _44092_ (.A(_15803_),
    .B(_17075_),
    .Y(_17076_));
 sky130_fd_sc_hd__o21ba_1 _44093_ (.A1(_16781_),
    .A2(_16796_),
    .B1_N(_16795_),
    .X(_17077_));
 sky130_fd_sc_hd__xnor2_1 _44094_ (.A(_17076_),
    .B(_17077_),
    .Y(_17078_));
 sky130_fd_sc_hd__o211ai_1 _44095_ (.A1(_16737_),
    .A2(_16428_),
    .B1(_17071_),
    .C1(_17078_),
    .Y(_17079_));
 sky130_fd_sc_hd__a21o_1 _44096_ (.A1(_17071_),
    .A2(_16738_),
    .B1(_17078_),
    .X(_17080_));
 sky130_fd_sc_hd__and2_1 _44097_ (.A(_17079_),
    .B(_17080_),
    .X(_17081_));
 sky130_fd_sc_hd__or2_1 _44098_ (.A(_17070_),
    .B(_17081_),
    .X(_17082_));
 sky130_fd_sc_hd__o21ai_1 _44099_ (.A1(_17069_),
    .A2(_17070_),
    .B1(_17081_),
    .Y(_17083_));
 sky130_fd_sc_hd__o21a_1 _44100_ (.A1(_17069_),
    .A2(_17082_),
    .B1(_17083_),
    .X(_17085_));
 sky130_fd_sc_hd__o211a_1 _44101_ (.A1(_16747_),
    .A2(_16804_),
    .B1(_16805_),
    .C1(_17085_),
    .X(_17086_));
 sky130_fd_sc_hd__o21a_1 _44102_ (.A1(_16747_),
    .A2(_16804_),
    .B1(_16805_),
    .X(_17087_));
 sky130_fd_sc_hd__or2_1 _44103_ (.A(_17087_),
    .B(_17085_),
    .X(_17088_));
 sky130_fd_sc_hd__or2b_1 _44104_ (.A(_17086_),
    .B_N(_17088_),
    .X(_17089_));
 sky130_fd_sc_hd__or3b_4 _44105_ (.A(_15615_),
    .B(_15614_),
    .C_N(_16456_),
    .X(_17090_));
 sky130_fd_sc_hd__o21a_1 _44106_ (.A1(_15599_),
    .A2(net70),
    .B1(_17090_),
    .X(_17091_));
 sky130_fd_sc_hd__clkbuf_2 _44107_ (.A(_17091_),
    .X(_17092_));
 sky130_fd_sc_hd__nor2_1 _44108_ (.A(_16743_),
    .B(_16742_),
    .Y(_17093_));
 sky130_fd_sc_hd__inv_2 _44109_ (.A(_16815_),
    .Y(_17094_));
 sky130_fd_sc_hd__clkbuf_2 _44110_ (.A(_17094_),
    .X(_17096_));
 sky130_fd_sc_hd__o21ai_4 _44111_ (.A1(_16741_),
    .A2(_17093_),
    .B1(_17096_),
    .Y(_17097_));
 sky130_fd_sc_hd__or3_1 _44112_ (.A(_16741_),
    .B(_17096_),
    .C(_17093_),
    .X(_17098_));
 sky130_fd_sc_hd__nand2_1 _44113_ (.A(_17097_),
    .B(_17098_),
    .Y(_17099_));
 sky130_fd_sc_hd__and2b_2 _44114_ (.A_N(_17091_),
    .B(_17098_),
    .X(_17100_));
 sky130_fd_sc_hd__a22oi_4 _44115_ (.A1(_17092_),
    .A2(_17099_),
    .B1(_17100_),
    .B2(_17097_),
    .Y(_17101_));
 sky130_fd_sc_hd__xnor2_2 _44116_ (.A(_17089_),
    .B(_17101_),
    .Y(_17102_));
 sky130_fd_sc_hd__xor2_1 _44117_ (.A(_17035_),
    .B(_17102_),
    .X(_17103_));
 sky130_fd_sc_hd__o21ai_1 _44118_ (.A1(_17032_),
    .A2(_17034_),
    .B1(_17103_),
    .Y(_17104_));
 sky130_fd_sc_hd__xnor2_1 _44119_ (.A(_17035_),
    .B(_17102_),
    .Y(_17105_));
 sky130_fd_sc_hd__a21o_1 _44120_ (.A1(_17026_),
    .A2(_17031_),
    .B1(_17033_),
    .X(_17107_));
 sky130_fd_sc_hd__nand3_1 _44121_ (.A(_17031_),
    .B(_17033_),
    .C(_17026_),
    .Y(_17108_));
 sky130_fd_sc_hd__nand3_1 _44122_ (.A(_17105_),
    .B(_17107_),
    .C(_17108_),
    .Y(_17109_));
 sky130_fd_sc_hd__nand2_1 _44123_ (.A(_17104_),
    .B(_17109_),
    .Y(_17110_));
 sky130_fd_sc_hd__and2_1 _44124_ (.A(_16823_),
    .B(_16824_),
    .X(_17111_));
 sky130_fd_sc_hd__a21oi_1 _44125_ (.A1(_16726_),
    .A2(_16728_),
    .B1(_16826_),
    .Y(_17112_));
 sky130_fd_sc_hd__a22oi_1 _44126_ (.A1(_16730_),
    .A2(_17111_),
    .B1(_17112_),
    .B2(_16723_),
    .Y(_17113_));
 sky130_fd_sc_hd__nand2_2 _44127_ (.A(_17110_),
    .B(_17113_),
    .Y(_17114_));
 sky130_fd_sc_hd__o22ai_2 _44128_ (.A1(_16828_),
    .A2(_16825_),
    .B1(_16833_),
    .B2(_16835_),
    .Y(_17115_));
 sky130_fd_sc_hd__nand3_2 _44129_ (.A(_17115_),
    .B(_17104_),
    .C(_17109_),
    .Y(_17116_));
 sky130_fd_sc_hd__a22oi_1 _44130_ (.A1(_16931_),
    .A2(_16932_),
    .B1(_17114_),
    .B2(_17116_),
    .Y(_17118_));
 sky130_fd_sc_hd__nand2_1 _44131_ (.A(_16931_),
    .B(_16932_),
    .Y(_17119_));
 sky130_fd_sc_hd__nand2_1 _44132_ (.A(_17114_),
    .B(_17116_),
    .Y(_17120_));
 sky130_fd_sc_hd__nor2_1 _44133_ (.A(_17119_),
    .B(_17120_),
    .Y(_17121_));
 sky130_fd_sc_hd__nand2_1 _44134_ (.A(_17112_),
    .B(_16723_),
    .Y(_17122_));
 sky130_fd_sc_hd__a21oi_1 _44135_ (.A1(_16839_),
    .A2(_17122_),
    .B1(_16837_),
    .Y(_17123_));
 sky130_fd_sc_hd__o21a_1 _44136_ (.A1(_16866_),
    .A2(_17123_),
    .B1(_16841_),
    .X(_17124_));
 sky130_fd_sc_hd__o21ai_2 _44137_ (.A1(_17118_),
    .A2(_17121_),
    .B1(_17124_),
    .Y(_17125_));
 sky130_fd_sc_hd__o21ai_2 _44138_ (.A1(_16866_),
    .A2(_17123_),
    .B1(_16841_),
    .Y(_17126_));
 sky130_fd_sc_hd__a22o_1 _44139_ (.A1(_16931_),
    .A2(_16932_),
    .B1(_17114_),
    .B2(_17116_),
    .X(_17127_));
 sky130_fd_sc_hd__nand4_2 _44140_ (.A(_16931_),
    .B(_16932_),
    .C(_17114_),
    .D(_17116_),
    .Y(_17129_));
 sky130_fd_sc_hd__nand3_1 _44141_ (.A(_17126_),
    .B(_17127_),
    .C(_17129_),
    .Y(_17130_));
 sky130_fd_sc_hd__o41a_1 _44142_ (.A1(_09012_),
    .A2(_07548_),
    .A3(_16846_),
    .A4(_16847_),
    .B1(_16875_),
    .X(_17131_));
 sky130_fd_sc_hd__nor4b_1 _44143_ (.A(_09012_),
    .B(_16875_),
    .C(_07548_),
    .D_N(_16849_),
    .Y(_17132_));
 sky130_fd_sc_hd__or2_2 _44144_ (.A(_17131_),
    .B(_17132_),
    .X(_17133_));
 sky130_fd_sc_hd__a21oi_4 _44145_ (.A1(_16874_),
    .A2(_16880_),
    .B1(_16879_),
    .Y(_17134_));
 sky130_fd_sc_hd__xnor2_1 _44146_ (.A(_17133_),
    .B(_17134_),
    .Y(_17135_));
 sky130_fd_sc_hd__a21o_1 _44147_ (.A1(_16860_),
    .A2(_16864_),
    .B1(_17135_),
    .X(_17136_));
 sky130_fd_sc_hd__nand3_1 _44148_ (.A(_16860_),
    .B(_16864_),
    .C(_17135_),
    .Y(_17137_));
 sky130_fd_sc_hd__buf_1 _44149_ (.A(_17137_),
    .X(_17138_));
 sky130_fd_sc_hd__a21oi_1 _44150_ (.A1(_17136_),
    .A2(_17138_),
    .B1(_16884_),
    .Y(_17140_));
 sky130_fd_sc_hd__inv_2 _44151_ (.A(_16884_),
    .Y(_17141_));
 sky130_fd_sc_hd__a21oi_2 _44152_ (.A1(_16860_),
    .A2(_16864_),
    .B1(_17135_),
    .Y(_17142_));
 sky130_fd_sc_hd__nor3b_1 _44153_ (.A(_17141_),
    .B(_17142_),
    .C_N(_17137_),
    .Y(_17143_));
 sky130_fd_sc_hd__nor2_1 _44154_ (.A(_17140_),
    .B(_17143_),
    .Y(_17144_));
 sky130_fd_sc_hd__a21oi_2 _44155_ (.A1(_17125_),
    .A2(_17130_),
    .B1(_17144_),
    .Y(_17145_));
 sky130_fd_sc_hd__and3_1 _44156_ (.A(_17141_),
    .B(_17136_),
    .C(_17138_),
    .X(_17146_));
 sky130_fd_sc_hd__a21oi_1 _44157_ (.A1(_17136_),
    .A2(_17138_),
    .B1(_17141_),
    .Y(_17147_));
 sky130_fd_sc_hd__o211a_1 _44158_ (.A1(_17146_),
    .A2(_17147_),
    .B1(_17125_),
    .C1(_17130_),
    .X(_17148_));
 sky130_fd_sc_hd__nor3_1 _44159_ (.A(_16912_),
    .B(_17145_),
    .C(_17148_),
    .Y(_17149_));
 sky130_fd_sc_hd__o21a_1 _44160_ (.A1(_17145_),
    .A2(_17148_),
    .B1(_16912_),
    .X(_17151_));
 sky130_fd_sc_hd__o22ai_1 _44161_ (.A1(_16909_),
    .A2(_16911_),
    .B1(_17149_),
    .B2(_17151_),
    .Y(_17152_));
 sky130_fd_sc_hd__nand2_1 _44162_ (.A(_16873_),
    .B(_16892_),
    .Y(_17153_));
 sky130_fd_sc_hd__a211o_1 _44163_ (.A1(_16869_),
    .A2(_17153_),
    .B1(_17145_),
    .C1(_17148_),
    .X(_17154_));
 sky130_fd_sc_hd__o21ai_1 _44164_ (.A1(_17145_),
    .A2(_17148_),
    .B1(_16912_),
    .Y(_17155_));
 sky130_fd_sc_hd__nor2_1 _44165_ (.A(_16909_),
    .B(_16911_),
    .Y(_17156_));
 sky130_fd_sc_hd__nand3_1 _44166_ (.A(_17154_),
    .B(_17155_),
    .C(_17156_),
    .Y(_17157_));
 sky130_fd_sc_hd__nand2_1 _44167_ (.A(_17152_),
    .B(_17157_),
    .Y(_17158_));
 sky130_fd_sc_hd__xor2_2 _44168_ (.A(_16907_),
    .B(_17158_),
    .X(_17159_));
 sky130_fd_sc_hd__o21bai_1 _44169_ (.A1(_16903_),
    .A2(_16901_),
    .B1_N(_16546_),
    .Y(_17160_));
 sky130_fd_sc_hd__o2bb2a_1 _44170_ (.A1_N(_16903_),
    .A2_N(_16901_),
    .B1(_17160_),
    .B2(_16563_),
    .X(_17162_));
 sky130_fd_sc_hd__xor2_1 _44171_ (.A(_17159_),
    .B(_17162_),
    .X(_00020_));
 sky130_fd_sc_hd__and3_1 _44172_ (.A(_17115_),
    .B(_17104_),
    .C(_17109_),
    .X(_17163_));
 sky130_fd_sc_hd__a31o_1 _44173_ (.A1(_16931_),
    .A2(_16932_),
    .A3(_17114_),
    .B1(_17163_),
    .X(_17164_));
 sky130_fd_sc_hd__and2_1 _44174_ (.A(_17035_),
    .B(_17102_),
    .X(_17165_));
 sky130_fd_sc_hd__o22ai_1 _44175_ (.A1(_17035_),
    .A2(_17102_),
    .B1(_17032_),
    .B2(_17034_),
    .Y(_17166_));
 sky130_fd_sc_hd__nand2b_1 _44176_ (.A_N(_17165_),
    .B(_17166_),
    .Y(_17167_));
 sky130_fd_sc_hd__inv_2 _44177_ (.A(_17097_),
    .Y(_17168_));
 sky130_fd_sc_hd__inv_2 _44178_ (.A(_17024_),
    .Y(_17169_));
 sky130_fd_sc_hd__inv_2 _44179_ (.A(_16979_),
    .Y(_17170_));
 sky130_fd_sc_hd__o22ai_2 _44180_ (.A1(_16937_),
    .A2(_17170_),
    .B1(_16980_),
    .B2(_16983_),
    .Y(_17172_));
 sky130_fd_sc_hd__buf_6 _44181_ (.A(_17172_),
    .X(_17173_));
 sky130_fd_sc_hd__inv_2 _44182_ (.A(net63),
    .Y(_17174_));
 sky130_fd_sc_hd__nor2_2 _44183_ (.A(_16948_),
    .B(_16950_),
    .Y(_17175_));
 sky130_fd_sc_hd__a21o_1 _44184_ (.A1(_16964_),
    .A2(_16962_),
    .B1(_16961_),
    .X(_17176_));
 sky130_fd_sc_hd__o221a_1 _44185_ (.A1(_16257_),
    .A2(_15370_),
    .B1(_15304_),
    .B2(_15299_),
    .C1(_16945_),
    .X(_17177_));
 sky130_fd_sc_hd__or3b_2 _44186_ (.A(_16221_),
    .B(_15299_),
    .C_N(_16575_),
    .X(_17178_));
 sky130_fd_sc_hd__o32a_1 _44187_ (.A1(_15332_),
    .A2(_15329_),
    .A3(_17178_),
    .B1(_16946_),
    .B2(_16943_),
    .X(_17179_));
 sky130_fd_sc_hd__nor2_1 _44188_ (.A(_17177_),
    .B(_17179_),
    .Y(_17180_));
 sky130_fd_sc_hd__xor2_1 _44189_ (.A(_17176_),
    .B(_17180_),
    .X(_17181_));
 sky130_fd_sc_hd__a32oi_2 _44190_ (.A1(_16619_),
    .A2(_16632_),
    .A3(_16633_),
    .B1(_16954_),
    .B2(_16965_),
    .Y(_17183_));
 sky130_fd_sc_hd__a211o_1 _44191_ (.A1(_16616_),
    .A2(_16593_),
    .B1(_16201_),
    .C1(_16197_),
    .X(_17184_));
 sky130_fd_sc_hd__and3_1 _44192_ (.A(_16222_),
    .B(_16575_),
    .C(_16602_),
    .X(_17185_));
 sky130_fd_sc_hd__or3b_1 _44193_ (.A(_16596_),
    .B(_17185_),
    .C_N(_16234_),
    .X(_17186_));
 sky130_fd_sc_hd__or4b_1 _44194_ (.A(_16593_),
    .B(_07702_),
    .C(_17178_),
    .D_N(_16616_),
    .X(_17187_));
 sky130_fd_sc_hd__and3_1 _44195_ (.A(_17184_),
    .B(_17186_),
    .C(_17187_),
    .X(_17188_));
 sky130_fd_sc_hd__a22oi_1 _44196_ (.A1(_15843_),
    .A2(_16594_),
    .B1(_16635_),
    .B2(_17184_),
    .Y(_17189_));
 sky130_fd_sc_hd__xnor2_1 _44197_ (.A(_17188_),
    .B(_17189_),
    .Y(_17190_));
 sky130_fd_sc_hd__xnor2_1 _44198_ (.A(_17183_),
    .B(_17190_),
    .Y(_17191_));
 sky130_fd_sc_hd__xor2_2 _44199_ (.A(_17181_),
    .B(_17191_),
    .X(_17192_));
 sky130_fd_sc_hd__o21ai_2 _44200_ (.A1(_16953_),
    .A2(_16972_),
    .B1(_16971_),
    .Y(_17194_));
 sky130_fd_sc_hd__xor2_2 _44201_ (.A(_17192_),
    .B(_17194_),
    .X(_17195_));
 sky130_fd_sc_hd__xor2_4 _44202_ (.A(_17175_),
    .B(_17195_),
    .X(_17196_));
 sky130_fd_sc_hd__a211o_1 _44203_ (.A1(_16938_),
    .A2(_17174_),
    .B1(_17196_),
    .C1(_16975_),
    .X(_17197_));
 sky130_fd_sc_hd__a21oi_2 _44204_ (.A1(_16938_),
    .A2(_17174_),
    .B1(_16975_),
    .Y(_17198_));
 sky130_fd_sc_hd__inv_2 _44205_ (.A(_17196_),
    .Y(_17199_));
 sky130_fd_sc_hd__or2_2 _44206_ (.A(_17198_),
    .B(_17199_),
    .X(_17200_));
 sky130_fd_sc_hd__nand2_1 _44207_ (.A(_17197_),
    .B(_17200_),
    .Y(_17201_));
 sky130_fd_sc_hd__nand2_1 _44208_ (.A(_17173_),
    .B(_17201_),
    .Y(_17202_));
 sky130_fd_sc_hd__and2_1 _44209_ (.A(_17197_),
    .B(_17200_),
    .X(_17203_));
 sky130_fd_sc_hd__o221ai_4 _44210_ (.A1(_16937_),
    .A2(_17170_),
    .B1(_16980_),
    .B2(_16983_),
    .C1(_17203_),
    .Y(_17205_));
 sky130_fd_sc_hd__and3_1 _44211_ (.A(_17202_),
    .B(_17205_),
    .C(_16669_),
    .X(_17206_));
 sky130_fd_sc_hd__a21oi_1 _44212_ (.A1(_17202_),
    .A2(_17205_),
    .B1(_16999_),
    .Y(_17207_));
 sky130_fd_sc_hd__o21ai_2 _44213_ (.A1(_17206_),
    .A2(_17207_),
    .B1(_16058_),
    .Y(_17208_));
 sky130_fd_sc_hd__nand3_1 _44214_ (.A(_17202_),
    .B(_17205_),
    .C(_16999_),
    .Y(_17209_));
 sky130_fd_sc_hd__nand3b_1 _44215_ (.A_N(_17207_),
    .B(_16501_),
    .C(_17209_),
    .Y(_17210_));
 sky130_fd_sc_hd__a21o_1 _44216_ (.A1(_17208_),
    .A2(_17210_),
    .B1(_17005_),
    .X(_17211_));
 sky130_fd_sc_hd__clkbuf_2 _44217_ (.A(_17207_),
    .X(_17212_));
 sky130_fd_sc_hd__a31o_1 _44218_ (.A1(_17202_),
    .A2(_17205_),
    .A3(_16999_),
    .B1(_16058_),
    .X(_17213_));
 sky130_fd_sc_hd__o221ai_4 _44219_ (.A1(_17011_),
    .A2(_17012_),
    .B1(_17212_),
    .B2(_17213_),
    .C1(_17208_),
    .Y(_17214_));
 sky130_fd_sc_hd__o211ai_4 _44220_ (.A1(_16992_),
    .A2(_17013_),
    .B1(_17211_),
    .C1(_17214_),
    .Y(_17216_));
 sky130_fd_sc_hd__a21oi_1 _44221_ (.A1(_17208_),
    .A2(_17210_),
    .B1(_17005_),
    .Y(_17217_));
 sky130_fd_sc_hd__o221a_1 _44222_ (.A1(_17011_),
    .A2(_17012_),
    .B1(_17212_),
    .B2(_17213_),
    .C1(_17208_),
    .X(_17218_));
 sky130_fd_sc_hd__a31o_1 _44223_ (.A1(_16171_),
    .A2(_16984_),
    .A3(_16990_),
    .B1(_16992_),
    .X(_17219_));
 sky130_fd_sc_hd__inv_2 _44224_ (.A(_17219_),
    .Y(_17220_));
 sky130_fd_sc_hd__o21ai_2 _44225_ (.A1(_17217_),
    .A2(_17218_),
    .B1(_17220_),
    .Y(_17221_));
 sky130_fd_sc_hd__o211ai_4 _44226_ (.A1(_17021_),
    .A2(_17169_),
    .B1(_17216_),
    .C1(_17221_),
    .Y(_17222_));
 sky130_fd_sc_hd__o21ai_1 _44227_ (.A1(_17022_),
    .A2(_17023_),
    .B1(_17024_),
    .Y(_17223_));
 sky130_fd_sc_hd__a21o_1 _44228_ (.A1(_17216_),
    .A2(_17221_),
    .B1(_17223_),
    .X(_17224_));
 sky130_fd_sc_hd__o211ai_4 _44229_ (.A1(_17168_),
    .A2(_17100_),
    .B1(_17222_),
    .C1(_17224_),
    .Y(_17225_));
 sky130_fd_sc_hd__o211a_1 _44230_ (.A1(_17021_),
    .A2(_17169_),
    .B1(_17216_),
    .C1(_17221_),
    .X(_17227_));
 sky130_fd_sc_hd__a21oi_1 _44231_ (.A1(_17216_),
    .A2(_17221_),
    .B1(_17223_),
    .Y(_17228_));
 sky130_fd_sc_hd__nor2_1 _44232_ (.A(_17168_),
    .B(_17100_),
    .Y(_17229_));
 sky130_fd_sc_hd__o21ai_2 _44233_ (.A1(_17227_),
    .A2(_17228_),
    .B1(_17229_),
    .Y(_17230_));
 sky130_fd_sc_hd__inv_2 _44234_ (.A(_17019_),
    .Y(_17231_));
 sky130_fd_sc_hd__o21ai_1 _44235_ (.A1(_17021_),
    .A2(_17024_),
    .B1(_17010_),
    .Y(_17232_));
 sky130_fd_sc_hd__o2bb2ai_2 _44236_ (.A1_N(_17225_),
    .A2_N(_17230_),
    .B1(_17231_),
    .B2(_17232_),
    .Y(_17233_));
 sky130_fd_sc_hd__buf_1 _44237_ (.A(_17076_),
    .X(_17234_));
 sky130_fd_sc_hd__or2_1 _44238_ (.A(_17234_),
    .B(_17077_),
    .X(_17235_));
 sky130_fd_sc_hd__a21oi_2 _44239_ (.A1(_17235_),
    .A2(_17080_),
    .B1(_16816_),
    .Y(_17236_));
 sky130_fd_sc_hd__a31o_1 _44240_ (.A1(_16816_),
    .A2(_17235_),
    .A3(_17080_),
    .B1(_17092_),
    .X(_17238_));
 sky130_fd_sc_hd__and2_1 _44241_ (.A(_16816_),
    .B(_17080_),
    .X(_17239_));
 sky130_fd_sc_hd__a21o_1 _44242_ (.A1(_17239_),
    .A2(_17235_),
    .B1(_17236_),
    .X(_17240_));
 sky130_fd_sc_hd__a2bb2o_1 _44243_ (.A1_N(_17236_),
    .A2_N(_17238_),
    .B1(_17092_),
    .B2(_17240_),
    .X(_17241_));
 sky130_fd_sc_hd__o21ba_1 _44244_ (.A1(_17063_),
    .A2(_17061_),
    .B1_N(_17060_),
    .X(_17242_));
 sky130_fd_sc_hd__nor2_1 _44245_ (.A(_17242_),
    .B(_17234_),
    .Y(_17243_));
 sky130_fd_sc_hd__and2_1 _44246_ (.A(_17234_),
    .B(_17242_),
    .X(_17244_));
 sky130_fd_sc_hd__o21bai_2 _44247_ (.A1(_17074_),
    .A2(_16428_),
    .B1_N(_17072_),
    .Y(_17245_));
 sky130_fd_sc_hd__o21ba_1 _44248_ (.A1(_17243_),
    .A2(_17244_),
    .B1_N(_17245_),
    .X(_17246_));
 sky130_fd_sc_hd__a21boi_1 _44249_ (.A1(_17234_),
    .A2(_17242_),
    .B1_N(_17245_),
    .Y(_17247_));
 sky130_fd_sc_hd__o21a_1 _44250_ (.A1(_17234_),
    .A2(_17242_),
    .B1(_17247_),
    .X(_17249_));
 sky130_fd_sc_hd__o21ai_2 _44251_ (.A1(_10045_),
    .A2(_14290_),
    .B1(_17057_),
    .Y(_17250_));
 sky130_fd_sc_hd__and3_1 _44252_ (.A(_17059_),
    .B(_17043_),
    .C(_17044_),
    .X(_17251_));
 sky130_fd_sc_hd__a21oi_1 _44253_ (.A1(_17043_),
    .A2(_17044_),
    .B1(_17059_),
    .Y(_17252_));
 sky130_fd_sc_hd__nor2_1 _44254_ (.A(_17251_),
    .B(_17252_),
    .Y(_17253_));
 sky130_fd_sc_hd__xnor2_1 _44255_ (.A(_17250_),
    .B(_17253_),
    .Y(_17254_));
 sky130_fd_sc_hd__nor2_1 _44256_ (.A(_17046_),
    .B(_17041_),
    .Y(_17255_));
 sky130_fd_sc_hd__nor3_1 _44257_ (.A(_16761_),
    .B(_16762_),
    .C(_16370_),
    .Y(_17256_));
 sky130_fd_sc_hd__and3_4 _44258_ (.A(_16761_),
    .B(_16762_),
    .C(_16370_),
    .X(_17257_));
 sky130_fd_sc_hd__or3_1 _44259_ (.A(net215),
    .B(_17257_),
    .C(_17046_),
    .X(_17258_));
 sky130_fd_sc_hd__o21ai_1 _44260_ (.A1(net215),
    .A2(_17257_),
    .B1(_17046_),
    .Y(_17260_));
 sky130_fd_sc_hd__o211a_4 _44261_ (.A1(_17255_),
    .A2(_17047_),
    .B1(_17258_),
    .C1(_17260_),
    .X(_17261_));
 sky130_fd_sc_hd__a211o_4 _44262_ (.A1(_17258_),
    .A2(_17260_),
    .B1(_17255_),
    .C1(_17047_),
    .X(_17262_));
 sky130_fd_sc_hd__and2b_1 _44263_ (.A_N(_17261_),
    .B(_17262_),
    .X(_17263_));
 sky130_fd_sc_hd__xor2_1 _44264_ (.A(_17254_),
    .B(_17263_),
    .X(_17264_));
 sky130_fd_sc_hd__nand3_1 _44265_ (.A(_17264_),
    .B(_17068_),
    .C(_17054_),
    .Y(_17265_));
 sky130_fd_sc_hd__a21o_1 _44266_ (.A1(_17054_),
    .A2(_17068_),
    .B1(_17264_),
    .X(_17266_));
 sky130_fd_sc_hd__nand2_1 _44267_ (.A(_17265_),
    .B(_17266_),
    .Y(_17267_));
 sky130_fd_sc_hd__o21a_1 _44268_ (.A1(_17246_),
    .A2(_17249_),
    .B1(_17267_),
    .X(_17268_));
 sky130_fd_sc_hd__and2b_1 _44269_ (.A_N(_17069_),
    .B(_17081_),
    .X(_17269_));
 sky130_fd_sc_hd__or2_1 _44270_ (.A(_17070_),
    .B(_17269_),
    .X(_17271_));
 sky130_fd_sc_hd__or3_2 _44271_ (.A(_17246_),
    .B(_17249_),
    .C(_17267_),
    .X(_17272_));
 sky130_fd_sc_hd__nand2_1 _44272_ (.A(_17271_),
    .B(_17272_),
    .Y(_17273_));
 sky130_fd_sc_hd__inv_2 _44273_ (.A(_17268_),
    .Y(_17274_));
 sky130_fd_sc_hd__a21oi_1 _44274_ (.A1(_17272_),
    .A2(_17274_),
    .B1(_17271_),
    .Y(_17275_));
 sky130_fd_sc_hd__o21ba_1 _44275_ (.A1(_17268_),
    .A2(_17273_),
    .B1_N(_17275_),
    .X(_17276_));
 sky130_fd_sc_hd__xnor2_1 _44276_ (.A(_17241_),
    .B(_17276_),
    .Y(_17277_));
 sky130_fd_sc_hd__inv_2 _44277_ (.A(_17101_),
    .Y(_17278_));
 sky130_fd_sc_hd__a21oi_1 _44278_ (.A1(_17088_),
    .A2(_17278_),
    .B1(_17086_),
    .Y(_17279_));
 sky130_fd_sc_hd__nand2_1 _44279_ (.A(_17277_),
    .B(_17279_),
    .Y(_17280_));
 sky130_fd_sc_hd__or2_1 _44280_ (.A(_17279_),
    .B(_17277_),
    .X(_17282_));
 sky130_fd_sc_hd__and2_1 _44281_ (.A(_17280_),
    .B(_17282_),
    .X(_17283_));
 sky130_fd_sc_hd__nand3_2 _44282_ (.A(_17230_),
    .B(_17028_),
    .C(_17225_),
    .Y(_17284_));
 sky130_fd_sc_hd__nand3_2 _44283_ (.A(_17233_),
    .B(_17283_),
    .C(_17284_),
    .Y(_17285_));
 sky130_fd_sc_hd__a21o_1 _44284_ (.A1(_17284_),
    .A2(_17233_),
    .B1(_17283_),
    .X(_17286_));
 sky130_fd_sc_hd__nand3_1 _44285_ (.A(_17167_),
    .B(_17285_),
    .C(_17286_),
    .Y(_17287_));
 sky130_fd_sc_hd__and3_1 _44286_ (.A(_17233_),
    .B(_17283_),
    .C(_17284_),
    .X(_17288_));
 sky130_fd_sc_hd__a21oi_1 _44287_ (.A1(_17284_),
    .A2(_17233_),
    .B1(_17283_),
    .Y(_17289_));
 sky130_fd_sc_hd__o21bai_2 _44288_ (.A1(_17288_),
    .A2(_17289_),
    .B1_N(_17167_),
    .Y(_17290_));
 sky130_fd_sc_hd__a21oi_2 _44289_ (.A1(_17020_),
    .A2(_17025_),
    .B1(_16936_),
    .Y(_17291_));
 sky130_fd_sc_hd__o21ai_1 _44290_ (.A1(_17033_),
    .A2(_17291_),
    .B1(_17026_),
    .Y(_17293_));
 sky130_fd_sc_hd__o21ai_2 _44291_ (.A1(_15574_),
    .A2(_16507_),
    .B1(_12882_),
    .Y(_17294_));
 sky130_fd_sc_hd__and3_1 _44292_ (.A(_16507_),
    .B(_16915_),
    .C(_16500_),
    .X(_17295_));
 sky130_fd_sc_hd__o21a_2 _44293_ (.A1(_17294_),
    .A2(_17295_),
    .B1(_16845_),
    .X(_17296_));
 sky130_fd_sc_hd__a311oi_4 _44294_ (.A1(_16707_),
    .A2(_16509_),
    .A3(_16915_),
    .B1(_16845_),
    .C1(_17294_),
    .Y(_17297_));
 sky130_fd_sc_hd__or2_1 _44295_ (.A(_17296_),
    .B(_17297_),
    .X(_17298_));
 sky130_fd_sc_hd__inv_2 _44296_ (.A(_17298_),
    .Y(_17299_));
 sky130_fd_sc_hd__nand2_2 _44297_ (.A(_17293_),
    .B(_17299_),
    .Y(_17300_));
 sky130_fd_sc_hd__o221ai_4 _44298_ (.A1(_17033_),
    .A2(_17291_),
    .B1(_17296_),
    .B2(_17297_),
    .C1(_17026_),
    .Y(_17301_));
 sky130_fd_sc_hd__a21oi_1 _44299_ (.A1(_17300_),
    .A2(_17301_),
    .B1(_16923_),
    .Y(_17302_));
 sky130_fd_sc_hd__nand3_2 _44300_ (.A(_16923_),
    .B(_17300_),
    .C(_17301_),
    .Y(_17304_));
 sky130_fd_sc_hd__inv_2 _44301_ (.A(_17304_),
    .Y(_17305_));
 sky130_fd_sc_hd__o2bb2ai_1 _44302_ (.A1_N(_17287_),
    .A2_N(_17290_),
    .B1(_17302_),
    .B2(_17305_),
    .Y(_17306_));
 sky130_fd_sc_hd__nor2_1 _44303_ (.A(_17302_),
    .B(_17305_),
    .Y(_17307_));
 sky130_fd_sc_hd__nand3_1 _44304_ (.A(_17287_),
    .B(_17290_),
    .C(_17307_),
    .Y(_17308_));
 sky130_fd_sc_hd__and3_1 _44305_ (.A(_17164_),
    .B(_17306_),
    .C(_17308_),
    .X(_17309_));
 sky130_fd_sc_hd__a21oi_1 _44306_ (.A1(_17306_),
    .A2(_17308_),
    .B1(_17164_),
    .Y(_17310_));
 sky130_fd_sc_hd__clkbuf_2 _44307_ (.A(_09012_),
    .X(_17311_));
 sky130_fd_sc_hd__clkbuf_2 _44308_ (.A(_16846_),
    .X(_17312_));
 sky130_fd_sc_hd__o21ai_1 _44309_ (.A1(_16913_),
    .A2(_16925_),
    .B1(_16929_),
    .Y(_17313_));
 sky130_fd_sc_hd__o311a_1 _44310_ (.A1(_17311_),
    .A2(_17312_),
    .A3(net143),
    .B1(_17313_),
    .C1(_16926_),
    .X(_17315_));
 sky130_fd_sc_hd__or3_1 _44311_ (.A(_17311_),
    .B(_16846_),
    .C(net143),
    .X(_17316_));
 sky130_fd_sc_hd__a21oi_1 _44312_ (.A1(_16926_),
    .A2(_17313_),
    .B1(_17316_),
    .Y(_17317_));
 sky130_fd_sc_hd__o21bai_4 _44313_ (.A1(_17133_),
    .A2(_17134_),
    .B1_N(_17317_),
    .Y(_17318_));
 sky130_fd_sc_hd__a2111o_1 _44314_ (.A1(_16926_),
    .A2(_17313_),
    .B1(_17316_),
    .C1(_17133_),
    .D1(_17134_),
    .X(_17319_));
 sky130_fd_sc_hd__o21ai_1 _44315_ (.A1(_17315_),
    .A2(_17318_),
    .B1(_17319_),
    .Y(_17320_));
 sky130_fd_sc_hd__o21ai_1 _44316_ (.A1(_17309_),
    .A2(_17310_),
    .B1(_17320_),
    .Y(_17321_));
 sky130_fd_sc_hd__nand3_1 _44317_ (.A(_17164_),
    .B(_17306_),
    .C(_17308_),
    .Y(_17322_));
 sky130_fd_sc_hd__a21o_1 _44318_ (.A1(_17306_),
    .A2(_17308_),
    .B1(_17164_),
    .X(_17323_));
 sky130_fd_sc_hd__o2111ai_2 _44319_ (.A1(_17315_),
    .A2(_17318_),
    .B1(_17322_),
    .C1(_17323_),
    .D1(_17319_),
    .Y(_17324_));
 sky130_fd_sc_hd__a32oi_4 _44320_ (.A1(_17126_),
    .A2(_17127_),
    .A3(_17129_),
    .B1(_17144_),
    .B2(_17125_),
    .Y(_17326_));
 sky130_fd_sc_hd__a21o_1 _44321_ (.A1(_17321_),
    .A2(_17324_),
    .B1(_17326_),
    .X(_17327_));
 sky130_fd_sc_hd__nand3_2 _44322_ (.A(_17321_),
    .B(_17324_),
    .C(_17326_),
    .Y(_17328_));
 sky130_fd_sc_hd__o21a_1 _44323_ (.A1(_16884_),
    .A2(_17142_),
    .B1(_17138_),
    .X(_17329_));
 sky130_fd_sc_hd__a21o_1 _44324_ (.A1(_17327_),
    .A2(_17328_),
    .B1(_17329_),
    .X(_17330_));
 sky130_fd_sc_hd__o2111ai_2 _44325_ (.A1(_16884_),
    .A2(_17142_),
    .B1(_17138_),
    .C1(_17327_),
    .D1(_17328_),
    .Y(_17331_));
 sky130_fd_sc_hd__o21ai_1 _44326_ (.A1(_17156_),
    .A2(_17151_),
    .B1(_17154_),
    .Y(_17332_));
 sky130_fd_sc_hd__a21o_1 _44327_ (.A1(_17330_),
    .A2(_17331_),
    .B1(_17332_),
    .X(_17333_));
 sky130_fd_sc_hd__nand3_1 _44328_ (.A(_17332_),
    .B(_17330_),
    .C(_17331_),
    .Y(_17334_));
 sky130_fd_sc_hd__nand2_1 _44329_ (.A(_17333_),
    .B(_17334_),
    .Y(_17335_));
 sky130_fd_sc_hd__nand2_1 _44330_ (.A(_16907_),
    .B(_17158_),
    .Y(_17337_));
 sky130_fd_sc_hd__a21bo_1 _44331_ (.A1(_17159_),
    .A2(_17162_),
    .B1_N(_17337_),
    .X(_17338_));
 sky130_fd_sc_hd__xnor2_1 _44332_ (.A(_17335_),
    .B(_17338_),
    .Y(_00021_));
 sky130_fd_sc_hd__inv_2 _44333_ (.A(_17327_),
    .Y(_17339_));
 sky130_fd_sc_hd__a21oi_4 _44334_ (.A1(_17328_),
    .A2(_17329_),
    .B1(_17339_),
    .Y(_17340_));
 sky130_fd_sc_hd__inv_2 _44335_ (.A(net143),
    .Y(_17341_));
 sky130_fd_sc_hd__o211ai_1 _44336_ (.A1(_17311_),
    .A2(_17312_),
    .B1(_17300_),
    .C1(_17304_),
    .Y(_17342_));
 sky130_fd_sc_hd__a211o_1 _44337_ (.A1(_17300_),
    .A2(_17304_),
    .B1(_17311_),
    .C1(_17312_),
    .X(_17343_));
 sky130_fd_sc_hd__nand2_1 _44338_ (.A(_17342_),
    .B(_17343_),
    .Y(_17344_));
 sky130_fd_sc_hd__xor2_2 _44339_ (.A(_17341_),
    .B(_17344_),
    .X(_17345_));
 sky130_fd_sc_hd__nor2_1 _44340_ (.A(_16059_),
    .B(_17206_),
    .Y(_17347_));
 sky130_fd_sc_hd__inv_2 _44341_ (.A(_17200_),
    .Y(_17348_));
 sky130_fd_sc_hd__a211oi_2 _44342_ (.A1(_17173_),
    .A2(_17197_),
    .B1(_17348_),
    .C1(_16668_),
    .Y(_17349_));
 sky130_fd_sc_hd__nand2_1 _44343_ (.A(_17172_),
    .B(_17197_),
    .Y(_17350_));
 sky130_fd_sc_hd__a21oi_1 _44344_ (.A1(_17200_),
    .A2(_17350_),
    .B1(_16010_),
    .Y(_17351_));
 sky130_fd_sc_hd__o21bai_2 _44345_ (.A1(_17349_),
    .A2(_17351_),
    .B1_N(_12876_),
    .Y(_17352_));
 sky130_fd_sc_hd__a211o_1 _44346_ (.A1(_17173_),
    .A2(_17197_),
    .B1(_17348_),
    .C1(_16668_),
    .X(_17353_));
 sky130_fd_sc_hd__or2_1 _44347_ (.A(_16937_),
    .B(_17170_),
    .X(_17354_));
 sky130_fd_sc_hd__a22oi_1 _44348_ (.A1(_17199_),
    .A2(_17198_),
    .B1(_16990_),
    .B2(_17354_),
    .Y(_17355_));
 sky130_fd_sc_hd__o21ai_1 _44349_ (.A1(_17348_),
    .A2(_17355_),
    .B1(_16669_),
    .Y(_17356_));
 sky130_fd_sc_hd__nand3_2 _44350_ (.A(_12876_),
    .B(_17353_),
    .C(_17356_),
    .Y(_17358_));
 sky130_fd_sc_hd__nand3_2 _44351_ (.A(_17352_),
    .B(_17358_),
    .C(_16681_),
    .Y(_17359_));
 sky130_fd_sc_hd__o21ai_2 _44352_ (.A1(_17212_),
    .A2(_17347_),
    .B1(_17359_),
    .Y(_17360_));
 sky130_fd_sc_hd__a21oi_4 _44353_ (.A1(_17352_),
    .A2(_17358_),
    .B1(_16681_),
    .Y(_17361_));
 sky130_fd_sc_hd__a21o_1 _44354_ (.A1(_16043_),
    .A2(_17209_),
    .B1(_17212_),
    .X(_17362_));
 sky130_fd_sc_hd__inv_2 _44355_ (.A(_17359_),
    .Y(_17363_));
 sky130_fd_sc_hd__nor2_1 _44356_ (.A(_17363_),
    .B(_17361_),
    .Y(_17364_));
 sky130_fd_sc_hd__o21ai_2 _44357_ (.A1(_17220_),
    .A2(_17217_),
    .B1(_17214_),
    .Y(_17365_));
 sky130_fd_sc_hd__o221ai_4 _44358_ (.A1(_17360_),
    .A2(_17361_),
    .B1(_17362_),
    .B2(_17364_),
    .C1(_17365_),
    .Y(_17366_));
 sky130_fd_sc_hd__buf_6 _44359_ (.A(_17359_),
    .X(_17367_));
 sky130_fd_sc_hd__a21o_1 _44360_ (.A1(_17352_),
    .A2(_17358_),
    .B1(_17022_),
    .X(_17369_));
 sky130_fd_sc_hd__a21oi_1 _44361_ (.A1(_17367_),
    .A2(_17369_),
    .B1(_17362_),
    .Y(_17370_));
 sky130_fd_sc_hd__o211a_1 _44362_ (.A1(_17212_),
    .A2(_17347_),
    .B1(_17359_),
    .C1(_17369_),
    .X(_17371_));
 sky130_fd_sc_hd__o21bai_2 _44363_ (.A1(_17370_),
    .A2(_17371_),
    .B1_N(_17365_),
    .Y(_17372_));
 sky130_fd_sc_hd__inv_2 _44364_ (.A(_17238_),
    .Y(_17373_));
 sky130_fd_sc_hd__or2_1 _44365_ (.A(_17236_),
    .B(_17373_),
    .X(_17374_));
 sky130_fd_sc_hd__a21oi_2 _44366_ (.A1(_17366_),
    .A2(_17372_),
    .B1(_17374_),
    .Y(_17375_));
 sky130_fd_sc_hd__buf_6 _44367_ (.A(_17366_),
    .X(_17376_));
 sky130_fd_sc_hd__o211ai_2 _44368_ (.A1(_17236_),
    .A2(_17373_),
    .B1(_17376_),
    .C1(_17372_),
    .Y(_17377_));
 sky130_fd_sc_hd__nand3b_2 _44369_ (.A_N(_17375_),
    .B(_17377_),
    .C(_17227_),
    .Y(_17378_));
 sky130_fd_sc_hd__o211a_1 _44370_ (.A1(_17236_),
    .A2(_17373_),
    .B1(_17376_),
    .C1(_17372_),
    .X(_17380_));
 sky130_fd_sc_hd__o21ai_2 _44371_ (.A1(_17375_),
    .A2(_17380_),
    .B1(_17222_),
    .Y(_17381_));
 sky130_fd_sc_hd__or2_1 _44372_ (.A(_17268_),
    .B(_17273_),
    .X(_17382_));
 sky130_fd_sc_hd__or2_1 _44373_ (.A(_17241_),
    .B(_17275_),
    .X(_17383_));
 sky130_fd_sc_hd__or3_1 _44374_ (.A(_17094_),
    .B(_17243_),
    .C(_17247_),
    .X(_17384_));
 sky130_fd_sc_hd__o21ai_2 _44375_ (.A1(_17243_),
    .A2(_17247_),
    .B1(_17096_),
    .Y(_17385_));
 sky130_fd_sc_hd__nand2_1 _44376_ (.A(_17384_),
    .B(_17385_),
    .Y(_17386_));
 sky130_fd_sc_hd__nor2_1 _44377_ (.A(_17091_),
    .B(_17386_),
    .Y(_17387_));
 sky130_fd_sc_hd__o211a_1 _44378_ (.A1(_15599_),
    .A2(net70),
    .B1(_17090_),
    .C1(_17386_),
    .X(_17388_));
 sky130_fd_sc_hd__nor2_1 _44379_ (.A(_17387_),
    .B(_17388_),
    .Y(_17389_));
 sky130_fd_sc_hd__clkbuf_2 _44380_ (.A(_17254_),
    .X(_17391_));
 sky130_fd_sc_hd__mux2_1 _44381_ (.A0(_17257_),
    .A1(net214),
    .S(_17049_),
    .X(_17392_));
 sky130_fd_sc_hd__xnor2_1 _44382_ (.A(_17391_),
    .B(_17392_),
    .Y(_17393_));
 sky130_fd_sc_hd__inv_2 _44383_ (.A(_17391_),
    .Y(_17394_));
 sky130_fd_sc_hd__a21oi_2 _44384_ (.A1(_17262_),
    .A2(_17394_),
    .B1(_17261_),
    .Y(_17395_));
 sky130_fd_sc_hd__nor2_1 _44385_ (.A(_17393_),
    .B(_17395_),
    .Y(_17396_));
 sky130_fd_sc_hd__and2_1 _44386_ (.A(_17395_),
    .B(_17393_),
    .X(_17397_));
 sky130_fd_sc_hd__a21oi_2 _44387_ (.A1(_17253_),
    .A2(_17250_),
    .B1(_17252_),
    .Y(_17398_));
 sky130_fd_sc_hd__nand2_1 _44388_ (.A(_17076_),
    .B(_17398_),
    .Y(_17399_));
 sky130_fd_sc_hd__inv_2 _44389_ (.A(_17399_),
    .Y(_17400_));
 sky130_fd_sc_hd__nor2_1 _44390_ (.A(_17398_),
    .B(_17076_),
    .Y(_17402_));
 sky130_fd_sc_hd__a21o_1 _44391_ (.A1(_17245_),
    .A2(_17399_),
    .B1(_17402_),
    .X(_17403_));
 sky130_fd_sc_hd__o21ai_1 _44392_ (.A1(_17402_),
    .A2(_17400_),
    .B1(_17245_),
    .Y(_17404_));
 sky130_fd_sc_hd__o21a_1 _44393_ (.A1(_17400_),
    .A2(_17403_),
    .B1(_17404_),
    .X(_17405_));
 sky130_fd_sc_hd__buf_1 _44394_ (.A(_17405_),
    .X(_17406_));
 sky130_fd_sc_hd__o21a_1 _44395_ (.A1(_17396_),
    .A2(_17397_),
    .B1(_17406_),
    .X(_17407_));
 sky130_fd_sc_hd__a21oi_1 _44396_ (.A1(_17393_),
    .A2(_17395_),
    .B1(_17405_),
    .Y(_17408_));
 sky130_fd_sc_hd__o21a_1 _44397_ (.A1(_17393_),
    .A2(_17395_),
    .B1(_17408_),
    .X(_17409_));
 sky130_fd_sc_hd__a211oi_2 _44398_ (.A1(_17266_),
    .A2(_17272_),
    .B1(_17407_),
    .C1(_17409_),
    .Y(_17410_));
 sky130_fd_sc_hd__o211a_1 _44399_ (.A1(_17407_),
    .A2(_17409_),
    .B1(_17266_),
    .C1(_17272_),
    .X(_17411_));
 sky130_fd_sc_hd__nor2_1 _44400_ (.A(_17410_),
    .B(_17411_),
    .Y(_17413_));
 sky130_fd_sc_hd__or3b_1 _44401_ (.A(_17410_),
    .B(_17411_),
    .C_N(_17389_),
    .X(_17414_));
 sky130_fd_sc_hd__o21ai_1 _44402_ (.A1(_17389_),
    .A2(_17413_),
    .B1(_17414_),
    .Y(_17415_));
 sky130_fd_sc_hd__a21oi_1 _44403_ (.A1(_17382_),
    .A2(_17383_),
    .B1(_17415_),
    .Y(_17416_));
 sky130_fd_sc_hd__and3_1 _44404_ (.A(_17382_),
    .B(_17383_),
    .C(_17415_),
    .X(_17417_));
 sky130_fd_sc_hd__o2bb2ai_1 _44405_ (.A1_N(_17378_),
    .A2_N(_17381_),
    .B1(_17416_),
    .B2(_17417_),
    .Y(_17418_));
 sky130_fd_sc_hd__nor2_1 _44406_ (.A(_17416_),
    .B(_17417_),
    .Y(_17419_));
 sky130_fd_sc_hd__nand3_1 _44407_ (.A(_17378_),
    .B(_17381_),
    .C(_17419_),
    .Y(_17420_));
 sky130_fd_sc_hd__nand2_1 _44408_ (.A(_17418_),
    .B(_17420_),
    .Y(_17421_));
 sky130_fd_sc_hd__a32oi_1 _44409_ (.A1(_17233_),
    .A2(_17283_),
    .A3(_17284_),
    .B1(_17277_),
    .B2(_17279_),
    .Y(_17422_));
 sky130_fd_sc_hd__nand2_1 _44410_ (.A(_17421_),
    .B(_17422_),
    .Y(_17424_));
 sky130_fd_sc_hd__clkbuf_2 _44411_ (.A(_17420_),
    .X(_17425_));
 sky130_fd_sc_hd__nand2_1 _44412_ (.A(_17280_),
    .B(_17285_),
    .Y(_17426_));
 sky130_fd_sc_hd__nand3_2 _44413_ (.A(_17418_),
    .B(_17425_),
    .C(_17426_),
    .Y(_17427_));
 sky130_fd_sc_hd__and4_1 _44414_ (.A(_16716_),
    .B(_16519_),
    .C(_16322_),
    .D(_13293_),
    .X(_17428_));
 sky130_fd_sc_hd__nand2_1 _44415_ (.A(_17230_),
    .B(_17028_),
    .Y(_17429_));
 sky130_fd_sc_hd__xnor2_2 _44416_ (.A(_16849_),
    .B(_16917_),
    .Y(_17430_));
 sky130_fd_sc_hd__nand3_1 _44417_ (.A(_17225_),
    .B(_17429_),
    .C(_17430_),
    .Y(_17431_));
 sky130_fd_sc_hd__a21o_1 _44418_ (.A1(_17225_),
    .A2(_17429_),
    .B1(_17430_),
    .X(_17432_));
 sky130_fd_sc_hd__o211ai_1 _44419_ (.A1(_17296_),
    .A2(_17428_),
    .B1(_17431_),
    .C1(_17432_),
    .Y(_17433_));
 sky130_fd_sc_hd__o311a_1 _44420_ (.A1(_17229_),
    .A2(_17227_),
    .A3(_17228_),
    .B1(_17430_),
    .C1(_17429_),
    .X(_17435_));
 sky130_fd_sc_hd__a21oi_1 _44421_ (.A1(_17225_),
    .A2(_17429_),
    .B1(_17430_),
    .Y(_17436_));
 sky130_fd_sc_hd__nor2_1 _44422_ (.A(_17296_),
    .B(_17428_),
    .Y(_17437_));
 sky130_fd_sc_hd__o21ai_1 _44423_ (.A1(_17435_),
    .A2(_17436_),
    .B1(_17437_),
    .Y(_17438_));
 sky130_fd_sc_hd__nand2_1 _44424_ (.A(_17433_),
    .B(_17438_),
    .Y(_17439_));
 sky130_fd_sc_hd__a21oi_1 _44425_ (.A1(_17424_),
    .A2(_17427_),
    .B1(_17439_),
    .Y(_17440_));
 sky130_fd_sc_hd__nor3_1 _44426_ (.A(_17437_),
    .B(_17435_),
    .C(_17436_),
    .Y(_17441_));
 sky130_fd_sc_hd__o21a_1 _44427_ (.A1(_17435_),
    .A2(_17436_),
    .B1(_17437_),
    .X(_17442_));
 sky130_fd_sc_hd__o211a_1 _44428_ (.A1(_17441_),
    .A2(_17442_),
    .B1(_17424_),
    .C1(_17427_),
    .X(_17443_));
 sky130_fd_sc_hd__a32o_1 _44429_ (.A1(_17167_),
    .A2(_17285_),
    .A3(_17286_),
    .B1(_17290_),
    .B2(_17307_),
    .X(_17444_));
 sky130_fd_sc_hd__o21ai_1 _44430_ (.A1(_17440_),
    .A2(_17443_),
    .B1(_17444_),
    .Y(_17446_));
 sky130_fd_sc_hd__o211ai_1 _44431_ (.A1(_17441_),
    .A2(_17442_),
    .B1(_17424_),
    .C1(_17427_),
    .Y(_17447_));
 sky130_fd_sc_hd__a32oi_2 _44432_ (.A1(_17167_),
    .A2(_17285_),
    .A3(_17286_),
    .B1(_17290_),
    .B2(_17307_),
    .Y(_17448_));
 sky130_fd_sc_hd__nand3b_2 _44433_ (.A_N(_17440_),
    .B(_17447_),
    .C(_17448_),
    .Y(_17449_));
 sky130_fd_sc_hd__nand3b_1 _44434_ (.A_N(_17345_),
    .B(_17446_),
    .C(_17449_),
    .Y(_17450_));
 sky130_fd_sc_hd__nand2_1 _44435_ (.A(_17446_),
    .B(_17449_),
    .Y(_17451_));
 sky130_fd_sc_hd__nand2_1 _44436_ (.A(_17451_),
    .B(_17345_),
    .Y(_17452_));
 sky130_fd_sc_hd__o21ai_1 _44437_ (.A1(_17320_),
    .A2(_17309_),
    .B1(_17323_),
    .Y(_17453_));
 sky130_fd_sc_hd__a21oi_1 _44438_ (.A1(_17450_),
    .A2(_17452_),
    .B1(_17453_),
    .Y(_17454_));
 sky130_fd_sc_hd__and3_1 _44439_ (.A(_17453_),
    .B(_17450_),
    .C(_17452_),
    .X(_17455_));
 sky130_fd_sc_hd__nor2_2 _44440_ (.A(_17454_),
    .B(_17455_),
    .Y(_17457_));
 sky130_fd_sc_hd__xnor2_4 _44441_ (.A(_17318_),
    .B(_17457_),
    .Y(_17458_));
 sky130_fd_sc_hd__xor2_2 _44442_ (.A(_17340_),
    .B(_17458_),
    .X(_17459_));
 sky130_fd_sc_hd__nand3_1 _44443_ (.A(_17333_),
    .B(_17334_),
    .C(_17159_),
    .Y(_17460_));
 sky130_fd_sc_hd__a21oi_2 _44444_ (.A1(_16564_),
    .A2(_16548_),
    .B1(_17160_),
    .Y(_17461_));
 sky130_fd_sc_hd__a21bo_1 _44445_ (.A1(_17337_),
    .A2(_17334_),
    .B1_N(_17333_),
    .X(_17462_));
 sky130_fd_sc_hd__o31ai_4 _44446_ (.A1(_16902_),
    .A2(_17460_),
    .A3(_17461_),
    .B1(_17462_),
    .Y(_17463_));
 sky130_fd_sc_hd__nor2_1 _44447_ (.A(_17459_),
    .B(_17463_),
    .Y(_17464_));
 sky130_fd_sc_hd__nand2_1 _44448_ (.A(_17463_),
    .B(_17459_),
    .Y(_17465_));
 sky130_fd_sc_hd__and2b_1 _44449_ (.A_N(_17464_),
    .B(_17465_),
    .X(_17466_));
 sky130_fd_sc_hd__clkbuf_1 _44450_ (.A(_17466_),
    .X(_00022_));
 sky130_fd_sc_hd__a21oi_1 _44451_ (.A1(_17418_),
    .A2(_17425_),
    .B1(_17426_),
    .Y(_17468_));
 sky130_fd_sc_hd__o21ai_2 _44452_ (.A1(_17468_),
    .A2(_17439_),
    .B1(_17427_),
    .Y(_17469_));
 sky130_fd_sc_hd__nand2_1 _44453_ (.A(_17378_),
    .B(_17381_),
    .Y(_17470_));
 sky130_fd_sc_hd__inv_2 _44454_ (.A(_17385_),
    .Y(_17471_));
 sky130_fd_sc_hd__clkbuf_2 _44455_ (.A(_17351_),
    .X(_17472_));
 sky130_fd_sc_hd__nor2_1 _44456_ (.A(_16059_),
    .B(_17472_),
    .Y(_17473_));
 sky130_fd_sc_hd__a2bb2o_1 _44457_ (.A1_N(_17349_),
    .A2_N(_17473_),
    .B1(_17367_),
    .B2(_17369_),
    .X(_17474_));
 sky130_fd_sc_hd__o2111ai_1 _44458_ (.A1(_17472_),
    .A2(_16716_),
    .B1(_17353_),
    .C1(_17367_),
    .D1(_17369_),
    .Y(_17475_));
 sky130_fd_sc_hd__a21oi_1 _44459_ (.A1(_17367_),
    .A2(_17362_),
    .B1(_17361_),
    .Y(_17476_));
 sky130_fd_sc_hd__nand3_2 _44460_ (.A(_17474_),
    .B(_17475_),
    .C(_17476_),
    .Y(_17478_));
 sky130_fd_sc_hd__inv_2 _44461_ (.A(_17360_),
    .Y(_17479_));
 sky130_fd_sc_hd__a2bb2oi_1 _44462_ (.A1_N(_17349_),
    .A2_N(_17473_),
    .B1(_17367_),
    .B2(_17369_),
    .Y(_17480_));
 sky130_fd_sc_hd__a31o_1 _44463_ (.A1(_17008_),
    .A2(_17200_),
    .A3(_17350_),
    .B1(_17473_),
    .X(_17481_));
 sky130_fd_sc_hd__nor3_1 _44464_ (.A(_17361_),
    .B(_17481_),
    .C(_17363_),
    .Y(_17482_));
 sky130_fd_sc_hd__o22ai_2 _44465_ (.A1(_17361_),
    .A2(_17479_),
    .B1(_17480_),
    .B2(_17482_),
    .Y(_17483_));
 sky130_fd_sc_hd__o211a_1 _44466_ (.A1(_17471_),
    .A2(_17387_),
    .B1(_17478_),
    .C1(_17483_),
    .X(_17484_));
 sky130_fd_sc_hd__buf_4 _44467_ (.A(_17483_),
    .X(_17485_));
 sky130_fd_sc_hd__o21ai_2 _44468_ (.A1(_17092_),
    .A2(_17386_),
    .B1(_17385_),
    .Y(_17486_));
 sky130_fd_sc_hd__a21oi_2 _44469_ (.A1(_17478_),
    .A2(_17485_),
    .B1(_17486_),
    .Y(_17487_));
 sky130_fd_sc_hd__o21bai_4 _44470_ (.A1(_17484_),
    .A2(_17487_),
    .B1_N(_17376_),
    .Y(_17489_));
 sky130_fd_sc_hd__o211ai_2 _44471_ (.A1(_17471_),
    .A2(_17387_),
    .B1(_17478_),
    .C1(_17485_),
    .Y(_17490_));
 sky130_fd_sc_hd__a21o_1 _44472_ (.A1(_17478_),
    .A2(_17485_),
    .B1(_17486_),
    .X(_17491_));
 sky130_fd_sc_hd__nand3_2 _44473_ (.A(_17376_),
    .B(_17490_),
    .C(_17491_),
    .Y(_17492_));
 sky130_fd_sc_hd__inv_2 _44474_ (.A(_17411_),
    .Y(_17493_));
 sky130_fd_sc_hd__a21oi_2 _44475_ (.A1(_17493_),
    .A2(_17389_),
    .B1(_17410_),
    .Y(_17494_));
 sky130_fd_sc_hd__and3_1 _44476_ (.A(_17049_),
    .B(_17391_),
    .C(net214),
    .X(_17495_));
 sky130_fd_sc_hd__a41o_1 _44477_ (.A1(_17044_),
    .A2(_17045_),
    .A3(_17394_),
    .A4(_17257_),
    .B1(_17495_),
    .X(_17496_));
 sky130_fd_sc_hd__xor2_1 _44478_ (.A(_17406_),
    .B(_17496_),
    .X(_17497_));
 sky130_fd_sc_hd__nor3_1 _44479_ (.A(_17396_),
    .B(_17408_),
    .C(_17497_),
    .Y(_17498_));
 sky130_fd_sc_hd__inv_2 _44480_ (.A(_17498_),
    .Y(_17500_));
 sky130_fd_sc_hd__nand2_1 _44481_ (.A(_17096_),
    .B(_17403_),
    .Y(_17501_));
 sky130_fd_sc_hd__a211o_1 _44482_ (.A1(_17245_),
    .A2(_17399_),
    .B1(_17402_),
    .C1(_17094_),
    .X(_17502_));
 sky130_fd_sc_hd__nand2_1 _44483_ (.A(_17501_),
    .B(_17502_),
    .Y(_17503_));
 sky130_fd_sc_hd__xnor2_1 _44484_ (.A(_17091_),
    .B(_17503_),
    .Y(_17504_));
 sky130_fd_sc_hd__clkbuf_2 _44485_ (.A(_17504_),
    .X(_17505_));
 sky130_fd_sc_hd__o21ai_1 _44486_ (.A1(_17396_),
    .A2(_17408_),
    .B1(_17497_),
    .Y(_17506_));
 sky130_fd_sc_hd__o21a_1 _44487_ (.A1(_17505_),
    .A2(_17498_),
    .B1(_17506_),
    .X(_17507_));
 sky130_fd_sc_hd__a21oi_1 _44488_ (.A1(_17506_),
    .A2(_17500_),
    .B1(_17505_),
    .Y(_17508_));
 sky130_fd_sc_hd__a21oi_2 _44489_ (.A1(_17500_),
    .A2(_17507_),
    .B1(_17508_),
    .Y(_17509_));
 sky130_fd_sc_hd__nor2_2 _44490_ (.A(_17494_),
    .B(_17509_),
    .Y(_17511_));
 sky130_fd_sc_hd__and2_1 _44491_ (.A(_17494_),
    .B(_17509_),
    .X(_17512_));
 sky130_fd_sc_hd__or2_1 _44492_ (.A(_17511_),
    .B(_17512_),
    .X(_17513_));
 sky130_fd_sc_hd__a21oi_4 _44493_ (.A1(_17489_),
    .A2(_17492_),
    .B1(_17513_),
    .Y(_17514_));
 sky130_fd_sc_hd__o211a_2 _44494_ (.A1(_17511_),
    .A2(_17512_),
    .B1(_17489_),
    .C1(_17492_),
    .X(_17515_));
 sky130_fd_sc_hd__a21o_1 _44495_ (.A1(_17382_),
    .A2(_17383_),
    .B1(_17415_),
    .X(_17516_));
 sky130_fd_sc_hd__o221ai_2 _44496_ (.A1(_17417_),
    .A2(_17470_),
    .B1(_17514_),
    .B2(_17515_),
    .C1(_17516_),
    .Y(_17517_));
 sky130_fd_sc_hd__a211o_1 _44497_ (.A1(_17516_),
    .A2(_17425_),
    .B1(_17515_),
    .C1(_17514_),
    .X(_17518_));
 sky130_fd_sc_hd__o21ai_2 _44498_ (.A1(_17222_),
    .A2(_17375_),
    .B1(_17377_),
    .Y(_17519_));
 sky130_fd_sc_hd__clkbuf_2 _44499_ (.A(_16934_),
    .X(_17520_));
 sky130_fd_sc_hd__or2_1 _44500_ (.A(_16519_),
    .B(_16914_),
    .X(_17522_));
 sky130_fd_sc_hd__nor2_2 _44501_ (.A(_17520_),
    .B(_17522_),
    .Y(_17523_));
 sky130_fd_sc_hd__xnor2_2 _44502_ (.A(_17519_),
    .B(_17523_),
    .Y(_17524_));
 sky130_fd_sc_hd__nand3_1 _44503_ (.A(_17517_),
    .B(_17518_),
    .C(_17524_),
    .Y(_17525_));
 sky130_fd_sc_hd__o211ai_1 _44504_ (.A1(_17511_),
    .A2(_17512_),
    .B1(_17489_),
    .C1(_17492_),
    .Y(_17526_));
 sky130_fd_sc_hd__a21o_2 _44505_ (.A1(_17489_),
    .A2(_17492_),
    .B1(_17513_),
    .X(_17527_));
 sky130_fd_sc_hd__nand2_1 _44506_ (.A(_17516_),
    .B(_17425_),
    .Y(_17528_));
 sky130_fd_sc_hd__a21oi_1 _44507_ (.A1(_17526_),
    .A2(_17527_),
    .B1(_17528_),
    .Y(_17529_));
 sky130_fd_sc_hd__a211oi_4 _44508_ (.A1(_17516_),
    .A2(_17425_),
    .B1(_17515_),
    .C1(_17514_),
    .Y(_17530_));
 sky130_fd_sc_hd__o21bai_2 _44509_ (.A1(_17529_),
    .A2(_17530_),
    .B1_N(_17524_),
    .Y(_17531_));
 sky130_fd_sc_hd__and3_1 _44510_ (.A(_17469_),
    .B(_17525_),
    .C(_17531_),
    .X(_17533_));
 sky130_fd_sc_hd__a21oi_1 _44511_ (.A1(_17525_),
    .A2(_17531_),
    .B1(_17469_),
    .Y(_17534_));
 sky130_fd_sc_hd__a21o_1 _44512_ (.A1(_10304_),
    .A2(_16914_),
    .B1(_16519_),
    .X(_17535_));
 sky130_fd_sc_hd__o21ai_2 _44513_ (.A1(_17437_),
    .A2(_17435_),
    .B1(_17432_),
    .Y(_17536_));
 sky130_fd_sc_hd__xnor2_1 _44514_ (.A(_17535_),
    .B(_17536_),
    .Y(_17537_));
 sky130_fd_sc_hd__o21ai_1 _44515_ (.A1(_17533_),
    .A2(_17534_),
    .B1(_17537_),
    .Y(_17538_));
 sky130_fd_sc_hd__a21o_1 _44516_ (.A1(_17525_),
    .A2(_17531_),
    .B1(_17469_),
    .X(_17539_));
 sky130_fd_sc_hd__nand3_1 _44517_ (.A(_17469_),
    .B(_17525_),
    .C(_17531_),
    .Y(_17540_));
 sky130_fd_sc_hd__nand3b_1 _44518_ (.A_N(_17537_),
    .B(_17539_),
    .C(_17540_),
    .Y(_17541_));
 sky130_fd_sc_hd__nand2_2 _44519_ (.A(_17538_),
    .B(_17541_),
    .Y(_17542_));
 sky130_fd_sc_hd__a21boi_4 _44520_ (.A1(_17345_),
    .A2(_17449_),
    .B1_N(_17446_),
    .Y(_17544_));
 sky130_fd_sc_hd__nand2_1 _44521_ (.A(_17542_),
    .B(_17544_),
    .Y(_17545_));
 sky130_fd_sc_hd__nand3b_1 _44522_ (.A_N(_17544_),
    .B(_17538_),
    .C(_17541_),
    .Y(_17546_));
 sky130_fd_sc_hd__o21ai_2 _44523_ (.A1(_17341_),
    .A2(_17344_),
    .B1(_17343_),
    .Y(_17547_));
 sky130_fd_sc_hd__a21o_1 _44524_ (.A1(_17545_),
    .A2(_17546_),
    .B1(_17547_),
    .X(_17548_));
 sky130_fd_sc_hd__a21boi_1 _44525_ (.A1(_17542_),
    .A2(_17544_),
    .B1_N(_17547_),
    .Y(_17549_));
 sky130_fd_sc_hd__o21ai_2 _44526_ (.A1(_17544_),
    .A2(_17542_),
    .B1(_17549_),
    .Y(_17550_));
 sky130_fd_sc_hd__nand3_1 _44527_ (.A(_17453_),
    .B(_17450_),
    .C(_17452_),
    .Y(_17551_));
 sky130_fd_sc_hd__a21oi_1 _44528_ (.A1(_17318_),
    .A2(_17551_),
    .B1(_17454_),
    .Y(_17552_));
 sky130_fd_sc_hd__a21boi_1 _44529_ (.A1(_17548_),
    .A2(_17550_),
    .B1_N(_17552_),
    .Y(_17553_));
 sky130_fd_sc_hd__nand3b_2 _44530_ (.A_N(_17552_),
    .B(_17548_),
    .C(_17550_),
    .Y(_17555_));
 sky130_fd_sc_hd__o211ai_2 _44531_ (.A1(_17458_),
    .A2(_17340_),
    .B1(_17555_),
    .C1(_17465_),
    .Y(_17556_));
 sky130_fd_sc_hd__o21ai_1 _44532_ (.A1(_17340_),
    .A2(_17458_),
    .B1(_17465_),
    .Y(_17557_));
 sky130_fd_sc_hd__a21bo_1 _44533_ (.A1(_17548_),
    .A2(_17550_),
    .B1_N(_17552_),
    .X(_17558_));
 sky130_fd_sc_hd__nand2_1 _44534_ (.A(_17558_),
    .B(_17555_),
    .Y(_17559_));
 sky130_fd_sc_hd__a2bb2o_1 _44535_ (.A1_N(_17553_),
    .A2_N(_17556_),
    .B1(_17557_),
    .B2(_17559_),
    .X(_00023_));
 sky130_fd_sc_hd__inv_2 _44536_ (.A(_17546_),
    .Y(_17560_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44537_ (.A(_16519_),
    .X(_17561_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44538_ (.A(_16914_),
    .X(_17562_));
 sky130_fd_sc_hd__o22a_1 _44539_ (.A1(_17561_),
    .A2(_17562_),
    .B1(_17311_),
    .B2(_17536_),
    .X(_17563_));
 sky130_fd_sc_hd__o311a_2 _44540_ (.A1(_14857_),
    .A2(_14605_),
    .A3(_14607_),
    .B1(_16018_),
    .C1(_16707_),
    .X(_17565_));
 sky130_fd_sc_hd__o21a_1 _44541_ (.A1(_17011_),
    .A2(_17012_),
    .B1(_16934_),
    .X(_17566_));
 sky130_fd_sc_hd__nor2_1 _44542_ (.A(_17403_),
    .B(_17096_),
    .Y(_17567_));
 sky130_fd_sc_hd__o21a_1 _44543_ (.A1(_17092_),
    .A2(_17567_),
    .B1(_17501_),
    .X(_17568_));
 sky130_fd_sc_hd__a221o_2 _44544_ (.A1(_17472_),
    .A2(_17565_),
    .B1(_17566_),
    .B2(_17349_),
    .C1(_17568_),
    .X(_17569_));
 sky130_fd_sc_hd__or4_1 _44545_ (.A(_16043_),
    .B(_17011_),
    .C(_17012_),
    .D(_17356_),
    .X(_17570_));
 sky130_fd_sc_hd__or3_1 _44546_ (.A(_16707_),
    .B(_17022_),
    .C(_17353_),
    .X(_17571_));
 sky130_fd_sc_hd__a21bo_1 _44547_ (.A1(_17570_),
    .A2(_17571_),
    .B1_N(_17568_),
    .X(_17572_));
 sky130_fd_sc_hd__nand2_1 _44548_ (.A(_17569_),
    .B(_17572_),
    .Y(_17573_));
 sky130_fd_sc_hd__nand2_1 _44549_ (.A(_17485_),
    .B(_17573_),
    .Y(_17574_));
 sky130_fd_sc_hd__nand3b_2 _44550_ (.A_N(_17483_),
    .B(_17569_),
    .C(_17572_),
    .Y(_17576_));
 sky130_fd_sc_hd__and4_2 _44551_ (.A(_17406_),
    .B(_17391_),
    .C(_17049_),
    .D(net214),
    .X(_17577_));
 sky130_fd_sc_hd__or3b_1 _44552_ (.A(_17049_),
    .B(_17391_),
    .C_N(_17257_),
    .X(_17578_));
 sky130_fd_sc_hd__nor2_1 _44553_ (.A(_17578_),
    .B(_17406_),
    .Y(_17579_));
 sky130_fd_sc_hd__o21ai_1 _44554_ (.A1(_17577_),
    .A2(_17579_),
    .B1(_17504_),
    .Y(_17580_));
 sky130_fd_sc_hd__or3_1 _44555_ (.A(_17577_),
    .B(_17579_),
    .C(_17504_),
    .X(_17581_));
 sky130_fd_sc_hd__nand2_1 _44556_ (.A(_17580_),
    .B(_17581_),
    .Y(_17582_));
 sky130_fd_sc_hd__or2_1 _44557_ (.A(_17507_),
    .B(_17582_),
    .X(_17583_));
 sky130_fd_sc_hd__nand2_1 _44558_ (.A(_17582_),
    .B(_17507_),
    .Y(_17584_));
 sky130_fd_sc_hd__and2_1 _44559_ (.A(_17583_),
    .B(_17584_),
    .X(_17585_));
 sky130_fd_sc_hd__a21o_1 _44560_ (.A1(_17574_),
    .A2(_17576_),
    .B1(_17585_),
    .X(_17587_));
 sky130_fd_sc_hd__nand3_2 _44561_ (.A(_17574_),
    .B(_17576_),
    .C(_17585_),
    .Y(_17588_));
 sky130_fd_sc_hd__nand2_2 _44562_ (.A(_17587_),
    .B(_17588_),
    .Y(_17589_));
 sky130_fd_sc_hd__o211ai_2 _44563_ (.A1(_17494_),
    .A2(_17509_),
    .B1(_17527_),
    .C1(_17589_),
    .Y(_17590_));
 sky130_fd_sc_hd__o21bai_2 _44564_ (.A1(_17511_),
    .A2(_17514_),
    .B1_N(_17589_),
    .Y(_17591_));
 sky130_fd_sc_hd__o21a_1 _44565_ (.A1(_17376_),
    .A2(_17487_),
    .B1(_17490_),
    .X(_17592_));
 sky130_fd_sc_hd__a22oi_1 _44566_ (.A1(_16597_),
    .A2(_17178_),
    .B1(_17176_),
    .B2(_17187_),
    .Y(_17593_));
 sky130_fd_sc_hd__o32a_2 _44567_ (.A1(_15332_),
    .A2(_15329_),
    .A3(_17178_),
    .B1(_17177_),
    .B2(_17593_),
    .X(_17594_));
 sky130_fd_sc_hd__o21ai_1 _44568_ (.A1(_16943_),
    .A2(_16946_),
    .B1(_17175_),
    .Y(_17595_));
 sky130_fd_sc_hd__xnor2_1 _44569_ (.A(_17194_),
    .B(_17595_),
    .Y(_17596_));
 sky130_fd_sc_hd__xor2_2 _44570_ (.A(_16966_),
    .B(_17596_),
    .X(_17598_));
 sky130_fd_sc_hd__xnor2_4 _44571_ (.A(_17594_),
    .B(_17598_),
    .Y(_17599_));
 sky130_fd_sc_hd__nand2_1 _44572_ (.A(_17599_),
    .B(_17198_),
    .Y(_17600_));
 sky130_fd_sc_hd__or2_1 _44573_ (.A(_17198_),
    .B(_17599_),
    .X(_17601_));
 sky130_fd_sc_hd__nand2_1 _44574_ (.A(_17600_),
    .B(_17601_),
    .Y(_17602_));
 sky130_fd_sc_hd__xnor2_1 _44575_ (.A(_17173_),
    .B(_17602_),
    .Y(_17603_));
 sky130_fd_sc_hd__o21ai_2 _44576_ (.A1(_16671_),
    .A2(_16672_),
    .B1(_17603_),
    .Y(_17604_));
 sky130_fd_sc_hd__o21ai_1 _44577_ (.A1(_17008_),
    .A2(_17603_),
    .B1(_16934_),
    .Y(_17605_));
 sky130_fd_sc_hd__nand2_1 _44578_ (.A(_17173_),
    .B(_17600_),
    .Y(_17606_));
 sky130_fd_sc_hd__a21oi_1 _44579_ (.A1(_17601_),
    .A2(_17606_),
    .B1(_17008_),
    .Y(_17607_));
 sky130_fd_sc_hd__o221a_1 _44580_ (.A1(_16671_),
    .A2(_16672_),
    .B1(_17198_),
    .B2(_17599_),
    .C1(_17606_),
    .X(_17609_));
 sky130_fd_sc_hd__nor2_1 _44581_ (.A(_17607_),
    .B(_17609_),
    .Y(_17610_));
 sky130_fd_sc_hd__or3b_1 _44582_ (.A(_17565_),
    .B(_17566_),
    .C_N(_17610_),
    .X(_17611_));
 sky130_fd_sc_hd__o21bai_1 _44583_ (.A1(_17565_),
    .A2(_17566_),
    .B1_N(_17610_),
    .Y(_17612_));
 sky130_fd_sc_hd__a22o_1 _44584_ (.A1(_17604_),
    .A2(_17605_),
    .B1(_17611_),
    .B2(_17612_),
    .X(_17613_));
 sky130_fd_sc_hd__nand4_1 _44585_ (.A(_17604_),
    .B(_17605_),
    .C(_17611_),
    .D(_17612_),
    .Y(_17614_));
 sky130_fd_sc_hd__inv_2 _44586_ (.A(_17604_),
    .Y(_17615_));
 sky130_fd_sc_hd__nor2_1 _44587_ (.A(_17008_),
    .B(_17603_),
    .Y(_17616_));
 sky130_fd_sc_hd__nor2_1 _44588_ (.A(_17615_),
    .B(_17616_),
    .Y(_17617_));
 sky130_fd_sc_hd__o221a_1 _44589_ (.A1(_17605_),
    .A2(_17615_),
    .B1(_16934_),
    .B2(_17617_),
    .C1(_17005_),
    .X(_17618_));
 sky130_fd_sc_hd__a21oi_1 _44590_ (.A1(_17219_),
    .A2(_17211_),
    .B1(_17618_),
    .Y(_17620_));
 sky130_fd_sc_hd__a21oi_1 _44591_ (.A1(_17613_),
    .A2(_17614_),
    .B1(_17620_),
    .Y(_17621_));
 sky130_fd_sc_hd__o21ai_1 _44592_ (.A1(_17484_),
    .A2(_17621_),
    .B1(_17491_),
    .Y(_17622_));
 sky130_fd_sc_hd__nand2_1 _44593_ (.A(_17622_),
    .B(_17523_),
    .Y(_17623_));
 sky130_fd_sc_hd__o21ai_2 _44594_ (.A1(_17592_),
    .A2(_17523_),
    .B1(_17623_),
    .Y(_17624_));
 sky130_fd_sc_hd__nand3_2 _44595_ (.A(_17590_),
    .B(_17591_),
    .C(_17624_),
    .Y(_17625_));
 sky130_fd_sc_hd__a21o_1 _44596_ (.A1(_17590_),
    .A2(_17591_),
    .B1(_17624_),
    .X(_17626_));
 sky130_fd_sc_hd__nor2_1 _44597_ (.A(_17515_),
    .B(_17514_),
    .Y(_17627_));
 sky130_fd_sc_hd__o21a_1 _44598_ (.A1(_17528_),
    .A2(_17627_),
    .B1(_17524_),
    .X(_17628_));
 sky130_fd_sc_hd__o2bb2ai_4 _44599_ (.A1_N(_17625_),
    .A2_N(_17626_),
    .B1(_17628_),
    .B2(_17530_),
    .Y(_17629_));
 sky130_fd_sc_hd__a21oi_1 _44600_ (.A1(_17517_),
    .A2(_17524_),
    .B1(_17530_),
    .Y(_17631_));
 sky130_fd_sc_hd__nand3_2 _44601_ (.A(_17631_),
    .B(_17626_),
    .C(_17625_),
    .Y(_17632_));
 sky130_fd_sc_hd__clkbuf_2 _44602_ (.A(_17522_),
    .X(_17633_));
 sky130_fd_sc_hd__clkbuf_2 _44603_ (.A(_17519_),
    .X(_17634_));
 sky130_fd_sc_hd__a21oi_1 _44604_ (.A1(_17634_),
    .A2(_17520_),
    .B1(_17633_),
    .Y(_17635_));
 sky130_fd_sc_hd__a21oi_2 _44605_ (.A1(_17633_),
    .A2(_17634_),
    .B1(_17635_),
    .Y(_17636_));
 sky130_fd_sc_hd__a21oi_1 _44606_ (.A1(_17629_),
    .A2(_17632_),
    .B1(_17636_),
    .Y(_17637_));
 sky130_fd_sc_hd__and3_1 _44607_ (.A(_17629_),
    .B(_17632_),
    .C(_17636_),
    .X(_17638_));
 sky130_fd_sc_hd__o21a_1 _44608_ (.A1(_17537_),
    .A2(_17534_),
    .B1(_17540_),
    .X(_17639_));
 sky130_fd_sc_hd__o21ai_2 _44609_ (.A1(_17637_),
    .A2(_17638_),
    .B1(_17639_),
    .Y(_17640_));
 sky130_fd_sc_hd__o2bb2a_1 _44610_ (.A1_N(_17625_),
    .A2_N(_17626_),
    .B1(_17628_),
    .B2(_17530_),
    .X(_17642_));
 sky130_fd_sc_hd__nand2_2 _44611_ (.A(_17632_),
    .B(_17636_),
    .Y(_17643_));
 sky130_fd_sc_hd__a21o_1 _44612_ (.A1(_17629_),
    .A2(_17632_),
    .B1(_17636_),
    .X(_17644_));
 sky130_fd_sc_hd__o21ai_1 _44613_ (.A1(_17537_),
    .A2(_17534_),
    .B1(_17540_),
    .Y(_17645_));
 sky130_fd_sc_hd__o211ai_2 _44614_ (.A1(_17642_),
    .A2(_17643_),
    .B1(_17644_),
    .C1(_17645_),
    .Y(_17646_));
 sky130_fd_sc_hd__nand3b_2 _44615_ (.A_N(_17563_),
    .B(_17640_),
    .C(_17646_),
    .Y(_17647_));
 sky130_fd_sc_hd__a21bo_1 _44616_ (.A1(_17640_),
    .A2(_17646_),
    .B1_N(_17563_),
    .X(_17648_));
 sky130_fd_sc_hd__nand2_1 _44617_ (.A(_17647_),
    .B(_17648_),
    .Y(_17649_));
 sky130_fd_sc_hd__o21ai_1 _44618_ (.A1(_17560_),
    .A2(_17549_),
    .B1(_17649_),
    .Y(_17650_));
 sky130_fd_sc_hd__clkbuf_2 _44619_ (.A(_17650_),
    .X(_17651_));
 sky130_fd_sc_hd__nand2_1 _44620_ (.A(_17547_),
    .B(_17545_),
    .Y(_17653_));
 sky130_fd_sc_hd__o2111ai_4 _44621_ (.A1(_17542_),
    .A2(_17544_),
    .B1(_17647_),
    .C1(_17653_),
    .D1(_17648_),
    .Y(_17654_));
 sky130_fd_sc_hd__a22oi_1 _44622_ (.A1(_17558_),
    .A2(_17556_),
    .B1(_17651_),
    .B2(_17654_),
    .Y(_17655_));
 sky130_fd_sc_hd__nand4_1 _44623_ (.A(_17558_),
    .B(_17556_),
    .C(_17651_),
    .D(_17654_),
    .Y(_17656_));
 sky130_fd_sc_hd__nor2b_1 _44624_ (.A(_17655_),
    .B_N(_17656_),
    .Y(_17657_));
 sky130_fd_sc_hd__clkbuf_1 _44625_ (.A(_17657_),
    .X(_00024_));
 sky130_fd_sc_hd__o21ai_4 _44626_ (.A1(_17485_),
    .A2(_17573_),
    .B1(_17569_),
    .Y(_17658_));
 sky130_fd_sc_hd__xnor2_1 _44627_ (.A(_17523_),
    .B(_17658_),
    .Y(_17659_));
 sky130_fd_sc_hd__mux2_1 _44628_ (.A0(_17579_),
    .A1(_17577_),
    .S(_17505_),
    .X(_17660_));
 sky130_fd_sc_hd__a21oi_2 _44629_ (.A1(_17472_),
    .A2(_17565_),
    .B1(_17568_),
    .Y(_17661_));
 sky130_fd_sc_hd__and4_1 _44630_ (.A(_17472_),
    .B(_16716_),
    .C(_17022_),
    .D(_17568_),
    .X(_17663_));
 sky130_fd_sc_hd__or2_1 _44631_ (.A(_17661_),
    .B(_17663_),
    .X(_17664_));
 sky130_fd_sc_hd__xnor2_1 _44632_ (.A(_17660_),
    .B(_17664_),
    .Y(_17665_));
 sky130_fd_sc_hd__o211ai_2 _44633_ (.A1(_17507_),
    .A2(_17582_),
    .B1(_17665_),
    .C1(_17588_),
    .Y(_17666_));
 sky130_fd_sc_hd__nand2_2 _44634_ (.A(_17659_),
    .B(_17666_),
    .Y(_17667_));
 sky130_fd_sc_hd__a21o_1 _44635_ (.A1(_17583_),
    .A2(_17588_),
    .B1(_17665_),
    .X(_17668_));
 sky130_fd_sc_hd__inv_2 _44636_ (.A(_17668_),
    .Y(_17669_));
 sky130_fd_sc_hd__inv_2 _44637_ (.A(_17511_),
    .Y(_17670_));
 sky130_fd_sc_hd__a21oi_2 _44638_ (.A1(_17670_),
    .A2(_17527_),
    .B1(_17589_),
    .Y(_17671_));
 sky130_fd_sc_hd__a31oi_2 _44639_ (.A1(_17670_),
    .A2(_17527_),
    .A3(_17589_),
    .B1(_17624_),
    .Y(_17672_));
 sky130_fd_sc_hd__a21o_1 _44640_ (.A1(_17668_),
    .A2(_17666_),
    .B1(_17659_),
    .X(_17674_));
 sky130_fd_sc_hd__o221ai_4 _44641_ (.A1(_17667_),
    .A2(_17669_),
    .B1(_17671_),
    .B2(_17672_),
    .C1(_17674_),
    .Y(_17675_));
 sky130_fd_sc_hd__o21ai_1 _44642_ (.A1(_17669_),
    .A2(_17667_),
    .B1(_17674_),
    .Y(_17676_));
 sky130_fd_sc_hd__a31o_1 _44643_ (.A1(_17670_),
    .A2(_17527_),
    .A3(_17589_),
    .B1(_17624_),
    .X(_17677_));
 sky130_fd_sc_hd__nand3_1 _44644_ (.A(_17591_),
    .B(_17676_),
    .C(_17677_),
    .Y(_17678_));
 sky130_fd_sc_hd__nor2_1 _44645_ (.A(_16716_),
    .B(_17592_),
    .Y(_17679_));
 sky130_fd_sc_hd__or2_1 _44646_ (.A(_17312_),
    .B(_17622_),
    .X(_17680_));
 sky130_fd_sc_hd__o31a_1 _44647_ (.A1(_17561_),
    .A2(_17562_),
    .A3(_17679_),
    .B1(_17680_),
    .X(_17681_));
 sky130_fd_sc_hd__a21oi_2 _44648_ (.A1(_17675_),
    .A2(_17678_),
    .B1(_17681_),
    .Y(_17682_));
 sky130_fd_sc_hd__and3_2 _44649_ (.A(_17675_),
    .B(_17678_),
    .C(_17681_),
    .X(_17683_));
 sky130_fd_sc_hd__a211o_1 _44650_ (.A1(_17629_),
    .A2(_17643_),
    .B1(_17682_),
    .C1(_17683_),
    .X(_17685_));
 sky130_fd_sc_hd__o211ai_4 _44651_ (.A1(_17682_),
    .A2(_17683_),
    .B1(_17629_),
    .C1(_17643_),
    .Y(_17686_));
 sky130_fd_sc_hd__o21a_1 _44652_ (.A1(_17561_),
    .A2(_17562_),
    .B1(_17634_),
    .X(_17687_));
 sky130_fd_sc_hd__and3_1 _44653_ (.A(_17685_),
    .B(_17686_),
    .C(_17687_),
    .X(_17688_));
 sky130_fd_sc_hd__a21oi_1 _44654_ (.A1(_17685_),
    .A2(_17686_),
    .B1(_17687_),
    .Y(_17689_));
 sky130_fd_sc_hd__o211a_1 _44655_ (.A1(_17642_),
    .A2(_17643_),
    .B1(_17644_),
    .C1(_17645_),
    .X(_17690_));
 sky130_fd_sc_hd__a21oi_1 _44656_ (.A1(_17563_),
    .A2(_17640_),
    .B1(_17690_),
    .Y(_17691_));
 sky130_fd_sc_hd__o21ai_2 _44657_ (.A1(_17688_),
    .A2(_17689_),
    .B1(_17691_),
    .Y(_17692_));
 sky130_fd_sc_hd__inv_2 _44658_ (.A(_17692_),
    .Y(_17693_));
 sky130_fd_sc_hd__o21ai_1 _44659_ (.A1(_17642_),
    .A2(_17643_),
    .B1(_17644_),
    .Y(_17694_));
 sky130_fd_sc_hd__a21boi_1 _44660_ (.A1(_17694_),
    .A2(_17639_),
    .B1_N(_17563_),
    .Y(_17696_));
 sky130_fd_sc_hd__o2111ai_2 _44661_ (.A1(_17561_),
    .A2(_17562_),
    .B1(_17634_),
    .C1(_17685_),
    .D1(_17686_),
    .Y(_17697_));
 sky130_fd_sc_hd__clkbuf_2 _44662_ (.A(_17633_),
    .X(_17698_));
 sky130_fd_sc_hd__a22o_1 _44663_ (.A1(_17698_),
    .A2(_17634_),
    .B1(_17685_),
    .B2(_17686_),
    .X(_17699_));
 sky130_fd_sc_hd__o211a_1 _44664_ (.A1(_17690_),
    .A2(_17696_),
    .B1(_17697_),
    .C1(_17699_),
    .X(_17700_));
 sky130_fd_sc_hd__o2bb2ai_1 _44665_ (.A1_N(_17651_),
    .A2_N(_17656_),
    .B1(_17693_),
    .B2(_17700_),
    .Y(_17701_));
 sky130_fd_sc_hd__o211ai_2 _44666_ (.A1(_17690_),
    .A2(_17696_),
    .B1(_17697_),
    .C1(_17699_),
    .Y(_17702_));
 sky130_fd_sc_hd__nand4_1 _44667_ (.A(_17651_),
    .B(_17656_),
    .C(_17692_),
    .D(_17702_),
    .Y(_17703_));
 sky130_fd_sc_hd__nand2_1 _44668_ (.A(_17701_),
    .B(_17703_),
    .Y(_00025_));
 sky130_fd_sc_hd__a21boi_1 _44669_ (.A1(_17687_),
    .A2(_17686_),
    .B1_N(_17685_),
    .Y(_17704_));
 sky130_fd_sc_hd__o221a_1 _44670_ (.A1(_17667_),
    .A2(_17669_),
    .B1(_17671_),
    .B2(_17672_),
    .C1(_17674_),
    .X(_17706_));
 sky130_fd_sc_hd__a21oi_1 _44671_ (.A1(_17658_),
    .A2(_17520_),
    .B1(_17633_),
    .Y(_17707_));
 sky130_fd_sc_hd__a21o_1 _44672_ (.A1(_17633_),
    .A2(_17658_),
    .B1(_17707_),
    .X(_17708_));
 sky130_fd_sc_hd__o211ai_4 _44673_ (.A1(_17661_),
    .A2(_17663_),
    .B1(_17505_),
    .C1(_17577_),
    .Y(_17709_));
 sky130_fd_sc_hd__or4_2 _44674_ (.A(_17406_),
    .B(_17505_),
    .C(_17578_),
    .D(_17664_),
    .X(_17710_));
 sky130_fd_sc_hd__clkbuf_2 _44675_ (.A(_17661_),
    .X(_17711_));
 sky130_fd_sc_hd__xor2_1 _44676_ (.A(_17523_),
    .B(_17711_),
    .X(_17712_));
 sky130_fd_sc_hd__a21boi_1 _44677_ (.A1(_17709_),
    .A2(_17710_),
    .B1_N(_17712_),
    .Y(_17713_));
 sky130_fd_sc_hd__and3b_1 _44678_ (.A_N(_17712_),
    .B(_17709_),
    .C(_17710_),
    .X(_17714_));
 sky130_fd_sc_hd__a211oi_1 _44679_ (.A1(_17668_),
    .A2(_17667_),
    .B1(_17713_),
    .C1(_17714_),
    .Y(_17715_));
 sky130_fd_sc_hd__o211ai_1 _44680_ (.A1(_17713_),
    .A2(_17714_),
    .B1(_17668_),
    .C1(_17667_),
    .Y(_17717_));
 sky130_fd_sc_hd__nand2b_1 _44681_ (.A_N(_17715_),
    .B(_17717_),
    .Y(_17718_));
 sky130_fd_sc_hd__xor2_2 _44682_ (.A(_17708_),
    .B(_17718_),
    .X(_17719_));
 sky130_fd_sc_hd__o21ai_2 _44683_ (.A1(_17706_),
    .A2(_17683_),
    .B1(_17719_),
    .Y(_17720_));
 sky130_fd_sc_hd__or3_1 _44684_ (.A(_17706_),
    .B(_17683_),
    .C(_17719_),
    .X(_17721_));
 sky130_fd_sc_hd__nand2_1 _44685_ (.A(_17720_),
    .B(_17721_),
    .Y(_17722_));
 sky130_fd_sc_hd__xnor2_1 _44686_ (.A(_17680_),
    .B(_17722_),
    .Y(_17723_));
 sky130_fd_sc_hd__nand2_1 _44687_ (.A(_17704_),
    .B(_17723_),
    .Y(_17724_));
 sky130_fd_sc_hd__or2_2 _44688_ (.A(_17704_),
    .B(_17723_),
    .X(_17725_));
 sky130_fd_sc_hd__nand2_2 _44689_ (.A(_17724_),
    .B(_17725_),
    .Y(_17726_));
 sky130_fd_sc_hd__nand2_1 _44690_ (.A(_17650_),
    .B(_17654_),
    .Y(_17728_));
 sky130_fd_sc_hd__nand2_1 _44691_ (.A(_17692_),
    .B(_17702_),
    .Y(_17729_));
 sky130_fd_sc_hd__and4bb_1 _44692_ (.A_N(_17728_),
    .B_N(_17729_),
    .C(_17558_),
    .D(_17555_),
    .X(_17730_));
 sky130_fd_sc_hd__nand2_1 _44693_ (.A(_17651_),
    .B(_17702_),
    .Y(_17731_));
 sky130_fd_sc_hd__o21ai_1 _44694_ (.A1(_17340_),
    .A2(_17458_),
    .B1(_17555_),
    .Y(_17732_));
 sky130_fd_sc_hd__nor3_1 _44695_ (.A(_17729_),
    .B(_17553_),
    .C(_17728_),
    .Y(_17733_));
 sky130_fd_sc_hd__a22o_1 _44696_ (.A1(_17692_),
    .A2(_17731_),
    .B1(_17732_),
    .B2(_17733_),
    .X(_17734_));
 sky130_fd_sc_hd__a31oi_4 _44697_ (.A1(_17463_),
    .A2(_17730_),
    .A3(_17459_),
    .B1(_17734_),
    .Y(_17735_));
 sky130_fd_sc_hd__xor2_1 _44698_ (.A(_17726_),
    .B(_17735_),
    .X(_00026_));
 sky130_fd_sc_hd__o21bai_2 _44699_ (.A1(_17706_),
    .A2(_17719_),
    .B1_N(_17680_),
    .Y(_17736_));
 sky130_fd_sc_hd__a21oi_2 _44700_ (.A1(_17569_),
    .A2(_17576_),
    .B1(_17312_),
    .Y(_17738_));
 sky130_fd_sc_hd__a211o_1 _44701_ (.A1(_17520_),
    .A2(_17711_),
    .B1(_17562_),
    .C1(_17561_),
    .X(_17739_));
 sky130_fd_sc_hd__a21bo_1 _44702_ (.A1(_17698_),
    .A2(_17711_),
    .B1_N(_17739_),
    .X(_17740_));
 sky130_fd_sc_hd__mux2_1 _44703_ (.A0(_17710_),
    .A1(_17709_),
    .S(_17712_),
    .X(_17741_));
 sky130_fd_sc_hd__xnor2_1 _44704_ (.A(_17740_),
    .B(_17741_),
    .Y(_17742_));
 sky130_fd_sc_hd__nor3b_1 _44705_ (.A(_17738_),
    .B(_17707_),
    .C_N(_17717_),
    .Y(_17743_));
 sky130_fd_sc_hd__nor3_1 _44706_ (.A(_17715_),
    .B(_17742_),
    .C(_17743_),
    .Y(_17744_));
 sky130_fd_sc_hd__o21a_1 _44707_ (.A1(_17715_),
    .A2(_17743_),
    .B1(_17742_),
    .X(_17745_));
 sky130_fd_sc_hd__nor2_1 _44708_ (.A(_17744_),
    .B(_17745_),
    .Y(_17746_));
 sky130_fd_sc_hd__xnor2_2 _44709_ (.A(_17738_),
    .B(_17746_),
    .Y(_17747_));
 sky130_fd_sc_hd__a21o_1 _44710_ (.A1(_17720_),
    .A2(_17736_),
    .B1(_17747_),
    .X(_17749_));
 sky130_fd_sc_hd__nand3_4 _44711_ (.A(_17720_),
    .B(_17736_),
    .C(_17747_),
    .Y(_17750_));
 sky130_fd_sc_hd__nand2_1 _44712_ (.A(_17749_),
    .B(_17750_),
    .Y(_17751_));
 sky130_fd_sc_hd__o21ai_1 _44713_ (.A1(_17726_),
    .A2(_17735_),
    .B1(_17725_),
    .Y(_17752_));
 sky130_fd_sc_hd__xnor2_1 _44714_ (.A(_17751_),
    .B(_17752_),
    .Y(_00027_));
 sky130_fd_sc_hd__o211ai_4 _44715_ (.A1(_17726_),
    .A2(_17735_),
    .B1(_17749_),
    .C1(_17725_),
    .Y(_17753_));
 sky130_fd_sc_hd__nor4_2 _44716_ (.A(_17520_),
    .B(_17698_),
    .C(_17711_),
    .D(_17709_),
    .Y(_17754_));
 sky130_fd_sc_hd__a31o_4 _44717_ (.A1(_17746_),
    .A2(_17658_),
    .A3(_17698_),
    .B1(_17745_),
    .X(_17755_));
 sky130_fd_sc_hd__nor2_1 _44718_ (.A(net58),
    .B(_17755_),
    .Y(_17756_));
 sky130_fd_sc_hd__and3_1 _44719_ (.A(_17698_),
    .B(_17709_),
    .C(_17711_),
    .X(_17757_));
 sky130_fd_sc_hd__o21ba_4 _44720_ (.A1(_17710_),
    .A2(_17740_),
    .B1_N(_17757_),
    .X(_17759_));
 sky130_fd_sc_hd__inv_2 _44721_ (.A(_17759_),
    .Y(_17760_));
 sky130_fd_sc_hd__o2bb2ai_1 _44722_ (.A1_N(_17750_),
    .A2_N(_17753_),
    .B1(_17756_),
    .B2(_17760_),
    .Y(_17761_));
 sky130_fd_sc_hd__o2111ai_1 _44723_ (.A1(_17755_),
    .A2(net58),
    .B1(_17759_),
    .C1(_17750_),
    .D1(_17753_),
    .Y(_17762_));
 sky130_fd_sc_hd__nand2_1 _44724_ (.A(_17761_),
    .B(_17762_),
    .Y(_00028_));
 sky130_fd_sc_hd__buf_1 _44725_ (.A(_17750_),
    .X(_17763_));
 sky130_fd_sc_hd__buf_6 _44726_ (.A(_17753_),
    .X(_17764_));
 sky130_fd_sc_hd__o2bb2a_1 _44727_ (.A1_N(_17763_),
    .A2_N(_17764_),
    .B1(_17756_),
    .B2(_17760_),
    .X(_00029_));
 sky130_fd_sc_hd__o2bb2a_1 _44728_ (.A1_N(_17763_),
    .A2_N(_17764_),
    .B1(_17756_),
    .B2(_17760_),
    .X(_00030_));
 sky130_fd_sc_hd__o2bb2a_1 _44729_ (.A1_N(_17763_),
    .A2_N(_17764_),
    .B1(_17756_),
    .B2(_17760_),
    .X(_00031_));
 sky130_fd_sc_hd__a221oi_1 _44730_ (.A1(_17759_),
    .A2(_17755_),
    .B1(_17764_),
    .B2(_17763_),
    .C1(net58),
    .Y(_00032_));
 sky130_fd_sc_hd__a221oi_1 _44731_ (.A1(_17759_),
    .A2(_17755_),
    .B1(_17764_),
    .B2(_17763_),
    .C1(net58),
    .Y(_00033_));
 sky130_fd_sc_hd__a221oi_1 _44732_ (.A1(_17759_),
    .A2(_17755_),
    .B1(_17753_),
    .B2(_17750_),
    .C1(net58),
    .Y(_00034_));
 sky130_fd_sc_hd__and2_1 _44733_ (.A(_11207_),
    .B(_11218_),
    .X(_17766_));
 sky130_fd_sc_hd__nor2_1 _44734_ (.A(_17892_),
    .B(_17766_),
    .Y(_00003_));
 sky130_fd_sc_hd__inv_2 _44735_ (.A(net378),
    .Y(_22139_));
 sky130_fd_sc_hd__buf_2 _44736_ (.A(_22139_),
    .X(_22150_));
 sky130_fd_sc_hd__buf_1 _44737_ (.A(\delay_line[20][0] ),
    .X(_22161_));
 sky130_fd_sc_hd__buf_2 _44738_ (.A(_22161_),
    .X(_22172_));
 sky130_fd_sc_hd__buf_1 _44739_ (.A(_22172_),
    .X(_22183_));
 sky130_fd_sc_hd__clkbuf_2 _44740_ (.A(_22183_),
    .X(_22194_));
 sky130_fd_sc_hd__clkbuf_4 _44741_ (.A(_22194_),
    .X(_22205_));
 sky130_fd_sc_hd__buf_1 _44742_ (.A(\delay_line[31][0] ),
    .X(_22215_));
 sky130_fd_sc_hd__inv_2 _44743_ (.A(_22215_),
    .Y(_22226_));
 sky130_fd_sc_hd__clkbuf_4 _44744_ (.A(_22226_),
    .X(_22237_));
 sky130_fd_sc_hd__buf_1 _44745_ (.A(\delay_line[28][0] ),
    .X(_22248_));
 sky130_fd_sc_hd__clkbuf_2 _44746_ (.A(_22248_),
    .X(_22259_));
 sky130_fd_sc_hd__buf_4 _44747_ (.A(_22259_),
    .X(_22270_));
 sky130_fd_sc_hd__buf_1 _44748_ (.A(\delay_line[30][0] ),
    .X(_22281_));
 sky130_fd_sc_hd__buf_1 _44749_ (.A(_22281_),
    .X(_22292_));
 sky130_fd_sc_hd__clkbuf_4 _44750_ (.A(_22292_),
    .X(_22303_));
 sky130_fd_sc_hd__nor2_1 _44751_ (.A(_22270_),
    .B(_22303_),
    .Y(_22314_));
 sky130_fd_sc_hd__and2_1 _44752_ (.A(_22270_),
    .B(_22303_),
    .X(_22325_));
 sky130_fd_sc_hd__or3_1 _44753_ (.A(_22237_),
    .B(_22314_),
    .C(_22325_),
    .X(_22336_));
 sky130_fd_sc_hd__o21ai_1 _44754_ (.A1(_22314_),
    .A2(_22325_),
    .B1(_22237_),
    .Y(_22347_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44755_ (.A(\delay_line[25][0] ),
    .X(_22358_));
 sky130_fd_sc_hd__buf_1 _44756_ (.A(_22358_),
    .X(_22369_));
 sky130_fd_sc_hd__clkbuf_4 _44757_ (.A(_22369_),
    .X(_22380_));
 sky130_fd_sc_hd__buf_1 _44758_ (.A(\delay_line[15][0] ),
    .X(_22391_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44759_ (.A(_22391_),
    .X(_22402_));
 sky130_fd_sc_hd__clkbuf_2 _44760_ (.A(_22402_),
    .X(_22413_));
 sky130_fd_sc_hd__buf_4 _44761_ (.A(_22413_),
    .X(_22424_));
 sky130_fd_sc_hd__and2_1 _44762_ (.A(_22380_),
    .B(_22424_),
    .X(_22435_));
 sky130_fd_sc_hd__nor2_1 _44763_ (.A(_22380_),
    .B(_22424_),
    .Y(_22446_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44764_ (.A(\delay_line[27][0] ),
    .X(_22457_));
 sky130_fd_sc_hd__buf_4 _44765_ (.A(_22457_),
    .X(_22468_));
 sky130_fd_sc_hd__or3b_2 _44766_ (.A(_22435_),
    .B(_22446_),
    .C_N(_22468_),
    .X(_22479_));
 sky130_fd_sc_hd__o21bai_2 _44767_ (.A1(_22435_),
    .A2(_22446_),
    .B1_N(_22468_),
    .Y(_22490_));
 sky130_fd_sc_hd__and4_1 _44768_ (.A(_22336_),
    .B(_22347_),
    .C(_22479_),
    .D(_22490_),
    .X(_22501_));
 sky130_fd_sc_hd__a22oi_2 _44769_ (.A1(_22336_),
    .A2(_22347_),
    .B1(_22479_),
    .B2(_22490_),
    .Y(_22512_));
 sky130_fd_sc_hd__clkbuf_2 _44770_ (.A(net315),
    .X(_22523_));
 sky130_fd_sc_hd__clkbuf_2 _44771_ (.A(_22523_),
    .X(_22534_));
 sky130_fd_sc_hd__buf_1 _44772_ (.A(_22534_),
    .X(_22545_));
 sky130_fd_sc_hd__buf_1 _44773_ (.A(\delay_line[32][0] ),
    .X(_22556_));
 sky130_fd_sc_hd__buf_1 _44774_ (.A(_22556_),
    .X(_22567_));
 sky130_fd_sc_hd__buf_1 _44775_ (.A(_22567_),
    .X(_22578_));
 sky130_fd_sc_hd__nor2_1 _44776_ (.A(_22545_),
    .B(_22578_),
    .Y(_22589_));
 sky130_fd_sc_hd__and2_1 _44777_ (.A(_22545_),
    .B(_22578_),
    .X(_22600_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44778_ (.A(\delay_line[34][0] ),
    .X(_22611_));
 sky130_fd_sc_hd__buf_1 _44779_ (.A(_22611_),
    .X(_22622_));
 sky130_fd_sc_hd__or3b_1 _44780_ (.A(_22589_),
    .B(_22600_),
    .C_N(_22622_),
    .X(_22633_));
 sky130_fd_sc_hd__o21bai_1 _44781_ (.A1(_22589_),
    .A2(_22600_),
    .B1_N(_22622_),
    .Y(_22644_));
 sky130_fd_sc_hd__a2bb2oi_2 _44782_ (.A1_N(_22501_),
    .A2_N(_22512_),
    .B1(_22633_),
    .B2(_22644_),
    .Y(_22655_));
 sky130_fd_sc_hd__and4bb_2 _44783_ (.A_N(_22501_),
    .B_N(_22512_),
    .C(_22633_),
    .D(_22644_),
    .X(_22666_));
 sky130_fd_sc_hd__clkbuf_4 _44784_ (.A(net302),
    .X(_22677_));
 sky130_fd_sc_hd__clkbuf_4 _44785_ (.A(\delay_line[37][0] ),
    .X(_22688_));
 sky130_fd_sc_hd__nor2_1 _44786_ (.A(_22677_),
    .B(_22688_),
    .Y(_22699_));
 sky130_fd_sc_hd__and2_1 _44787_ (.A(_22677_),
    .B(_22688_),
    .X(_22710_));
 sky130_fd_sc_hd__buf_2 _44788_ (.A(\delay_line[38][0] ),
    .X(_22721_));
 sky130_fd_sc_hd__or3b_1 _44789_ (.A(_22699_),
    .B(_22710_),
    .C_N(_22721_),
    .X(_22732_));
 sky130_fd_sc_hd__o21bai_2 _44790_ (.A1(_22699_),
    .A2(_22710_),
    .B1_N(_22721_),
    .Y(_22743_));
 sky130_fd_sc_hd__buf_1 _44791_ (.A(\delay_line[39][0] ),
    .X(_22754_));
 sky130_fd_sc_hd__buf_1 _44792_ (.A(_22754_),
    .X(_22765_));
 sky130_fd_sc_hd__buf_1 _44793_ (.A(\delay_line[40][0] ),
    .X(_22776_));
 sky130_fd_sc_hd__buf_1 _44794_ (.A(_22776_),
    .X(_22787_));
 sky130_fd_sc_hd__nor2_1 _44795_ (.A(_22765_),
    .B(_22787_),
    .Y(_22798_));
 sky130_fd_sc_hd__and2_1 _44796_ (.A(_22765_),
    .B(_22787_),
    .X(_22809_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44797_ (.A(\delay_line[3][0] ),
    .X(_22820_));
 sky130_fd_sc_hd__clkbuf_2 _44798_ (.A(\delay_line[5][0] ),
    .X(_22831_));
 sky130_fd_sc_hd__clkbuf_2 _44799_ (.A(_22831_),
    .X(_22842_));
 sky130_fd_sc_hd__nor2_1 _44800_ (.A(_22820_),
    .B(_22842_),
    .Y(_22853_));
 sky130_fd_sc_hd__and2_1 _44801_ (.A(_22820_),
    .B(_22842_),
    .X(_22864_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44802_ (.A(\delay_line[2][0] ),
    .X(_22875_));
 sky130_fd_sc_hd__or3b_2 _44803_ (.A(_22853_),
    .B(_22864_),
    .C_N(_22875_),
    .X(_22886_));
 sky130_fd_sc_hd__buf_1 _44804_ (.A(\delay_line[6][0] ),
    .X(_22897_));
 sky130_fd_sc_hd__clkbuf_2 _44805_ (.A(_22897_),
    .X(_22908_));
 sky130_fd_sc_hd__buf_2 _44806_ (.A(_22908_),
    .X(_22919_));
 sky130_fd_sc_hd__o21bai_1 _44807_ (.A1(_22853_),
    .A2(_22864_),
    .B1_N(_22875_),
    .Y(_22930_));
 sky130_fd_sc_hd__and3_1 _44808_ (.A(_22886_),
    .B(_22919_),
    .C(_22930_),
    .X(_22941_));
 sky130_fd_sc_hd__a21oi_1 _44809_ (.A1(_22930_),
    .A2(_22886_),
    .B1(_22919_),
    .Y(_22952_));
 sky130_fd_sc_hd__inv_2 _44810_ (.A(\delay_line[7][0] ),
    .Y(_22963_));
 sky130_fd_sc_hd__clkbuf_4 _44811_ (.A(_22963_),
    .X(_22974_));
 sky130_fd_sc_hd__buf_1 _44812_ (.A(\delay_line[8][0] ),
    .X(_22985_));
 sky130_fd_sc_hd__inv_2 _44813_ (.A(_22985_),
    .Y(_22996_));
 sky130_fd_sc_hd__nor2_2 _44814_ (.A(_22974_),
    .B(_22996_),
    .Y(_23007_));
 sky130_fd_sc_hd__clkbuf_2 _44815_ (.A(\delay_line[7][0] ),
    .X(_23018_));
 sky130_fd_sc_hd__clkbuf_2 _44816_ (.A(_23018_),
    .X(_23029_));
 sky130_fd_sc_hd__buf_2 _44817_ (.A(_22985_),
    .X(_23040_));
 sky130_fd_sc_hd__buf_2 _44818_ (.A(_23040_),
    .X(_23051_));
 sky130_fd_sc_hd__nor2_1 _44819_ (.A(_23029_),
    .B(_23051_),
    .Y(_23062_));
 sky130_fd_sc_hd__buf_2 _44820_ (.A(\delay_line[9][0] ),
    .X(_23073_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44821_ (.A(_23073_),
    .X(_23084_));
 sky130_fd_sc_hd__buf_2 _44822_ (.A(_23084_),
    .X(_23095_));
 sky130_fd_sc_hd__clkbuf_2 _44823_ (.A(net415),
    .X(_23106_));
 sky130_fd_sc_hd__buf_2 _44824_ (.A(_23106_),
    .X(_23117_));
 sky130_fd_sc_hd__or2_1 _44825_ (.A(_23095_),
    .B(_23117_),
    .X(_23128_));
 sky130_fd_sc_hd__nand2_1 _44826_ (.A(_23095_),
    .B(_23117_),
    .Y(_23139_));
 sky130_fd_sc_hd__buf_1 _44827_ (.A(\delay_line[0][0] ),
    .X(_23150_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44828_ (.A(_23150_),
    .X(_23161_));
 sky130_fd_sc_hd__clkbuf_2 _44829_ (.A(_23161_),
    .X(_23172_));
 sky130_fd_sc_hd__nor2_1 _44830_ (.A(net398),
    .B(_23172_),
    .Y(_23183_));
 sky130_fd_sc_hd__inv_2 _44831_ (.A(net398),
    .Y(_23194_));
 sky130_fd_sc_hd__inv_2 _44832_ (.A(\delay_line[0][0] ),
    .Y(_23205_));
 sky130_fd_sc_hd__nor2_1 _44833_ (.A(_23194_),
    .B(_23205_),
    .Y(_23216_));
 sky130_fd_sc_hd__buf_1 _44834_ (.A(\delay_line[12][0] ),
    .X(_23227_));
 sky130_fd_sc_hd__buf_1 _44835_ (.A(_23227_),
    .X(_23238_));
 sky130_fd_sc_hd__or3b_2 _44836_ (.A(_23183_),
    .B(_23216_),
    .C_N(_23238_),
    .X(_23249_));
 sky130_fd_sc_hd__clkbuf_2 _44837_ (.A(_23238_),
    .X(_23260_));
 sky130_fd_sc_hd__o21bai_2 _44838_ (.A1(_23183_),
    .A2(_23216_),
    .B1_N(_23260_),
    .Y(_23271_));
 sky130_fd_sc_hd__a22oi_2 _44839_ (.A1(_23128_),
    .A2(_23139_),
    .B1(_23249_),
    .B2(_23271_),
    .Y(_23282_));
 sky130_fd_sc_hd__and4_1 _44840_ (.A(_23128_),
    .B(_23139_),
    .C(_23249_),
    .D(_23271_),
    .X(_23293_));
 sky130_fd_sc_hd__nor4_1 _44841_ (.A(_23007_),
    .B(_23062_),
    .C(_23282_),
    .D(_23293_),
    .Y(_23304_));
 sky130_fd_sc_hd__o22ai_1 _44842_ (.A1(_23007_),
    .A2(_23062_),
    .B1(_23282_),
    .B2(_23293_),
    .Y(_23315_));
 sky130_fd_sc_hd__inv_2 _44843_ (.A(_23315_),
    .Y(_23326_));
 sky130_fd_sc_hd__or4_2 _44844_ (.A(_22941_),
    .B(_22952_),
    .C(net185),
    .D(_23326_),
    .X(_23337_));
 sky130_fd_sc_hd__o22a_1 _44845_ (.A1(_22941_),
    .A2(_22952_),
    .B1(net185),
    .B2(_23326_),
    .X(_23348_));
 sky130_fd_sc_hd__inv_2 _44846_ (.A(_23348_),
    .Y(_23359_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44847_ (.A(\delay_line[1][0] ),
    .X(_23370_));
 sky130_fd_sc_hd__and3_2 _44848_ (.A(_23337_),
    .B(_23359_),
    .C(_23370_),
    .X(_23381_));
 sky130_fd_sc_hd__a21o_1 _44849_ (.A1(_23337_),
    .A2(_23359_),
    .B1(_23370_),
    .X(_23392_));
 sky130_fd_sc_hd__or4b_4 _44850_ (.A(_22798_),
    .B(_22809_),
    .C(_23381_),
    .D_N(_23392_),
    .X(_23403_));
 sky130_fd_sc_hd__inv_2 _44851_ (.A(\delay_line[1][0] ),
    .Y(_23414_));
 sky130_fd_sc_hd__or3b_4 _44852_ (.A(_23348_),
    .B(_23414_),
    .C_N(_23337_),
    .X(_23425_));
 sky130_fd_sc_hd__a2bb2o_2 _44853_ (.A1_N(_22798_),
    .A2_N(_22809_),
    .B1(_23425_),
    .B2(_23392_),
    .X(_23436_));
 sky130_fd_sc_hd__and4_2 _44854_ (.A(_22732_),
    .B(_22743_),
    .C(_23403_),
    .D(_23436_),
    .X(_23447_));
 sky130_fd_sc_hd__a22oi_4 _44855_ (.A1(_22732_),
    .A2(_22743_),
    .B1(_23403_),
    .B2(_23436_),
    .Y(_23458_));
 sky130_fd_sc_hd__or4_2 _44856_ (.A(_22655_),
    .B(_22666_),
    .C(_23447_),
    .D(_23458_),
    .X(_23469_));
 sky130_fd_sc_hd__buf_1 _44857_ (.A(_23469_),
    .X(_23480_));
 sky130_fd_sc_hd__o22ai_4 _44858_ (.A1(_22655_),
    .A2(_22666_),
    .B1(_23447_),
    .B2(_23458_),
    .Y(_23491_));
 sky130_fd_sc_hd__buf_1 _44859_ (.A(\delay_line[23][0] ),
    .X(_23502_));
 sky130_fd_sc_hd__buf_2 _44860_ (.A(_23502_),
    .X(_23513_));
 sky130_fd_sc_hd__buf_1 _44861_ (.A(_23513_),
    .X(_23524_));
 sky130_fd_sc_hd__and3_1 _44862_ (.A(_23480_),
    .B(_23491_),
    .C(_23524_),
    .X(_23535_));
 sky130_fd_sc_hd__a21oi_1 _44863_ (.A1(_23480_),
    .A2(_23491_),
    .B1(_23524_),
    .Y(_23546_));
 sky130_fd_sc_hd__nor2_1 _44864_ (.A(_23535_),
    .B(_23546_),
    .Y(_23557_));
 sky130_fd_sc_hd__xnor2_2 _44865_ (.A(_22205_),
    .B(_23557_),
    .Y(_23568_));
 sky130_fd_sc_hd__xor2_2 _44866_ (.A(_22150_),
    .B(_23568_),
    .X(_00000_));
 sky130_fd_sc_hd__or2_1 _44867_ (.A(_22150_),
    .B(_23568_),
    .X(_23589_));
 sky130_fd_sc_hd__clkbuf_2 _44868_ (.A(net368),
    .X(_23600_));
 sky130_fd_sc_hd__clkbuf_2 _44869_ (.A(_23600_),
    .X(_23611_));
 sky130_fd_sc_hd__clkbuf_2 _44870_ (.A(_23611_),
    .X(_23622_));
 sky130_fd_sc_hd__and2_1 _44871_ (.A(_23513_),
    .B(_23622_),
    .X(_23633_));
 sky130_fd_sc_hd__nor2_1 _44872_ (.A(_23524_),
    .B(_23622_),
    .Y(_23644_));
 sky130_fd_sc_hd__nor3_1 _44873_ (.A(_22237_),
    .B(_22314_),
    .C(_22325_),
    .Y(_23655_));
 sky130_fd_sc_hd__buf_1 _44874_ (.A(\delay_line[22][0] ),
    .X(_23666_));
 sky130_fd_sc_hd__buf_2 _44875_ (.A(_23666_),
    .X(_23676_));
 sky130_fd_sc_hd__clkbuf_2 _44876_ (.A(net346),
    .X(_23687_));
 sky130_fd_sc_hd__buf_2 _44877_ (.A(_23687_),
    .X(_23698_));
 sky130_fd_sc_hd__or2_1 _44878_ (.A(_23676_),
    .B(_23698_),
    .X(_23709_));
 sky130_fd_sc_hd__nand2_2 _44879_ (.A(_23676_),
    .B(_23698_),
    .Y(_23720_));
 sky130_fd_sc_hd__buf_1 _44880_ (.A(\delay_line[25][1] ),
    .X(_23731_));
 sky130_fd_sc_hd__buf_4 _44881_ (.A(_23731_),
    .X(_23742_));
 sky130_fd_sc_hd__nand3_1 _44882_ (.A(_23709_),
    .B(_23720_),
    .C(_23742_),
    .Y(_23753_));
 sky130_fd_sc_hd__a21o_1 _44883_ (.A1(_23709_),
    .A2(_23720_),
    .B1(_23742_),
    .X(_23764_));
 sky130_fd_sc_hd__o211a_1 _44884_ (.A1(_22325_),
    .A2(_23655_),
    .B1(_23753_),
    .C1(_23764_),
    .X(_23775_));
 sky130_fd_sc_hd__clkbuf_2 _44885_ (.A(_23753_),
    .X(_23786_));
 sky130_fd_sc_hd__a221oi_2 _44886_ (.A1(_22270_),
    .A2(_22303_),
    .B1(_23786_),
    .B2(_23764_),
    .C1(_23655_),
    .Y(_23797_));
 sky130_fd_sc_hd__nand2_1 _44887_ (.A(_22545_),
    .B(_22578_),
    .Y(_23808_));
 sky130_fd_sc_hd__o21ai_1 _44888_ (.A1(_22545_),
    .A2(_22578_),
    .B1(_22622_),
    .Y(_23819_));
 sky130_fd_sc_hd__o211ai_2 _44889_ (.A1(_23775_),
    .A2(_23797_),
    .B1(_23808_),
    .C1(_23819_),
    .Y(_23830_));
 sky130_fd_sc_hd__a211o_1 _44890_ (.A1(_23808_),
    .A2(_23819_),
    .B1(_23775_),
    .C1(_23797_),
    .X(_23841_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44891_ (.A(\delay_line[18][0] ),
    .X(_23852_));
 sky130_fd_sc_hd__clkbuf_4 _44892_ (.A(_23852_),
    .X(_23863_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44893_ (.A(\delay_line[19][0] ),
    .X(_23874_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44894_ (.A(_23874_),
    .X(_23885_));
 sky130_fd_sc_hd__buf_1 _44895_ (.A(_23885_),
    .X(_23896_));
 sky130_fd_sc_hd__buf_4 _44896_ (.A(_23896_),
    .X(_23907_));
 sky130_fd_sc_hd__nor2_1 _44897_ (.A(_23863_),
    .B(_23907_),
    .Y(_23918_));
 sky130_fd_sc_hd__inv_2 _44898_ (.A(\delay_line[18][0] ),
    .Y(_23929_));
 sky130_fd_sc_hd__clkbuf_2 _44899_ (.A(_23929_),
    .X(_23940_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44900_ (.A(_23940_),
    .X(_23951_));
 sky130_fd_sc_hd__inv_2 _44901_ (.A(_23885_),
    .Y(_23962_));
 sky130_fd_sc_hd__nor2_2 _44902_ (.A(_23951_),
    .B(_23962_),
    .Y(_23973_));
 sky130_fd_sc_hd__buf_1 _44903_ (.A(\delay_line[21][0] ),
    .X(_23984_));
 sky130_fd_sc_hd__clkbuf_2 _44904_ (.A(_23984_),
    .X(_23995_));
 sky130_fd_sc_hd__clkbuf_2 _44905_ (.A(_23995_),
    .X(_24006_));
 sky130_fd_sc_hd__buf_2 _44906_ (.A(_24006_),
    .X(_24017_));
 sky130_fd_sc_hd__nor3b_2 _44907_ (.A(_23918_),
    .B(_23973_),
    .C_N(_24017_),
    .Y(_24028_));
 sky130_fd_sc_hd__o21ba_1 _44908_ (.A1(_23918_),
    .A2(_23973_),
    .B1_N(_24017_),
    .X(_24039_));
 sky130_fd_sc_hd__a21bo_1 _44909_ (.A1(_22380_),
    .A2(_22424_),
    .B1_N(_22479_),
    .X(_24050_));
 sky130_fd_sc_hd__clkbuf_2 _44910_ (.A(net394),
    .X(_24061_));
 sky130_fd_sc_hd__buf_2 _44911_ (.A(_24061_),
    .X(_24072_));
 sky130_fd_sc_hd__buf_1 _44912_ (.A(\delay_line[15][1] ),
    .X(_24083_));
 sky130_fd_sc_hd__buf_2 _44913_ (.A(_24083_),
    .X(_24094_));
 sky130_fd_sc_hd__or2_2 _44914_ (.A(_24072_),
    .B(_24094_),
    .X(_24105_));
 sky130_fd_sc_hd__nand2_8 _44915_ (.A(_24072_),
    .B(_24094_),
    .Y(_24116_));
 sky130_fd_sc_hd__buf_2 _44916_ (.A(\delay_line[16][0] ),
    .X(_24127_));
 sky130_fd_sc_hd__buf_2 _44917_ (.A(_24127_),
    .X(_24138_));
 sky130_fd_sc_hd__a21o_2 _44918_ (.A1(_24105_),
    .A2(_24116_),
    .B1(_24138_),
    .X(_24149_));
 sky130_fd_sc_hd__nand3_4 _44919_ (.A(_24105_),
    .B(_24116_),
    .C(_24138_),
    .Y(_24160_));
 sky130_fd_sc_hd__nand3_2 _44920_ (.A(_24050_),
    .B(_24149_),
    .C(_24160_),
    .Y(_24171_));
 sky130_fd_sc_hd__a21o_1 _44921_ (.A1(_24149_),
    .A2(_24160_),
    .B1(_24050_),
    .X(_24182_));
 sky130_fd_sc_hd__or4bb_2 _44922_ (.A(_24028_),
    .B(_24039_),
    .C_N(_24171_),
    .D_N(_24182_),
    .X(_24193_));
 sky130_fd_sc_hd__a2bb2o_1 _44923_ (.A1_N(_24028_),
    .A2_N(_24039_),
    .B1(_24171_),
    .B2(_24182_),
    .X(_24204_));
 sky130_fd_sc_hd__nand3_1 _44924_ (.A(_24193_),
    .B(_24204_),
    .C(_22501_),
    .Y(_24215_));
 sky130_fd_sc_hd__a21o_1 _44925_ (.A1(_24193_),
    .A2(_24204_),
    .B1(_22501_),
    .X(_24226_));
 sky130_fd_sc_hd__and4_1 _44926_ (.A(_23830_),
    .B(_23841_),
    .C(_24215_),
    .D(_24226_),
    .X(_24237_));
 sky130_fd_sc_hd__a22oi_1 _44927_ (.A1(_23830_),
    .A2(_23841_),
    .B1(_24215_),
    .B2(_24226_),
    .Y(_24248_));
 sky130_fd_sc_hd__or3b_1 _44928_ (.A(_24237_),
    .B(_24248_),
    .C_N(_22666_),
    .X(_24259_));
 sky130_fd_sc_hd__o21bai_1 _44929_ (.A1(_24237_),
    .A2(_24248_),
    .B1_N(_22666_),
    .Y(_24270_));
 sky130_fd_sc_hd__nand2_1 _44930_ (.A(_24259_),
    .B(_24270_),
    .Y(_24281_));
 sky130_fd_sc_hd__nor3b_2 _44931_ (.A(_22699_),
    .B(_22710_),
    .C_N(_22721_),
    .Y(_24292_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44932_ (.A(\delay_line[27][1] ),
    .X(_24303_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44933_ (.A(\delay_line[26][0] ),
    .X(_24314_));
 sky130_fd_sc_hd__nor2_1 _44934_ (.A(_24303_),
    .B(_24314_),
    .Y(_24325_));
 sky130_fd_sc_hd__inv_2 _44935_ (.A(_24303_),
    .Y(_24336_));
 sky130_fd_sc_hd__inv_2 _44936_ (.A(\delay_line[26][0] ),
    .Y(_24347_));
 sky130_fd_sc_hd__nor2_1 _44937_ (.A(_24336_),
    .B(_24347_),
    .Y(_24358_));
 sky130_fd_sc_hd__buf_1 _44938_ (.A(\delay_line[28][1] ),
    .X(_24369_));
 sky130_fd_sc_hd__buf_2 _44939_ (.A(_24369_),
    .X(_24380_));
 sky130_fd_sc_hd__nor2_1 _44940_ (.A(_22270_),
    .B(_24380_),
    .Y(_24391_));
 sky130_fd_sc_hd__and2_1 _44941_ (.A(_22259_),
    .B(_24380_),
    .X(_24402_));
 sky130_fd_sc_hd__or4_4 _44942_ (.A(_24325_),
    .B(_24358_),
    .C(_24391_),
    .D(_24402_),
    .X(_24413_));
 sky130_fd_sc_hd__o22ai_2 _44943_ (.A1(_24325_),
    .A2(_24358_),
    .B1(_24391_),
    .B2(_24402_),
    .Y(_24424_));
 sky130_fd_sc_hd__o211a_2 _44944_ (.A1(_22710_),
    .A2(_24292_),
    .B1(_24413_),
    .C1(net242),
    .X(_24435_));
 sky130_fd_sc_hd__a221oi_4 _44945_ (.A1(_22677_),
    .A2(_22688_),
    .B1(_24413_),
    .B2(net242),
    .C1(_24292_),
    .Y(_24446_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _44946_ (.A(\delay_line[32][1] ),
    .X(_24457_));
 sky130_fd_sc_hd__clkbuf_2 _44947_ (.A(_24457_),
    .X(_24468_));
 sky130_fd_sc_hd__buf_1 _44948_ (.A(_24468_),
    .X(_24479_));
 sky130_fd_sc_hd__nor2_1 _44949_ (.A(_22578_),
    .B(_24479_),
    .Y(_24490_));
 sky130_fd_sc_hd__inv_2 _44950_ (.A(\delay_line[32][0] ),
    .Y(_24501_));
 sky130_fd_sc_hd__clkbuf_2 _44951_ (.A(_24501_),
    .X(_24512_));
 sky130_fd_sc_hd__inv_2 _44952_ (.A(\delay_line[32][1] ),
    .Y(_24523_));
 sky130_fd_sc_hd__buf_1 _44953_ (.A(_24523_),
    .X(_24534_));
 sky130_fd_sc_hd__clkbuf_2 _44954_ (.A(_24534_),
    .X(_24545_));
 sky130_fd_sc_hd__nor2_1 _44955_ (.A(_24512_),
    .B(_24545_),
    .Y(_24556_));
 sky130_fd_sc_hd__buf_1 _44956_ (.A(_22215_),
    .X(_24567_));
 sky130_fd_sc_hd__clkbuf_2 _44957_ (.A(\delay_line[31][1] ),
    .X(_24578_));
 sky130_fd_sc_hd__buf_1 _44958_ (.A(_24578_),
    .X(_24589_));
 sky130_fd_sc_hd__or2_1 _44959_ (.A(_24567_),
    .B(_24589_),
    .X(_24600_));
 sky130_fd_sc_hd__buf_1 _44960_ (.A(net320),
    .X(_24611_));
 sky130_fd_sc_hd__buf_2 _44961_ (.A(_24611_),
    .X(_24622_));
 sky130_fd_sc_hd__nand2_2 _44962_ (.A(\delay_line[31][0] ),
    .B(_24578_),
    .Y(_24633_));
 sky130_fd_sc_hd__nand3_4 _44963_ (.A(_24600_),
    .B(_24622_),
    .C(_24633_),
    .Y(_24644_));
 sky130_fd_sc_hd__a21o_2 _44964_ (.A1(_24633_),
    .A2(_24600_),
    .B1(_24622_),
    .X(_24655_));
 sky130_fd_sc_hd__a2bb2oi_1 _44965_ (.A1_N(_24490_),
    .A2_N(_24556_),
    .B1(_24644_),
    .B2(_24655_),
    .Y(_24666_));
 sky130_fd_sc_hd__or4bb_2 _44966_ (.A(_24490_),
    .B(_24556_),
    .C_N(_24644_),
    .D_N(_24655_),
    .X(_24677_));
 sky130_fd_sc_hd__inv_2 _44967_ (.A(_24677_),
    .Y(_24688_));
 sky130_fd_sc_hd__nor4_1 _44968_ (.A(_24435_),
    .B(_24446_),
    .C(_24666_),
    .D(_24688_),
    .Y(_24699_));
 sky130_fd_sc_hd__o22a_1 _44969_ (.A1(_24435_),
    .A2(_24446_),
    .B1(_24666_),
    .B2(_24688_),
    .X(_24710_));
 sky130_fd_sc_hd__nor3b_1 _44970_ (.A(_24699_),
    .B(_24710_),
    .C_N(_23447_),
    .Y(_24721_));
 sky130_fd_sc_hd__o21bai_1 _44971_ (.A1(_24699_),
    .A2(_24710_),
    .B1_N(_23447_),
    .Y(_24732_));
 sky130_fd_sc_hd__and2b_1 _44972_ (.A_N(_24721_),
    .B(_24732_),
    .X(_24743_));
 sky130_fd_sc_hd__xor2_2 _44973_ (.A(_24281_),
    .B(_24743_),
    .X(_24754_));
 sky130_fd_sc_hd__xnor2_1 _44974_ (.A(_23469_),
    .B(_24754_),
    .Y(_24765_));
 sky130_fd_sc_hd__buf_1 _44975_ (.A(\delay_line[40][1] ),
    .X(_24776_));
 sky130_fd_sc_hd__and2b_1 _44976_ (.A_N(_22776_),
    .B(_24776_),
    .X(_24787_));
 sky130_fd_sc_hd__and2b_1 _44977_ (.A_N(_24776_),
    .B(_22787_),
    .X(_24798_));
 sky130_fd_sc_hd__buf_1 _44978_ (.A(\delay_line[6][1] ),
    .X(_24809_));
 sky130_fd_sc_hd__buf_2 _44979_ (.A(_24809_),
    .X(_24820_));
 sky130_fd_sc_hd__a21oi_1 _44980_ (.A1(_23029_),
    .A2(_23051_),
    .B1(_24820_),
    .Y(_24831_));
 sky130_fd_sc_hd__and3_1 _44981_ (.A(_23029_),
    .B(_23051_),
    .C(_24820_),
    .X(_24842_));
 sky130_fd_sc_hd__nor2_1 _44982_ (.A(_22831_),
    .B(net437),
    .Y(_24853_));
 sky130_fd_sc_hd__inv_2 _44983_ (.A(\delay_line[5][1] ),
    .Y(_24864_));
 sky130_fd_sc_hd__clkbuf_2 _44984_ (.A(_24864_),
    .X(_24875_));
 sky130_fd_sc_hd__and2_1 _44985_ (.A(_22831_),
    .B(net437),
    .X(_24886_));
 sky130_fd_sc_hd__or3_2 _44986_ (.A(_24853_),
    .B(_24875_),
    .C(_24886_),
    .X(_24897_));
 sky130_fd_sc_hd__o21ai_1 _44987_ (.A1(_24886_),
    .A2(_24853_),
    .B1(_24875_),
    .Y(_24908_));
 sky130_fd_sc_hd__a22o_1 _44988_ (.A1(_22820_),
    .A2(_22842_),
    .B1(_24897_),
    .B2(_24908_),
    .X(_24919_));
 sky130_fd_sc_hd__clkbuf_2 _44989_ (.A(\delay_line[2][1] ),
    .X(_24930_));
 sky130_fd_sc_hd__nand4_2 _44990_ (.A(_24897_),
    .B(_24908_),
    .C(_22820_),
    .D(_22842_),
    .Y(_24941_));
 sky130_fd_sc_hd__and3_1 _44991_ (.A(_24919_),
    .B(_24930_),
    .C(_24941_),
    .X(_24952_));
 sky130_fd_sc_hd__a21oi_1 _44992_ (.A1(_24941_),
    .A2(_24919_),
    .B1(_24930_),
    .Y(_24963_));
 sky130_fd_sc_hd__nor4_1 _44993_ (.A(_24831_),
    .B(_24842_),
    .C(_24952_),
    .D(_24963_),
    .Y(_24974_));
 sky130_fd_sc_hd__inv_2 _44994_ (.A(net213),
    .Y(_24985_));
 sky130_fd_sc_hd__clkbuf_2 _44995_ (.A(_24985_),
    .X(_24996_));
 sky130_fd_sc_hd__o22ai_2 _44996_ (.A1(_24831_),
    .A2(_24842_),
    .B1(_24952_),
    .B2(_24963_),
    .Y(_25007_));
 sky130_fd_sc_hd__and3_1 _44997_ (.A(_24996_),
    .B(_25007_),
    .C(_22941_),
    .X(_25018_));
 sky130_fd_sc_hd__a21oi_1 _44998_ (.A1(_24996_),
    .A2(_25007_),
    .B1(_22941_),
    .Y(_25029_));
 sky130_fd_sc_hd__clkbuf_2 _44999_ (.A(\delay_line[10][1] ),
    .X(_25040_));
 sky130_fd_sc_hd__clkbuf_2 _45000_ (.A(_25040_),
    .X(_25051_));
 sky130_fd_sc_hd__clkbuf_2 _45001_ (.A(_25051_),
    .X(_25062_));
 sky130_fd_sc_hd__clkbuf_2 _45002_ (.A(\delay_line[9][1] ),
    .X(_25073_));
 sky130_fd_sc_hd__xor2_2 _45003_ (.A(_23073_),
    .B(_25073_),
    .X(_25084_));
 sky130_fd_sc_hd__or2_1 _45004_ (.A(_25062_),
    .B(_25084_),
    .X(_25095_));
 sky130_fd_sc_hd__buf_1 _45005_ (.A(_25084_),
    .X(_25106_));
 sky130_fd_sc_hd__nand2_1 _45006_ (.A(_25062_),
    .B(_25106_),
    .Y(_25117_));
 sky130_fd_sc_hd__and4_1 _45007_ (.A(_25095_),
    .B(_23106_),
    .C(_23095_),
    .D(_25117_),
    .X(_25128_));
 sky130_fd_sc_hd__buf_1 _45008_ (.A(_25128_),
    .X(_25139_));
 sky130_fd_sc_hd__a22oi_4 _45009_ (.A1(_23095_),
    .A2(_23117_),
    .B1(_25117_),
    .B2(_25095_),
    .Y(_25150_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45010_ (.A(\delay_line[0][1] ),
    .X(_25161_));
 sky130_fd_sc_hd__and2b_1 _45011_ (.A_N(_23150_),
    .B(_25161_),
    .X(_25172_));
 sky130_fd_sc_hd__and2b_1 _45012_ (.A_N(_25161_),
    .B(_23161_),
    .X(_25183_));
 sky130_fd_sc_hd__clkbuf_4 _45013_ (.A(\delay_line[13][1] ),
    .X(_25194_));
 sky130_fd_sc_hd__o21ai_2 _45014_ (.A1(_25172_),
    .A2(_25183_),
    .B1(_25194_),
    .Y(_25204_));
 sky130_fd_sc_hd__inv_2 _45015_ (.A(\delay_line[13][1] ),
    .Y(_25215_));
 sky130_fd_sc_hd__nand2_1 _45016_ (.A(_23205_),
    .B(\delay_line[0][1] ),
    .Y(_25226_));
 sky130_fd_sc_hd__inv_2 _45017_ (.A(\delay_line[0][1] ),
    .Y(_25237_));
 sky130_fd_sc_hd__nand2_1 _45018_ (.A(_25237_),
    .B(_23172_),
    .Y(_25248_));
 sky130_fd_sc_hd__nand3_2 _45019_ (.A(_25215_),
    .B(_25226_),
    .C(_25248_),
    .Y(_25259_));
 sky130_fd_sc_hd__nand4_2 _45020_ (.A(_25204_),
    .B(_23172_),
    .C(net398),
    .D(_25259_),
    .Y(_25270_));
 sky130_fd_sc_hd__o2bb2ai_2 _45021_ (.A1_N(_25259_),
    .A2_N(_25204_),
    .B1(_23194_),
    .B2(_23205_),
    .Y(_25281_));
 sky130_fd_sc_hd__clkbuf_2 _45022_ (.A(\delay_line[12][1] ),
    .X(_25292_));
 sky130_fd_sc_hd__xor2_2 _45023_ (.A(\delay_line[12][0] ),
    .B(_25292_),
    .X(_25303_));
 sky130_fd_sc_hd__clkbuf_2 _45024_ (.A(_25303_),
    .X(_25314_));
 sky130_fd_sc_hd__a21oi_1 _45025_ (.A1(_25270_),
    .A2(_25281_),
    .B1(_25314_),
    .Y(_25325_));
 sky130_fd_sc_hd__and3_1 _45026_ (.A(_25281_),
    .B(_25314_),
    .C(_25270_),
    .X(_25336_));
 sky130_fd_sc_hd__nor3_2 _45027_ (.A(_25325_),
    .B(_23249_),
    .C(_25336_),
    .Y(_25347_));
 sky130_fd_sc_hd__o21a_1 _45028_ (.A1(_25336_),
    .A2(_25325_),
    .B1(_23249_),
    .X(_25358_));
 sky130_fd_sc_hd__o22ai_2 _45029_ (.A1(_25139_),
    .A2(_25150_),
    .B1(_25347_),
    .B2(_25358_),
    .Y(_25369_));
 sky130_fd_sc_hd__nor2_1 _45030_ (.A(_25128_),
    .B(_25150_),
    .Y(_25380_));
 sky130_fd_sc_hd__or2_1 _45031_ (.A(_23183_),
    .B(_23216_),
    .X(_25391_));
 sky130_fd_sc_hd__nand3_1 _45032_ (.A(_25281_),
    .B(_25314_),
    .C(_25270_),
    .Y(_25402_));
 sky130_fd_sc_hd__or4bb_1 _45033_ (.A(_25325_),
    .B(_25391_),
    .C_N(_23260_),
    .D_N(_25402_),
    .X(_25413_));
 sky130_fd_sc_hd__nand3b_1 _45034_ (.A_N(_25358_),
    .B(_25380_),
    .C(_25413_),
    .Y(_25424_));
 sky130_fd_sc_hd__and3_1 _45035_ (.A(_25369_),
    .B(_25424_),
    .C(_23293_),
    .X(_25435_));
 sky130_fd_sc_hd__a21oi_1 _45036_ (.A1(_25369_),
    .A2(_25424_),
    .B1(_23293_),
    .Y(_25446_));
 sky130_fd_sc_hd__buf_1 _45037_ (.A(\delay_line[7][1] ),
    .X(_00051_));
 sky130_fd_sc_hd__inv_2 _45038_ (.A(_00051_),
    .Y(_00062_));
 sky130_fd_sc_hd__buf_4 _45039_ (.A(_00062_),
    .X(_00073_));
 sky130_fd_sc_hd__nor2_1 _45040_ (.A(\delay_line[8][0] ),
    .B(\delay_line[8][1] ),
    .Y(_00084_));
 sky130_fd_sc_hd__and2_1 _45041_ (.A(\delay_line[8][0] ),
    .B(\delay_line[8][1] ),
    .X(_00095_));
 sky130_fd_sc_hd__nor2_1 _45042_ (.A(_00084_),
    .B(_00095_),
    .Y(_00106_));
 sky130_fd_sc_hd__buf_2 _45043_ (.A(_00106_),
    .X(_00117_));
 sky130_fd_sc_hd__xor2_2 _45044_ (.A(_00073_),
    .B(_00117_),
    .X(_00128_));
 sky130_fd_sc_hd__o21ai_2 _45045_ (.A1(_25435_),
    .A2(_25446_),
    .B1(_00128_),
    .Y(_00139_));
 sky130_fd_sc_hd__o41a_1 _45046_ (.A1(_25139_),
    .A2(_25150_),
    .A3(_25347_),
    .A4(_25358_),
    .B1(_23293_),
    .X(_00150_));
 sky130_fd_sc_hd__a211o_1 _45047_ (.A1(_00150_),
    .A2(_25369_),
    .B1(_00128_),
    .C1(_25446_),
    .X(_00161_));
 sky130_fd_sc_hd__a21o_1 _45048_ (.A1(_00139_),
    .A2(_00161_),
    .B1(net185),
    .X(_00172_));
 sky130_fd_sc_hd__nand3_2 _45049_ (.A(_00161_),
    .B(_23304_),
    .C(_00139_),
    .Y(_00183_));
 sky130_fd_sc_hd__a2bb2o_1 _45050_ (.A1_N(_25018_),
    .A2_N(_25029_),
    .B1(_00172_),
    .B2(_00183_),
    .X(_00194_));
 sky130_fd_sc_hd__nor2_1 _45051_ (.A(_25018_),
    .B(_25029_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand3_2 _45052_ (.A(_00172_),
    .B(_00183_),
    .C(_00205_),
    .Y(_00216_));
 sky130_fd_sc_hd__a21bo_1 _45053_ (.A1(_00194_),
    .A2(_00216_),
    .B1_N(_23337_),
    .X(_00227_));
 sky130_fd_sc_hd__nand3b_2 _45054_ (.A_N(_23337_),
    .B(_00194_),
    .C(_00216_),
    .Y(_00238_));
 sky130_fd_sc_hd__clkbuf_2 _45055_ (.A(\delay_line[1][1] ),
    .X(_00249_));
 sky130_fd_sc_hd__xor2_2 _45056_ (.A(\delay_line[1][0] ),
    .B(_00249_),
    .X(_00260_));
 sky130_fd_sc_hd__xnor2_2 _45057_ (.A(_22886_),
    .B(_00260_),
    .Y(_00271_));
 sky130_fd_sc_hd__a21oi_1 _45058_ (.A1(_00227_),
    .A2(_00238_),
    .B1(_00271_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand3_2 _45059_ (.A(_00227_),
    .B(_00238_),
    .C(_00271_),
    .Y(_00293_));
 sky130_fd_sc_hd__or2b_2 _45060_ (.A(_00282_),
    .B_N(_00293_),
    .X(_00304_));
 sky130_fd_sc_hd__xor2_4 _45061_ (.A(_23425_),
    .B(_00304_),
    .X(_00315_));
 sky130_fd_sc_hd__o21a_2 _45062_ (.A1(_24787_),
    .A2(_24798_),
    .B1(_00315_),
    .X(_00326_));
 sky130_fd_sc_hd__nor3_4 _45063_ (.A(_24787_),
    .B(_24798_),
    .C(_00315_),
    .Y(_00337_));
 sky130_fd_sc_hd__nor3b_1 _45064_ (.A(_00326_),
    .B(_00337_),
    .C_N(\delay_line[23][1] ),
    .Y(_00348_));
 sky130_fd_sc_hd__inv_2 _45065_ (.A(net93),
    .Y(_00359_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45066_ (.A(\delay_line[23][1] ),
    .X(_00370_));
 sky130_fd_sc_hd__o21bai_4 _45067_ (.A1(_00326_),
    .A2(_00337_),
    .B1_N(_00370_),
    .Y(_00381_));
 sky130_fd_sc_hd__buf_1 _45068_ (.A(\delay_line[39][1] ),
    .X(_00392_));
 sky130_fd_sc_hd__buf_1 _45069_ (.A(_00392_),
    .X(_00403_));
 sky130_fd_sc_hd__buf_1 _45070_ (.A(_00403_),
    .X(_00414_));
 sky130_fd_sc_hd__nor2_1 _45071_ (.A(_22765_),
    .B(_00414_),
    .Y(_00425_));
 sky130_fd_sc_hd__and2_1 _45072_ (.A(_22765_),
    .B(_00414_),
    .X(_00436_));
 sky130_fd_sc_hd__nor2_2 _45073_ (.A(_00425_),
    .B(_00436_),
    .Y(_00447_));
 sky130_fd_sc_hd__buf_2 _45074_ (.A(\delay_line[38][1] ),
    .X(_00458_));
 sky130_fd_sc_hd__xnor2_4 _45075_ (.A(_00458_),
    .B(net293),
    .Y(_00469_));
 sky130_fd_sc_hd__xnor2_4 _45076_ (.A(_00447_),
    .B(_00469_),
    .Y(_00480_));
 sky130_fd_sc_hd__a21oi_1 _45077_ (.A1(_00359_),
    .A2(_00381_),
    .B1(_00480_),
    .Y(_00491_));
 sky130_fd_sc_hd__and3_1 _45078_ (.A(_00359_),
    .B(_00381_),
    .C(_00480_),
    .X(_00502_));
 sky130_fd_sc_hd__nor2_1 _45079_ (.A(_00491_),
    .B(_00502_),
    .Y(_00513_));
 sky130_fd_sc_hd__a21bo_2 _45080_ (.A1(_22765_),
    .A2(_22787_),
    .B1_N(_23403_),
    .X(_00524_));
 sky130_fd_sc_hd__nor2_4 _45081_ (.A(net302),
    .B(\delay_line[35][1] ),
    .Y(_00535_));
 sky130_fd_sc_hd__and2_4 _45082_ (.A(net302),
    .B(\delay_line[35][1] ),
    .X(_00546_));
 sky130_fd_sc_hd__buf_1 _45083_ (.A(\delay_line[33][1] ),
    .X(_00557_));
 sky130_fd_sc_hd__clkbuf_2 _45084_ (.A(_00557_),
    .X(_00568_));
 sky130_fd_sc_hd__clkbuf_2 _45085_ (.A(_00568_),
    .X(_00579_));
 sky130_fd_sc_hd__clkbuf_2 _45086_ (.A(_00579_),
    .X(_00590_));
 sky130_fd_sc_hd__buf_2 _45087_ (.A(net308),
    .X(_00601_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45088_ (.A(_00601_),
    .X(_00612_));
 sky130_fd_sc_hd__and2_1 _45089_ (.A(_00590_),
    .B(_00612_),
    .X(_00623_));
 sky130_fd_sc_hd__nor2_1 _45090_ (.A(_00590_),
    .B(_00612_),
    .Y(_00634_));
 sky130_fd_sc_hd__or4_2 _45091_ (.A(_00535_),
    .B(_00546_),
    .C(_00623_),
    .D(_00634_),
    .X(_00645_));
 sky130_fd_sc_hd__o22ai_2 _45092_ (.A1(_00535_),
    .A2(_00546_),
    .B1(_00623_),
    .B2(_00634_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand3_1 _45093_ (.A(_00524_),
    .B(_00645_),
    .C(_00656_),
    .Y(_00667_));
 sky130_fd_sc_hd__a21o_1 _45094_ (.A1(_00645_),
    .A2(_00656_),
    .B1(_00524_),
    .X(_00678_));
 sky130_fd_sc_hd__and3_1 _45095_ (.A(_00513_),
    .B(_00667_),
    .C(_00678_),
    .X(_00689_));
 sky130_fd_sc_hd__o2bb2a_1 _45096_ (.A1_N(_00678_),
    .A2_N(_00667_),
    .B1(_00491_),
    .B2(_00502_),
    .X(_00700_));
 sky130_fd_sc_hd__or2_1 _45097_ (.A(_00689_),
    .B(_00700_),
    .X(_00711_));
 sky130_fd_sc_hd__nand2_1 _45098_ (.A(_24765_),
    .B(_00711_),
    .Y(_00722_));
 sky130_fd_sc_hd__or2_1 _45099_ (.A(_24765_),
    .B(_00711_),
    .X(_00733_));
 sky130_fd_sc_hd__and2_1 _45100_ (.A(_00722_),
    .B(_00733_),
    .X(_00744_));
 sky130_fd_sc_hd__buf_2 _45101_ (.A(_23513_),
    .X(_00755_));
 sky130_fd_sc_hd__and4_1 _45102_ (.A(_23480_),
    .B(_00744_),
    .C(_23491_),
    .D(_00755_),
    .X(_00766_));
 sky130_fd_sc_hd__a31o_1 _45103_ (.A1(_00755_),
    .A2(_23469_),
    .A3(_23491_),
    .B1(_00744_),
    .X(_00777_));
 sky130_fd_sc_hd__inv_2 _45104_ (.A(_00777_),
    .Y(_00788_));
 sky130_fd_sc_hd__nor4_1 _45105_ (.A(_23633_),
    .B(_23644_),
    .C(_00766_),
    .D(_00788_),
    .Y(_00799_));
 sky130_fd_sc_hd__o22a_1 _45106_ (.A1(_23633_),
    .A2(_23644_),
    .B1(_00766_),
    .B2(_00788_),
    .X(_00810_));
 sky130_fd_sc_hd__o2bb2a_1 _45107_ (.A1_N(_22205_),
    .A2_N(_23557_),
    .B1(net75),
    .B2(_00810_),
    .X(_00821_));
 sky130_fd_sc_hd__and4bb_1 _45108_ (.A_N(net75),
    .B_N(_00810_),
    .C(_22194_),
    .D(_23557_),
    .X(_00832_));
 sky130_fd_sc_hd__xor2_1 _45109_ (.A(\delay_line[17][1] ),
    .B(net378),
    .X(_00843_));
 sky130_fd_sc_hd__buf_2 _45110_ (.A(_00843_),
    .X(_00854_));
 sky130_fd_sc_hd__xor2_1 _45111_ (.A(_22205_),
    .B(_00854_),
    .X(_00865_));
 sky130_fd_sc_hd__o21a_1 _45112_ (.A1(_00821_),
    .A2(_00832_),
    .B1(_00865_),
    .X(_00876_));
 sky130_fd_sc_hd__nor3_1 _45113_ (.A(_00865_),
    .B(_00821_),
    .C(_00832_),
    .Y(_00887_));
 sky130_fd_sc_hd__nor2_1 _45114_ (.A(_00876_),
    .B(_00887_),
    .Y(_00898_));
 sky130_fd_sc_hd__xor2_1 _45115_ (.A(_23589_),
    .B(_00898_),
    .X(_00001_));
 sky130_fd_sc_hd__or3_2 _45116_ (.A(_22150_),
    .B(_23568_),
    .C(_00898_),
    .X(_00919_));
 sky130_fd_sc_hd__or3b_1 _45117_ (.A(_24281_),
    .B(net115),
    .C_N(_24732_),
    .X(_00930_));
 sky130_fd_sc_hd__o211ai_1 _45118_ (.A1(_22325_),
    .A2(_23655_),
    .B1(_23786_),
    .C1(_23764_),
    .Y(_00941_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45119_ (.A(\delay_line[31][2] ),
    .X(_00952_));
 sky130_fd_sc_hd__clkbuf_2 _45120_ (.A(_00952_),
    .X(_00963_));
 sky130_fd_sc_hd__o21ai_2 _45121_ (.A1(\delay_line[31][0] ),
    .A2(_24578_),
    .B1(_00963_),
    .Y(_00974_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45122_ (.A(_00963_),
    .X(_00985_));
 sky130_fd_sc_hd__or3_1 _45123_ (.A(_24567_),
    .B(_24589_),
    .C(_00985_),
    .X(_00996_));
 sky130_fd_sc_hd__clkbuf_2 _45124_ (.A(\delay_line[30][2] ),
    .X(_01007_));
 sky130_fd_sc_hd__buf_1 _45125_ (.A(_01007_),
    .X(_01018_));
 sky130_fd_sc_hd__buf_1 _45126_ (.A(_01018_),
    .X(_01029_));
 sky130_fd_sc_hd__buf_2 _45127_ (.A(_01029_),
    .X(_01040_));
 sky130_fd_sc_hd__buf_2 _45128_ (.A(\delay_line[29][0] ),
    .X(_01051_));
 sky130_fd_sc_hd__xor2_1 _45129_ (.A(_01040_),
    .B(_01051_),
    .X(_01062_));
 sky130_fd_sc_hd__a21o_1 _45130_ (.A1(_00974_),
    .A2(_00996_),
    .B1(_01062_),
    .X(_01073_));
 sky130_fd_sc_hd__nand3_1 _45131_ (.A(_00996_),
    .B(_01062_),
    .C(_00974_),
    .Y(_01084_));
 sky130_fd_sc_hd__nand2_2 _45132_ (.A(_01073_),
    .B(_01084_),
    .Y(_01095_));
 sky130_fd_sc_hd__inv_2 _45133_ (.A(\delay_line[28][1] ),
    .Y(_01106_));
 sky130_fd_sc_hd__buf_1 _45134_ (.A(\delay_line[28][2] ),
    .X(_01117_));
 sky130_fd_sc_hd__buf_2 _45135_ (.A(_01117_),
    .X(_01128_));
 sky130_fd_sc_hd__o21a_1 _45136_ (.A1(_22259_),
    .A2(_01106_),
    .B1(_01128_),
    .X(_01139_));
 sky130_fd_sc_hd__nor3_1 _45137_ (.A(_22270_),
    .B(_01128_),
    .C(_01106_),
    .Y(_01150_));
 sky130_fd_sc_hd__buf_1 _45138_ (.A(\delay_line[26][1] ),
    .X(_01161_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45139_ (.A(_01161_),
    .X(_01172_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45140_ (.A(\delay_line[27][2] ),
    .X(_01183_));
 sky130_fd_sc_hd__xor2_1 _45141_ (.A(\delay_line[27][0] ),
    .B(_01183_),
    .X(_01194_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45142_ (.A(_01194_),
    .X(_01205_));
 sky130_fd_sc_hd__or2_1 _45143_ (.A(_01172_),
    .B(_01205_),
    .X(_01216_));
 sky130_fd_sc_hd__nand2_1 _45144_ (.A(_01172_),
    .B(_01205_),
    .Y(_01227_));
 sky130_fd_sc_hd__o211a_1 _45145_ (.A1(_01139_),
    .A2(_01150_),
    .B1(_01216_),
    .C1(_01227_),
    .X(_01238_));
 sky130_fd_sc_hd__inv_2 _45146_ (.A(_01238_),
    .Y(_01249_));
 sky130_fd_sc_hd__a211o_1 _45147_ (.A1(_01216_),
    .A2(_01227_),
    .B1(_01139_),
    .C1(_01150_),
    .X(_01260_));
 sky130_fd_sc_hd__o21ai_1 _45148_ (.A1(_24336_),
    .A2(_24347_),
    .B1(_24413_),
    .Y(_01271_));
 sky130_fd_sc_hd__a21oi_2 _45149_ (.A1(_01249_),
    .A2(_01260_),
    .B1(_01271_),
    .Y(_01282_));
 sky130_fd_sc_hd__and3_1 _45150_ (.A(_01271_),
    .B(_01249_),
    .C(_01260_),
    .X(_01293_));
 sky130_fd_sc_hd__nor2_2 _45151_ (.A(_01282_),
    .B(_01293_),
    .Y(_01304_));
 sky130_fd_sc_hd__xor2_4 _45152_ (.A(_01095_),
    .B(_01304_),
    .X(_01315_));
 sky130_fd_sc_hd__a21oi_1 _45153_ (.A1(_00941_),
    .A2(_23841_),
    .B1(_01315_),
    .Y(_01326_));
 sky130_fd_sc_hd__and3_1 _45154_ (.A(_00941_),
    .B(_23841_),
    .C(_01315_),
    .X(_01337_));
 sky130_fd_sc_hd__nor2_1 _45155_ (.A(_01326_),
    .B(_01337_),
    .Y(_01348_));
 sky130_fd_sc_hd__o21a_1 _45156_ (.A1(_24435_),
    .A2(net184),
    .B1(_01348_),
    .X(_01359_));
 sky130_fd_sc_hd__nor3_1 _45157_ (.A(_24435_),
    .B(net184),
    .C(_01348_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _45158_ (.A(_01359_),
    .B(_01370_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand4_1 _45159_ (.A(_23830_),
    .B(_23841_),
    .C(_24215_),
    .D(_24226_),
    .Y(_01392_));
 sky130_fd_sc_hd__buf_1 _45160_ (.A(net356),
    .X(_01402_));
 sky130_fd_sc_hd__buf_1 _45161_ (.A(_01402_),
    .X(_01413_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45162_ (.A(_01413_),
    .X(_01424_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45163_ (.A(net345),
    .X(_01435_));
 sky130_fd_sc_hd__clkbuf_2 _45164_ (.A(_01435_),
    .X(_01446_));
 sky130_fd_sc_hd__buf_2 _45165_ (.A(_01446_),
    .X(_01457_));
 sky130_fd_sc_hd__nor2_1 _45166_ (.A(_01424_),
    .B(_01457_),
    .Y(_01468_));
 sky130_fd_sc_hd__and2_1 _45167_ (.A(_01424_),
    .B(_01457_),
    .X(_01479_));
 sky130_fd_sc_hd__buf_1 _45168_ (.A(\delay_line[25][2] ),
    .X(_01490_));
 sky130_fd_sc_hd__nor2_2 _45169_ (.A(\delay_line[25][0] ),
    .B(_01490_),
    .Y(_01501_));
 sky130_fd_sc_hd__and2_2 _45170_ (.A(\delay_line[25][0] ),
    .B(\delay_line[25][2] ),
    .X(_01512_));
 sky130_fd_sc_hd__or4_4 _45171_ (.A(_01468_),
    .B(_01479_),
    .C(_01501_),
    .D(_01512_),
    .X(_01523_));
 sky130_fd_sc_hd__o22ai_4 _45172_ (.A1(_01468_),
    .A2(_01479_),
    .B1(_01501_),
    .B2(_01512_),
    .Y(_01534_));
 sky130_fd_sc_hd__o211a_2 _45173_ (.A1(_23973_),
    .A2(_24028_),
    .B1(_01523_),
    .C1(_01534_),
    .X(_01545_));
 sky130_fd_sc_hd__a221oi_4 _45174_ (.A1(_23863_),
    .A2(_23907_),
    .B1(_01523_),
    .B2(_01534_),
    .C1(_24028_),
    .Y(_01556_));
 sky130_fd_sc_hd__o211ai_2 _45175_ (.A1(_01545_),
    .A2(_01556_),
    .B1(_23720_),
    .C1(_23786_),
    .Y(_01567_));
 sky130_fd_sc_hd__a211o_1 _45176_ (.A1(_23720_),
    .A2(_23786_),
    .B1(_01545_),
    .C1(_01556_),
    .X(_01578_));
 sky130_fd_sc_hd__and2b_2 _45177_ (.A_N(\delay_line[21][1] ),
    .B(\delay_line[21][0] ),
    .X(_01589_));
 sky130_fd_sc_hd__clkbuf_2 _45178_ (.A(\delay_line[21][1] ),
    .X(_01600_));
 sky130_fd_sc_hd__and2b_2 _45179_ (.A_N(_23984_),
    .B(_01600_),
    .X(_01611_));
 sky130_fd_sc_hd__nor2_2 _45180_ (.A(_01589_),
    .B(_01611_),
    .Y(_01622_));
 sky130_fd_sc_hd__and2b_2 _45181_ (.A_N(\delay_line[19][1] ),
    .B(\delay_line[19][0] ),
    .X(_01633_));
 sky130_fd_sc_hd__inv_2 _45182_ (.A(\delay_line[19][1] ),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_2 _45183_ (.A(\delay_line[19][0] ),
    .B(_01644_),
    .Y(_01655_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45184_ (.A(net375),
    .X(_01666_));
 sky130_fd_sc_hd__clkbuf_2 _45185_ (.A(_01666_),
    .X(_01677_));
 sky130_fd_sc_hd__clkbuf_4 _45186_ (.A(_01677_),
    .X(_01688_));
 sky130_fd_sc_hd__o21a_4 _45187_ (.A1(_01633_),
    .A2(_01655_),
    .B1(_01688_),
    .X(_01699_));
 sky130_fd_sc_hd__or2_4 _45188_ (.A(_01633_),
    .B(_01655_),
    .X(_01710_));
 sky130_fd_sc_hd__nor2_1 _45189_ (.A(_01688_),
    .B(_01710_),
    .Y(_01721_));
 sky130_fd_sc_hd__nor3_4 _45190_ (.A(_01622_),
    .B(_01699_),
    .C(_01721_),
    .Y(_01732_));
 sky130_fd_sc_hd__inv_2 _45191_ (.A(_01732_),
    .Y(_01743_));
 sky130_fd_sc_hd__o21ai_2 _45192_ (.A1(_01699_),
    .A2(_01721_),
    .B1(_01622_),
    .Y(_01754_));
 sky130_fd_sc_hd__clkbuf_2 _45193_ (.A(net393),
    .X(_01765_));
 sky130_fd_sc_hd__clkbuf_2 _45194_ (.A(_01765_),
    .X(_01776_));
 sky130_fd_sc_hd__buf_1 _45195_ (.A(\delay_line[15][2] ),
    .X(_01787_));
 sky130_fd_sc_hd__buf_1 _45196_ (.A(_01787_),
    .X(_01798_));
 sky130_fd_sc_hd__and2_1 _45197_ (.A(_22402_),
    .B(_01798_),
    .X(_01809_));
 sky130_fd_sc_hd__clkbuf_2 _45198_ (.A(_01798_),
    .X(_01820_));
 sky130_fd_sc_hd__nor2_1 _45199_ (.A(_22424_),
    .B(_01820_),
    .Y(_01831_));
 sky130_fd_sc_hd__nor2_1 _45200_ (.A(_01809_),
    .B(_01831_),
    .Y(_01842_));
 sky130_fd_sc_hd__or2_1 _45201_ (.A(_01776_),
    .B(_01842_),
    .X(_01853_));
 sky130_fd_sc_hd__buf_1 _45202_ (.A(\delay_line[16][1] ),
    .X(_01864_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45203_ (.A(_01864_),
    .X(_01875_));
 sky130_fd_sc_hd__buf_2 _45204_ (.A(_01875_),
    .X(_01886_));
 sky130_fd_sc_hd__or3b_2 _45205_ (.A(_01809_),
    .B(_01831_),
    .C_N(_01776_),
    .X(_01897_));
 sky130_fd_sc_hd__and3_4 _45206_ (.A(_01853_),
    .B(_01886_),
    .C(_01897_),
    .X(_01908_));
 sky130_fd_sc_hd__a21oi_4 _45207_ (.A1(_01897_),
    .A2(_01853_),
    .B1(_01886_),
    .Y(_01919_));
 sky130_fd_sc_hd__a211o_1 _45208_ (.A1(_24116_),
    .A2(_24160_),
    .B1(_01908_),
    .C1(_01919_),
    .X(_01930_));
 sky130_fd_sc_hd__o211ai_2 _45209_ (.A1(_01908_),
    .A2(_01919_),
    .B1(_24116_),
    .C1(_24160_),
    .Y(_01941_));
 sky130_fd_sc_hd__and4_2 _45210_ (.A(_01743_),
    .B(_01754_),
    .C(_01930_),
    .D(_01941_),
    .X(_01952_));
 sky130_fd_sc_hd__a22oi_4 _45211_ (.A1(_01743_),
    .A2(_01754_),
    .B1(_01930_),
    .B2(_01941_),
    .Y(_01963_));
 sky130_fd_sc_hd__a211o_1 _45212_ (.A1(_24171_),
    .A2(_24193_),
    .B1(_01952_),
    .C1(_01963_),
    .X(_01974_));
 sky130_fd_sc_hd__o211ai_2 _45213_ (.A1(_01952_),
    .A2(_01963_),
    .B1(_24171_),
    .C1(_24193_),
    .Y(_01985_));
 sky130_fd_sc_hd__and4_1 _45214_ (.A(_01567_),
    .B(_01578_),
    .C(_01974_),
    .D(_01985_),
    .X(_01996_));
 sky130_fd_sc_hd__a22oi_1 _45215_ (.A1(_01567_),
    .A2(_01578_),
    .B1(_01974_),
    .B2(_01985_),
    .Y(_02007_));
 sky130_fd_sc_hd__or2_1 _45216_ (.A(_01996_),
    .B(_02007_),
    .X(_02018_));
 sky130_fd_sc_hd__and3_1 _45217_ (.A(_24215_),
    .B(_01392_),
    .C(_02018_),
    .X(_02029_));
 sky130_fd_sc_hd__a21oi_1 _45218_ (.A1(_24215_),
    .A2(_01392_),
    .B1(_02018_),
    .Y(_02040_));
 sky130_fd_sc_hd__nor2_1 _45219_ (.A(_02029_),
    .B(_02040_),
    .Y(_02051_));
 sky130_fd_sc_hd__xnor2_1 _45220_ (.A(_01381_),
    .B(_02051_),
    .Y(_02062_));
 sky130_fd_sc_hd__a21o_1 _45221_ (.A1(_24259_),
    .A2(_00930_),
    .B1(_02062_),
    .X(_02073_));
 sky130_fd_sc_hd__inv_2 _45222_ (.A(_02073_),
    .Y(_02084_));
 sky130_fd_sc_hd__and3_1 _45223_ (.A(_24259_),
    .B(_00930_),
    .C(_02062_),
    .X(_02095_));
 sky130_fd_sc_hd__clkbuf_2 _45224_ (.A(\delay_line[32][2] ),
    .X(_02106_));
 sky130_fd_sc_hd__clkbuf_2 _45225_ (.A(_02106_),
    .X(_02117_));
 sky130_fd_sc_hd__clkbuf_2 _45226_ (.A(_02117_),
    .X(_02128_));
 sky130_fd_sc_hd__or3_1 _45227_ (.A(_22567_),
    .B(_24479_),
    .C(_02128_),
    .X(_02139_));
 sky130_fd_sc_hd__buf_1 _45228_ (.A(net314),
    .X(_02150_));
 sky130_fd_sc_hd__buf_1 _45229_ (.A(_02150_),
    .X(_02161_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45230_ (.A(_02161_),
    .X(_02172_));
 sky130_fd_sc_hd__clkbuf_2 _45231_ (.A(_02172_),
    .X(_02183_));
 sky130_fd_sc_hd__o21ai_1 _45232_ (.A1(_22567_),
    .A2(_24479_),
    .B1(_02128_),
    .Y(_02194_));
 sky130_fd_sc_hd__and3_1 _45233_ (.A(_02139_),
    .B(_02183_),
    .C(_02194_),
    .X(_02205_));
 sky130_fd_sc_hd__a21oi_1 _45234_ (.A1(_02194_),
    .A2(_02139_),
    .B1(_02183_),
    .Y(_02216_));
 sky130_fd_sc_hd__or2_1 _45235_ (.A(_02205_),
    .B(_02216_),
    .X(_02227_));
 sky130_fd_sc_hd__buf_1 _45236_ (.A(net307),
    .X(_02238_));
 sky130_fd_sc_hd__clkbuf_2 _45237_ (.A(_02238_),
    .X(_02249_));
 sky130_fd_sc_hd__clkbuf_2 _45238_ (.A(_02249_),
    .X(_02260_));
 sky130_fd_sc_hd__or2b_2 _45239_ (.A(_02260_),
    .B_N(_22611_),
    .X(_02271_));
 sky130_fd_sc_hd__or2b_1 _45240_ (.A(_22622_),
    .B_N(_02260_),
    .X(_02282_));
 sky130_fd_sc_hd__and3_1 _45241_ (.A(_02227_),
    .B(_02271_),
    .C(_02282_),
    .X(_02293_));
 sky130_fd_sc_hd__a21oi_2 _45242_ (.A1(_02271_),
    .A2(_02282_),
    .B1(_02227_),
    .Y(_02304_));
 sky130_fd_sc_hd__o211ai_1 _45243_ (.A1(_02293_),
    .A2(_02304_),
    .B1(_24644_),
    .C1(_24677_),
    .Y(_02315_));
 sky130_fd_sc_hd__a211o_1 _45244_ (.A1(_24644_),
    .A2(_24677_),
    .B1(_02293_),
    .C1(_02304_),
    .X(_02326_));
 sky130_fd_sc_hd__a21bo_1 _45245_ (.A1(_00590_),
    .A2(_00612_),
    .B1_N(_00645_),
    .X(_02337_));
 sky130_fd_sc_hd__a21oi_1 _45246_ (.A1(_02315_),
    .A2(_02326_),
    .B1(_02337_),
    .Y(_02348_));
 sky130_fd_sc_hd__and3_1 _45247_ (.A(_02337_),
    .B(_02315_),
    .C(_02326_),
    .X(_02359_));
 sky130_fd_sc_hd__or3_1 _45248_ (.A(_02348_),
    .B(_02359_),
    .C(_00667_),
    .X(_02370_));
 sky130_fd_sc_hd__o21ai_1 _45249_ (.A1(_02348_),
    .A2(_02359_),
    .B1(_00667_),
    .Y(_02381_));
 sky130_fd_sc_hd__nand2_1 _45250_ (.A(_00183_),
    .B(_00216_),
    .Y(_02392_));
 sky130_fd_sc_hd__inv_2 _45251_ (.A(_25424_),
    .Y(_02403_));
 sky130_fd_sc_hd__buf_1 _45252_ (.A(\delay_line[12][2] ),
    .X(_02414_));
 sky130_fd_sc_hd__clkbuf_2 _45253_ (.A(_02414_),
    .X(_02425_));
 sky130_fd_sc_hd__inv_2 _45254_ (.A(\delay_line[12][1] ),
    .Y(_02436_));
 sky130_fd_sc_hd__clkbuf_2 _45255_ (.A(_02436_),
    .X(_02447_));
 sky130_fd_sc_hd__nor3_2 _45256_ (.A(_23227_),
    .B(_02425_),
    .C(_02447_),
    .Y(_02458_));
 sky130_fd_sc_hd__o21a_1 _45257_ (.A1(_23227_),
    .A2(_02447_),
    .B1(_02425_),
    .X(_02469_));
 sky130_fd_sc_hd__clkbuf_2 _45258_ (.A(\delay_line[13][2] ),
    .X(_02480_));
 sky130_fd_sc_hd__inv_2 _45259_ (.A(_02480_),
    .Y(_02491_));
 sky130_fd_sc_hd__clkbuf_2 _45260_ (.A(\delay_line[11][0] ),
    .X(_02502_));
 sky130_fd_sc_hd__clkbuf_2 _45261_ (.A(_02502_),
    .X(_02513_));
 sky130_fd_sc_hd__buf_1 _45262_ (.A(\delay_line[0][2] ),
    .X(_02524_));
 sky130_fd_sc_hd__and2b_1 _45263_ (.A_N(_02513_),
    .B(_02524_),
    .X(_02535_));
 sky130_fd_sc_hd__nor2b_1 _45264_ (.A(_02524_),
    .B_N(_02513_),
    .Y(_02546_));
 sky130_fd_sc_hd__o21ai_1 _45265_ (.A1(_02535_),
    .A2(_02546_),
    .B1(_25172_),
    .Y(_02557_));
 sky130_fd_sc_hd__or2b_1 _45266_ (.A(\delay_line[0][2] ),
    .B_N(_02502_),
    .X(_02568_));
 sky130_fd_sc_hd__inv_2 _45267_ (.A(_02502_),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _45268_ (.A(_02579_),
    .B(_02524_),
    .Y(_02590_));
 sky130_fd_sc_hd__o211ai_1 _45269_ (.A1(_25237_),
    .A2(_23161_),
    .B1(_02568_),
    .C1(_02590_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand3_2 _45270_ (.A(_02491_),
    .B(_02557_),
    .C(_02601_),
    .Y(_02612_));
 sky130_fd_sc_hd__o21ai_1 _45271_ (.A1(_02535_),
    .A2(_02546_),
    .B1(_25226_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand4_2 _45272_ (.A(_23205_),
    .B(_02590_),
    .C(_02568_),
    .D(_25161_),
    .Y(_02634_));
 sky130_fd_sc_hd__nand3_2 _45273_ (.A(_02623_),
    .B(_02634_),
    .C(_02480_),
    .Y(_02645_));
 sky130_fd_sc_hd__a21oi_1 _45274_ (.A1(_25226_),
    .A2(_25248_),
    .B1(_25215_),
    .Y(_02656_));
 sky130_fd_sc_hd__a21o_1 _45275_ (.A1(_02612_),
    .A2(_02645_),
    .B1(_02656_),
    .X(_02667_));
 sky130_fd_sc_hd__o2111ai_4 _45276_ (.A1(_25172_),
    .A2(_25183_),
    .B1(_02645_),
    .C1(_25194_),
    .D1(_02612_),
    .Y(_02678_));
 sky130_fd_sc_hd__buf_1 _45277_ (.A(_23194_),
    .X(_02689_));
 sky130_fd_sc_hd__a31o_1 _45278_ (.A1(_25204_),
    .A2(_23172_),
    .A3(_25259_),
    .B1(_02689_),
    .X(_02700_));
 sky130_fd_sc_hd__a21oi_1 _45279_ (.A1(_02667_),
    .A2(_02678_),
    .B1(_02700_),
    .Y(_02711_));
 sky130_fd_sc_hd__and3_1 _45280_ (.A(_25204_),
    .B(_23216_),
    .C(_25259_),
    .X(_02722_));
 sky130_fd_sc_hd__o211a_1 _45281_ (.A1(_02722_),
    .A2(_02689_),
    .B1(_02678_),
    .C1(_02667_),
    .X(_02733_));
 sky130_fd_sc_hd__o22a_2 _45282_ (.A1(_02458_),
    .A2(_02469_),
    .B1(_02711_),
    .B2(_02733_),
    .X(_02744_));
 sky130_fd_sc_hd__a21oi_1 _45283_ (.A1(_02612_),
    .A2(_02645_),
    .B1(_02656_),
    .Y(_02755_));
 sky130_fd_sc_hd__and3_1 _45284_ (.A(_02612_),
    .B(_02645_),
    .C(_02656_),
    .X(_02766_));
 sky130_fd_sc_hd__o21bai_1 _45285_ (.A1(_02755_),
    .A2(_02766_),
    .B1_N(_02700_),
    .Y(_02777_));
 sky130_fd_sc_hd__o211ai_1 _45286_ (.A1(_02722_),
    .A2(_02689_),
    .B1(_02678_),
    .C1(_02667_),
    .Y(_02788_));
 sky130_fd_sc_hd__nor2_2 _45287_ (.A(_02458_),
    .B(_02469_),
    .Y(_02799_));
 sky130_fd_sc_hd__a31o_1 _45288_ (.A1(_02777_),
    .A2(_02788_),
    .A3(_02799_),
    .B1(_25402_),
    .X(_02810_));
 sky130_fd_sc_hd__buf_1 _45289_ (.A(net414),
    .X(_02821_));
 sky130_fd_sc_hd__buf_2 _45290_ (.A(_02821_),
    .X(_02832_));
 sky130_fd_sc_hd__clkbuf_2 _45291_ (.A(\delay_line[9][2] ),
    .X(_02843_));
 sky130_fd_sc_hd__buf_1 _45292_ (.A(_02843_),
    .X(_02854_));
 sky130_fd_sc_hd__and3b_2 _45293_ (.A_N(_02854_),
    .B(_25073_),
    .C(_23073_),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_2 _45294_ (.A(_25073_),
    .X(_02876_));
 sky130_fd_sc_hd__a21boi_2 _45295_ (.A1(_23073_),
    .A2(_02876_),
    .B1_N(_02854_),
    .Y(_02887_));
 sky130_fd_sc_hd__or3_1 _45296_ (.A(_02832_),
    .B(_02865_),
    .C(_02887_),
    .X(_02898_));
 sky130_fd_sc_hd__o21ai_2 _45297_ (.A1(_02865_),
    .A2(_02887_),
    .B1(_02832_),
    .Y(_02909_));
 sky130_fd_sc_hd__a22oi_1 _45298_ (.A1(_25062_),
    .A2(_25106_),
    .B1(_02898_),
    .B2(_02909_),
    .Y(_02920_));
 sky130_fd_sc_hd__and4_1 _45299_ (.A(_02898_),
    .B(_02909_),
    .C(_25062_),
    .D(_25106_),
    .X(_02931_));
 sky130_fd_sc_hd__nor2_1 _45300_ (.A(_02920_),
    .B(_02931_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand3_1 _45301_ (.A(_02777_),
    .B(_02788_),
    .C(_02799_),
    .Y(_02953_));
 sky130_fd_sc_hd__o22ai_2 _45302_ (.A1(_02458_),
    .A2(_02469_),
    .B1(_02711_),
    .B2(_02733_),
    .Y(_02964_));
 sky130_fd_sc_hd__a21o_1 _45303_ (.A1(_02953_),
    .A2(_02964_),
    .B1(_25336_),
    .X(_02975_));
 sky130_fd_sc_hd__o211ai_2 _45304_ (.A1(_02744_),
    .A2(_02810_),
    .B1(_02942_),
    .C1(_02975_),
    .Y(_02986_));
 sky130_fd_sc_hd__inv_2 _45305_ (.A(_25314_),
    .Y(_02996_));
 sky130_fd_sc_hd__nand2_1 _45306_ (.A(_25270_),
    .B(_25281_),
    .Y(_03007_));
 sky130_fd_sc_hd__a2bb2oi_1 _45307_ (.A1_N(_02996_),
    .A2_N(_03007_),
    .B1(_02953_),
    .B2(_02964_),
    .Y(_03018_));
 sky130_fd_sc_hd__nor2_1 _45308_ (.A(_02744_),
    .B(_02810_),
    .Y(_03029_));
 sky130_fd_sc_hd__or2_1 _45309_ (.A(_02920_),
    .B(_02931_),
    .X(_03040_));
 sky130_fd_sc_hd__o21ai_1 _45310_ (.A1(_03018_),
    .A2(_03029_),
    .B1(_03040_),
    .Y(_03051_));
 sky130_fd_sc_hd__o211ai_4 _45311_ (.A1(_25347_),
    .A2(_02403_),
    .B1(_02986_),
    .C1(_03051_),
    .Y(_03062_));
 sky130_fd_sc_hd__o21ai_1 _45312_ (.A1(_03018_),
    .A2(_03029_),
    .B1(_02942_),
    .Y(_03073_));
 sky130_fd_sc_hd__o31a_1 _45313_ (.A1(_25128_),
    .A2(_25150_),
    .A3(_25358_),
    .B1(_25413_),
    .X(_03084_));
 sky130_fd_sc_hd__nand3_1 _45314_ (.A(_02964_),
    .B(_25336_),
    .C(_02953_),
    .Y(_03095_));
 sky130_fd_sc_hd__nand3_1 _45315_ (.A(_02975_),
    .B(_03095_),
    .C(_03040_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand3_2 _45316_ (.A(_03073_),
    .B(_03084_),
    .C(_03106_),
    .Y(_03117_));
 sky130_fd_sc_hd__inv_2 _45317_ (.A(\delay_line[7][2] ),
    .Y(_03128_));
 sky130_fd_sc_hd__clkbuf_2 _45318_ (.A(_03128_),
    .X(_03139_));
 sky130_fd_sc_hd__clkbuf_2 _45319_ (.A(\delay_line[8][1] ),
    .X(_03150_));
 sky130_fd_sc_hd__clkbuf_2 _45320_ (.A(_03150_),
    .X(_03161_));
 sky130_fd_sc_hd__buf_1 _45321_ (.A(\delay_line[8][2] ),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_2 _45322_ (.A(_03172_),
    .X(_03183_));
 sky130_fd_sc_hd__o21a_1 _45323_ (.A1(_22985_),
    .A2(_03161_),
    .B1(_03183_),
    .X(_03194_));
 sky130_fd_sc_hd__clkbuf_2 _45324_ (.A(\delay_line[8][2] ),
    .X(_03205_));
 sky130_fd_sc_hd__nor3_1 _45325_ (.A(\delay_line[8][0] ),
    .B(_03150_),
    .C(_03205_),
    .Y(_03216_));
 sky130_fd_sc_hd__or3_4 _45326_ (.A(_03139_),
    .B(_03194_),
    .C(net280),
    .X(_03227_));
 sky130_fd_sc_hd__buf_2 _45327_ (.A(_03139_),
    .X(_03238_));
 sky130_fd_sc_hd__o21ai_2 _45328_ (.A1(_03194_),
    .A2(net280),
    .B1(_03238_),
    .Y(_03249_));
 sky130_fd_sc_hd__and3_1 _45329_ (.A(_03227_),
    .B(_03249_),
    .C(_25106_),
    .X(_03260_));
 sky130_fd_sc_hd__clkbuf_2 _45330_ (.A(_03260_),
    .X(_03271_));
 sky130_fd_sc_hd__a21oi_1 _45331_ (.A1(_03227_),
    .A2(_03249_),
    .B1(_25106_),
    .Y(_03282_));
 sky130_fd_sc_hd__nor3b_1 _45332_ (.A(_03271_),
    .B(_03282_),
    .C_N(_25139_),
    .Y(_03293_));
 sky130_fd_sc_hd__o21ba_1 _45333_ (.A1(_03260_),
    .A2(_03282_),
    .B1_N(_25139_),
    .X(_03304_));
 sky130_fd_sc_hd__nor2_1 _45334_ (.A(_03293_),
    .B(_03304_),
    .Y(_03315_));
 sky130_fd_sc_hd__a21oi_1 _45335_ (.A1(_03062_),
    .A2(_03117_),
    .B1(_03315_),
    .Y(_03326_));
 sky130_fd_sc_hd__and3_1 _45336_ (.A(_03062_),
    .B(_03117_),
    .C(_03315_),
    .X(_03337_));
 sky130_fd_sc_hd__a2bb2o_1 _45337_ (.A1_N(_00128_),
    .A2_N(_25446_),
    .B1(_00150_),
    .B2(_25369_),
    .X(_03348_));
 sky130_fd_sc_hd__o21bai_2 _45338_ (.A1(_03326_),
    .A2(_03337_),
    .B1_N(_03348_),
    .Y(_03359_));
 sky130_fd_sc_hd__a21o_1 _45339_ (.A1(_03062_),
    .A2(_03117_),
    .B1(_03315_),
    .X(_03370_));
 sky130_fd_sc_hd__nand3_1 _45340_ (.A(_03062_),
    .B(_03117_),
    .C(_03315_),
    .Y(_03381_));
 sky130_fd_sc_hd__nand3_1 _45341_ (.A(_03348_),
    .B(_03370_),
    .C(_03381_),
    .Y(_03392_));
 sky130_fd_sc_hd__buf_1 _45342_ (.A(\delay_line[6][2] ),
    .X(_03403_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45343_ (.A(_03403_),
    .X(_03414_));
 sky130_fd_sc_hd__buf_2 _45344_ (.A(_03414_),
    .X(_03425_));
 sky130_fd_sc_hd__or4b_4 _45345_ (.A(_00073_),
    .B(_00084_),
    .C(_00095_),
    .D_N(_03425_),
    .X(_03436_));
 sky130_fd_sc_hd__clkbuf_2 _45346_ (.A(_00051_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_4 _45347_ (.A(_03447_),
    .X(_03458_));
 sky130_fd_sc_hd__a21o_1 _45348_ (.A1(_03458_),
    .A2(_00117_),
    .B1(_03425_),
    .X(_03469_));
 sky130_fd_sc_hd__nand4_1 _45349_ (.A(_03436_),
    .B(_03469_),
    .C(_24820_),
    .D(_23007_),
    .Y(_03480_));
 sky130_fd_sc_hd__a32o_1 _45350_ (.A1(_23029_),
    .A2(_23051_),
    .A3(_24820_),
    .B1(_03436_),
    .B2(_03469_),
    .X(_03491_));
 sky130_fd_sc_hd__clkbuf_2 _45351_ (.A(\delay_line[3][2] ),
    .X(_03502_));
 sky130_fd_sc_hd__nor2_1 _45352_ (.A(_22831_),
    .B(_03502_),
    .Y(_03513_));
 sky130_fd_sc_hd__and2_1 _45353_ (.A(\delay_line[5][0] ),
    .B(_03502_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_2 _45354_ (.A(net431),
    .X(_03535_));
 sky130_fd_sc_hd__buf_4 _45355_ (.A(_03535_),
    .X(_03546_));
 sky130_fd_sc_hd__nand2_1 _45356_ (.A(_24875_),
    .B(_03546_),
    .Y(_03557_));
 sky130_fd_sc_hd__inv_2 _45357_ (.A(_03535_),
    .Y(_03568_));
 sky130_fd_sc_hd__buf_2 _45358_ (.A(\delay_line[5][1] ),
    .X(_03579_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45359_ (.A(_03579_),
    .X(_03590_));
 sky130_fd_sc_hd__nand2_1 _45360_ (.A(_03568_),
    .B(_03590_),
    .Y(_03601_));
 sky130_fd_sc_hd__o211ai_2 _45361_ (.A1(_03513_),
    .A2(_03524_),
    .B1(_03557_),
    .C1(_03601_),
    .Y(_03612_));
 sky130_fd_sc_hd__a211o_1 _45362_ (.A1(_03557_),
    .A2(_03601_),
    .B1(_03513_),
    .C1(_03524_),
    .X(_03623_));
 sky130_fd_sc_hd__a21oi_1 _45363_ (.A1(_03612_),
    .A2(_03623_),
    .B1(_22919_),
    .Y(_03634_));
 sky130_fd_sc_hd__and3_2 _45364_ (.A(_03623_),
    .B(_22908_),
    .C(_03612_),
    .X(_03645_));
 sky130_fd_sc_hd__or3_2 _45365_ (.A(_03634_),
    .B(_24897_),
    .C(_03645_),
    .X(_03656_));
 sky130_fd_sc_hd__o21ai_1 _45366_ (.A1(_03645_),
    .A2(_03634_),
    .B1(_24897_),
    .Y(_03667_));
 sky130_fd_sc_hd__inv_2 _45367_ (.A(\delay_line[2][2] ),
    .Y(_03678_));
 sky130_fd_sc_hd__or2_1 _45368_ (.A(\delay_line[3][0] ),
    .B(_03678_),
    .X(_03689_));
 sky130_fd_sc_hd__nand2_1 _45369_ (.A(_03678_),
    .B(_22820_),
    .Y(_03700_));
 sky130_fd_sc_hd__and3_1 _45370_ (.A(_03689_),
    .B(_03700_),
    .C(_24886_),
    .X(_03711_));
 sky130_fd_sc_hd__a21oi_1 _45371_ (.A1(_03689_),
    .A2(_03700_),
    .B1(_24886_),
    .Y(_03722_));
 sky130_fd_sc_hd__or2_1 _45372_ (.A(_03711_),
    .B(_03722_),
    .X(_03733_));
 sky130_fd_sc_hd__a21bo_1 _45373_ (.A1(_03656_),
    .A2(_03667_),
    .B1_N(_03733_),
    .X(_03744_));
 sky130_fd_sc_hd__nand3b_2 _45374_ (.A_N(_03733_),
    .B(_03656_),
    .C(_03667_),
    .Y(_03755_));
 sky130_fd_sc_hd__a22oi_1 _45375_ (.A1(_03480_),
    .A2(_03491_),
    .B1(_03744_),
    .B2(_03755_),
    .Y(_03766_));
 sky130_fd_sc_hd__nand4_1 _45376_ (.A(_03480_),
    .B(_03491_),
    .C(_03744_),
    .D(_03755_),
    .Y(_03777_));
 sky130_fd_sc_hd__or2b_2 _45377_ (.A(_03766_),
    .B_N(_03777_),
    .X(_03788_));
 sky130_fd_sc_hd__xor2_2 _45378_ (.A(_24996_),
    .B(_03788_),
    .X(_03799_));
 sky130_fd_sc_hd__a21o_1 _45379_ (.A1(_03359_),
    .A2(_03392_),
    .B1(_03799_),
    .X(_03810_));
 sky130_fd_sc_hd__nand2_1 _45380_ (.A(_03348_),
    .B(_03370_),
    .Y(_03821_));
 sky130_fd_sc_hd__o211ai_1 _45381_ (.A1(_03337_),
    .A2(_03821_),
    .B1(_03359_),
    .C1(_03799_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand3_2 _45382_ (.A(_02392_),
    .B(_03810_),
    .C(_03832_),
    .Y(_03843_));
 sky130_fd_sc_hd__a21oi_1 _45383_ (.A1(_03359_),
    .A2(_03392_),
    .B1(_03799_),
    .Y(_03854_));
 sky130_fd_sc_hd__o211a_1 _45384_ (.A1(_03337_),
    .A2(_03821_),
    .B1(_03359_),
    .C1(_03799_),
    .X(_03865_));
 sky130_fd_sc_hd__o21bai_1 _45385_ (.A1(_03854_),
    .A2(_03865_),
    .B1_N(_02392_),
    .Y(_03876_));
 sky130_fd_sc_hd__clkbuf_2 _45386_ (.A(_00249_),
    .X(_03887_));
 sky130_fd_sc_hd__buf_1 _45387_ (.A(\delay_line[1][2] ),
    .X(_03898_));
 sky130_fd_sc_hd__clkbuf_2 _45388_ (.A(_03898_),
    .X(_03909_));
 sky130_fd_sc_hd__o21a_1 _45389_ (.A1(_23370_),
    .A2(_03887_),
    .B1(_03909_),
    .X(_03920_));
 sky130_fd_sc_hd__nor3_1 _45390_ (.A(_23370_),
    .B(_03887_),
    .C(_03909_),
    .Y(_03931_));
 sky130_fd_sc_hd__nand3_1 _45391_ (.A(_24919_),
    .B(_24930_),
    .C(_24941_),
    .Y(_03942_));
 sky130_fd_sc_hd__o211a_1 _45392_ (.A1(_03920_),
    .A2(_03931_),
    .B1(_24941_),
    .C1(_03942_),
    .X(_03953_));
 sky130_fd_sc_hd__a211oi_2 _45393_ (.A1(_24941_),
    .A2(_03942_),
    .B1(_03920_),
    .C1(_03931_),
    .Y(_03964_));
 sky130_fd_sc_hd__or4b_4 _45394_ (.A(_22886_),
    .B(_03953_),
    .C(_03964_),
    .D_N(_00260_),
    .X(_03975_));
 sky130_fd_sc_hd__and4bb_1 _45395_ (.A_N(_22853_),
    .B_N(_22864_),
    .C(_00260_),
    .D(_22875_),
    .X(_03986_));
 sky130_fd_sc_hd__nor2_1 _45396_ (.A(_03953_),
    .B(_03964_),
    .Y(_03997_));
 sky130_fd_sc_hd__or2_1 _45397_ (.A(_03986_),
    .B(_03997_),
    .X(_04008_));
 sky130_fd_sc_hd__and3_1 _45398_ (.A(_03975_),
    .B(_04008_),
    .C(_25018_),
    .X(_04019_));
 sky130_fd_sc_hd__a21oi_2 _45399_ (.A1(_03975_),
    .A2(_04008_),
    .B1(_25018_),
    .Y(_04030_));
 sky130_fd_sc_hd__a211o_1 _45400_ (.A1(_03843_),
    .A2(_03876_),
    .B1(_04019_),
    .C1(_04030_),
    .X(_04041_));
 sky130_fd_sc_hd__buf_2 _45401_ (.A(_04019_),
    .X(_04052_));
 sky130_fd_sc_hd__o211ai_2 _45402_ (.A1(_04052_),
    .A2(_04030_),
    .B1(_03843_),
    .C1(_03876_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand4_2 _45403_ (.A(_00238_),
    .B(_00293_),
    .C(_04041_),
    .D(_04063_),
    .Y(_04074_));
 sky130_fd_sc_hd__nand4b_4 _45404_ (.A_N(_00282_),
    .B(_00293_),
    .C(_04074_),
    .D(_23381_),
    .Y(_04085_));
 sky130_fd_sc_hd__a22o_1 _45405_ (.A1(_00238_),
    .A2(_00293_),
    .B1(_04041_),
    .B2(_04063_),
    .X(_04096_));
 sky130_fd_sc_hd__a2bb2o_2 _45406_ (.A1_N(_23425_),
    .A2_N(_00304_),
    .B1(_04074_),
    .B2(_04096_),
    .X(_04107_));
 sky130_fd_sc_hd__buf_1 _45407_ (.A(\delay_line[39][2] ),
    .X(_04118_));
 sky130_fd_sc_hd__buf_1 _45408_ (.A(_04118_),
    .X(_04129_));
 sky130_fd_sc_hd__buf_1 _45409_ (.A(_04129_),
    .X(_04140_));
 sky130_fd_sc_hd__o21ai_1 _45410_ (.A1(_22754_),
    .A2(_00414_),
    .B1(_04140_),
    .Y(_04151_));
 sky130_fd_sc_hd__or3_1 _45411_ (.A(_22754_),
    .B(_00414_),
    .C(_04140_),
    .X(_04162_));
 sky130_fd_sc_hd__buf_1 _45412_ (.A(\delay_line[40][2] ),
    .X(_04173_));
 sky130_fd_sc_hd__nor2_1 _45413_ (.A(_04173_),
    .B(_24787_),
    .Y(_04184_));
 sky130_fd_sc_hd__and3b_1 _45414_ (.A_N(_22787_),
    .B(_24776_),
    .C(_04173_),
    .X(_04195_));
 sky130_fd_sc_hd__o2bb2a_1 _45415_ (.A1_N(_04151_),
    .A2_N(_04162_),
    .B1(_04184_),
    .B2(_04195_),
    .X(_04206_));
 sky130_fd_sc_hd__nor2_1 _45416_ (.A(_04184_),
    .B(_04195_),
    .Y(_04217_));
 sky130_fd_sc_hd__and3_1 _45417_ (.A(_04217_),
    .B(_04162_),
    .C(_04151_),
    .X(_04228_));
 sky130_fd_sc_hd__nor2_1 _45418_ (.A(_04206_),
    .B(_04228_),
    .Y(_04239_));
 sky130_fd_sc_hd__a21oi_1 _45419_ (.A1(_04085_),
    .A2(_04107_),
    .B1(_04239_),
    .Y(_04250_));
 sky130_fd_sc_hd__and3_1 _45420_ (.A(_04107_),
    .B(_04239_),
    .C(_04085_),
    .X(_04261_));
 sky130_fd_sc_hd__nand2_1 _45421_ (.A(_00458_),
    .B(net293),
    .Y(_04272_));
 sky130_fd_sc_hd__o31ai_2 _45422_ (.A1(_00425_),
    .A2(_00436_),
    .A3(_00469_),
    .B1(_04272_),
    .Y(_04283_));
 sky130_fd_sc_hd__buf_1 _45423_ (.A(\delay_line[37][2] ),
    .X(_04294_));
 sky130_fd_sc_hd__or2b_1 _45424_ (.A(_22688_),
    .B_N(_04294_),
    .X(_04305_));
 sky130_fd_sc_hd__nand2b_1 _45425_ (.A_N(_04294_),
    .B(_22688_),
    .Y(_04316_));
 sky130_fd_sc_hd__clkbuf_2 _45426_ (.A(\delay_line[35][2] ),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_2 _45427_ (.A(_04327_),
    .X(_04338_));
 sky130_fd_sc_hd__xor2_1 _45428_ (.A(_04338_),
    .B(_00535_),
    .X(_04349_));
 sky130_fd_sc_hd__a21o_1 _45429_ (.A1(_04305_),
    .A2(_04316_),
    .B1(_04349_),
    .X(_04360_));
 sky130_fd_sc_hd__nand3_1 _45430_ (.A(_04349_),
    .B(_04305_),
    .C(_04316_),
    .Y(_04371_));
 sky130_fd_sc_hd__nand3_2 _45431_ (.A(_04360_),
    .B(net290),
    .C(_04371_),
    .Y(_04382_));
 sky130_fd_sc_hd__a21o_1 _45432_ (.A1(_04371_),
    .A2(_04360_),
    .B1(net290),
    .X(_04393_));
 sky130_fd_sc_hd__and3_1 _45433_ (.A(_04283_),
    .B(_04382_),
    .C(_04393_),
    .X(_04404_));
 sky130_fd_sc_hd__a21oi_1 _45434_ (.A1(_04382_),
    .A2(_04393_),
    .B1(_04283_),
    .Y(_04415_));
 sky130_fd_sc_hd__o22a_1 _45435_ (.A1(_04250_),
    .A2(_04261_),
    .B1(_04404_),
    .B2(_04415_),
    .X(_04426_));
 sky130_fd_sc_hd__nor4_1 _45436_ (.A(_04250_),
    .B(_04261_),
    .C(_04404_),
    .D(_04415_),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_2 _45437_ (.A(_04426_),
    .B(net91),
    .Y(_04448_));
 sky130_fd_sc_hd__a21o_1 _45438_ (.A1(_02370_),
    .A2(_02381_),
    .B1(_04448_),
    .X(_04459_));
 sky130_fd_sc_hd__nand3_1 _45439_ (.A(_04448_),
    .B(_02381_),
    .C(_02370_),
    .Y(_04470_));
 sky130_fd_sc_hd__a21oi_1 _45440_ (.A1(_04459_),
    .A2(_04470_),
    .B1(net115),
    .Y(_04481_));
 sky130_fd_sc_hd__and3_1 _45441_ (.A(_04459_),
    .B(_04470_),
    .C(net115),
    .X(_04492_));
 sky130_fd_sc_hd__nor2_1 _45442_ (.A(_04481_),
    .B(_04492_),
    .Y(_04503_));
 sky130_fd_sc_hd__xnor2_1 _45443_ (.A(_00689_),
    .B(_04503_),
    .Y(_04514_));
 sky130_fd_sc_hd__o21a_1 _45444_ (.A1(_02084_),
    .A2(_02095_),
    .B1(_04514_),
    .X(_04524_));
 sky130_fd_sc_hd__nor3_1 _45445_ (.A(_02084_),
    .B(_02095_),
    .C(_04514_),
    .Y(_04535_));
 sky130_fd_sc_hd__o221a_1 _45446_ (.A1(_23480_),
    .A2(_24754_),
    .B1(_04524_),
    .B2(_04535_),
    .C1(_00733_),
    .X(_04546_));
 sky130_fd_sc_hd__nor2_1 _45447_ (.A(_04524_),
    .B(_04535_),
    .Y(_04557_));
 sky130_fd_sc_hd__o21ai_1 _45448_ (.A1(_23469_),
    .A2(_24754_),
    .B1(_00733_),
    .Y(_04568_));
 sky130_fd_sc_hd__buf_2 _45449_ (.A(\delay_line[23][2] ),
    .X(_04579_));
 sky130_fd_sc_hd__or2_1 _45450_ (.A(\delay_line[23][1] ),
    .B(_04579_),
    .X(_04590_));
 sky130_fd_sc_hd__nand2_2 _45451_ (.A(_00370_),
    .B(_04579_),
    .Y(_04601_));
 sky130_fd_sc_hd__a21o_1 _45452_ (.A1(_04590_),
    .A2(_04601_),
    .B1(_23502_),
    .X(_04612_));
 sky130_fd_sc_hd__and2_1 _45453_ (.A(_04590_),
    .B(_04601_),
    .X(_04623_));
 sky130_fd_sc_hd__nand2_1 _45454_ (.A(_23502_),
    .B(_04623_),
    .Y(_04634_));
 sky130_fd_sc_hd__a211oi_2 _45455_ (.A1(_04612_),
    .A2(_04634_),
    .B1(_00326_),
    .C1(net93),
    .Y(_04645_));
 sky130_fd_sc_hd__o211a_2 _45456_ (.A1(_00326_),
    .A2(_00348_),
    .B1(_04612_),
    .C1(_04634_),
    .X(_04656_));
 sky130_fd_sc_hd__or3b_1 _45457_ (.A(_04645_),
    .B(_04656_),
    .C_N(_00502_),
    .X(_04667_));
 sky130_fd_sc_hd__nor2_1 _45458_ (.A(_04645_),
    .B(_04656_),
    .Y(_04678_));
 sky130_fd_sc_hd__a31o_1 _45459_ (.A1(_00480_),
    .A2(_00359_),
    .A3(_00381_),
    .B1(_04678_),
    .X(_04689_));
 sky130_fd_sc_hd__and2_1 _45460_ (.A(_04667_),
    .B(_04689_),
    .X(_04700_));
 sky130_fd_sc_hd__nand2_2 _45461_ (.A(_23633_),
    .B(_04700_),
    .Y(_04711_));
 sky130_fd_sc_hd__a21o_1 _45462_ (.A1(_23524_),
    .A2(_23622_),
    .B1(_04700_),
    .X(_04722_));
 sky130_fd_sc_hd__nand2_1 _45463_ (.A(_04711_),
    .B(_04722_),
    .Y(_04733_));
 sky130_fd_sc_hd__a21o_1 _45464_ (.A1(_04557_),
    .A2(_04568_),
    .B1(_04733_),
    .X(_04744_));
 sky130_fd_sc_hd__and2_1 _45465_ (.A(_04557_),
    .B(_04568_),
    .X(_04755_));
 sky130_fd_sc_hd__o21ai_1 _45466_ (.A1(_04546_),
    .A2(_04755_),
    .B1(_04733_),
    .Y(_04766_));
 sky130_fd_sc_hd__o21a_1 _45467_ (.A1(_04546_),
    .A2(_04744_),
    .B1(_04766_),
    .X(_04777_));
 sky130_fd_sc_hd__o21ai_1 _45468_ (.A1(_00766_),
    .A2(net75),
    .B1(_04777_),
    .Y(_04788_));
 sky130_fd_sc_hd__or3_1 _45469_ (.A(_00766_),
    .B(net75),
    .C(_04777_),
    .X(_04799_));
 sky130_fd_sc_hd__nor2_1 _45470_ (.A(net368),
    .B(net367),
    .Y(_04810_));
 sky130_fd_sc_hd__and2_1 _45471_ (.A(net368),
    .B(net367),
    .X(_04821_));
 sky130_fd_sc_hd__or3b_4 _45472_ (.A(_04810_),
    .B(_04821_),
    .C_N(_22161_),
    .X(_04832_));
 sky130_fd_sc_hd__clkbuf_2 _45473_ (.A(_04832_),
    .X(_04843_));
 sky130_fd_sc_hd__o21bai_2 _45474_ (.A1(_04810_),
    .A2(_04821_),
    .B1_N(_22161_),
    .Y(_04854_));
 sky130_fd_sc_hd__buf_2 _45475_ (.A(_04854_),
    .X(_04865_));
 sky130_fd_sc_hd__buf_1 _45476_ (.A(\delay_line[17][1] ),
    .X(_04876_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45477_ (.A(\delay_line[17][2] ),
    .X(_04887_));
 sky130_fd_sc_hd__nor2_1 _45478_ (.A(_04876_),
    .B(_04887_),
    .Y(_04898_));
 sky130_fd_sc_hd__and2_1 _45479_ (.A(\delay_line[17][1] ),
    .B(\delay_line[17][2] ),
    .X(_04909_));
 sky130_fd_sc_hd__inv_2 _45480_ (.A(_04876_),
    .Y(_04920_));
 sky130_fd_sc_hd__buf_1 _45481_ (.A(net378),
    .X(_04931_));
 sky130_fd_sc_hd__a2bb2o_1 _45482_ (.A1_N(_04898_),
    .A2_N(_04909_),
    .B1(_04920_),
    .B2(_04931_),
    .X(_04942_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45483_ (.A(_04876_),
    .X(_04953_));
 sky130_fd_sc_hd__or4_1 _45484_ (.A(_04953_),
    .B(_22139_),
    .C(_04898_),
    .D(_04909_),
    .X(_04964_));
 sky130_fd_sc_hd__and4_1 _45485_ (.A(_04843_),
    .B(_04865_),
    .C(_04942_),
    .D(_04964_),
    .X(_04975_));
 sky130_fd_sc_hd__a22oi_1 _45486_ (.A1(_04843_),
    .A2(_04865_),
    .B1(_04942_),
    .B2(_04964_),
    .Y(_04986_));
 sky130_fd_sc_hd__nor2_1 _45487_ (.A(_04975_),
    .B(_04986_),
    .Y(_04997_));
 sky130_fd_sc_hd__and3_1 _45488_ (.A(_22194_),
    .B(_04997_),
    .C(_00854_),
    .X(_05008_));
 sky130_fd_sc_hd__o2bb2a_1 _45489_ (.A1_N(_00854_),
    .A2_N(_22194_),
    .B1(_04986_),
    .B2(_04975_),
    .X(_05019_));
 sky130_fd_sc_hd__or2_1 _45490_ (.A(_05008_),
    .B(_05019_),
    .X(_05030_));
 sky130_fd_sc_hd__a21boi_1 _45491_ (.A1(_04788_),
    .A2(_04799_),
    .B1_N(_05030_),
    .Y(_05041_));
 sky130_fd_sc_hd__a41o_1 _45492_ (.A1(_23524_),
    .A2(_23480_),
    .A3(_23491_),
    .A4(_00744_),
    .B1(_00799_),
    .X(_05052_));
 sky130_fd_sc_hd__nor2_1 _45493_ (.A(_05052_),
    .B(_04777_),
    .Y(_05063_));
 sky130_fd_sc_hd__or2_1 _45494_ (.A(_05030_),
    .B(_05063_),
    .X(_05074_));
 sky130_fd_sc_hd__a21oi_1 _45495_ (.A1(_04777_),
    .A2(_05052_),
    .B1(_05074_),
    .Y(_05085_));
 sky130_fd_sc_hd__inv_2 _45496_ (.A(_00821_),
    .Y(_05096_));
 sky130_fd_sc_hd__a21oi_1 _45497_ (.A1(_05096_),
    .A2(_00865_),
    .B1(_00832_),
    .Y(_05107_));
 sky130_fd_sc_hd__o21a_1 _45498_ (.A1(_05041_),
    .A2(_05085_),
    .B1(_05107_),
    .X(_05118_));
 sky130_fd_sc_hd__nor3_1 _45499_ (.A(_05107_),
    .B(_05041_),
    .C(_05085_),
    .Y(_05129_));
 sky130_fd_sc_hd__nor2_1 _45500_ (.A(_05118_),
    .B(_05129_),
    .Y(_05140_));
 sky130_fd_sc_hd__xnor2_2 _45501_ (.A(_00919_),
    .B(_05140_),
    .Y(_00002_));
 sky130_fd_sc_hd__clkbuf_2 _45502_ (.A(_04931_),
    .X(_05161_));
 sky130_fd_sc_hd__clkbuf_2 _45503_ (.A(_04909_),
    .X(_05172_));
 sky130_fd_sc_hd__a32o_1 _45504_ (.A1(_22205_),
    .A2(_04997_),
    .A3(_00854_),
    .B1(_05161_),
    .B2(_05172_),
    .X(_05183_));
 sky130_fd_sc_hd__a211oi_1 _45505_ (.A1(_24644_),
    .A2(_24677_),
    .B1(_02293_),
    .C1(_02304_),
    .Y(_05194_));
 sky130_fd_sc_hd__inv_2 _45506_ (.A(\delay_line[32][2] ),
    .Y(_05205_));
 sky130_fd_sc_hd__clkbuf_2 _45507_ (.A(_05205_),
    .X(_05216_));
 sky130_fd_sc_hd__buf_1 _45508_ (.A(_05216_),
    .X(_05227_));
 sky130_fd_sc_hd__inv_2 _45509_ (.A(\delay_line[32][3] ),
    .Y(_05238_));
 sky130_fd_sc_hd__clkbuf_2 _45510_ (.A(_05238_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_2 _45511_ (.A(_05249_),
    .X(_05260_));
 sky130_fd_sc_hd__buf_1 _45512_ (.A(_05260_),
    .X(_05271_));
 sky130_fd_sc_hd__a31o_1 _45513_ (.A1(_24512_),
    .A2(_24545_),
    .A3(_05227_),
    .B1(_05271_),
    .X(_05282_));
 sky130_fd_sc_hd__buf_1 _45514_ (.A(\delay_line[32][3] ),
    .X(_05293_));
 sky130_fd_sc_hd__clkbuf_2 _45515_ (.A(_05293_),
    .X(_05304_));
 sky130_fd_sc_hd__buf_1 _45516_ (.A(_05304_),
    .X(_05315_));
 sky130_fd_sc_hd__or4_1 _45517_ (.A(_22567_),
    .B(_24479_),
    .C(_02128_),
    .D(_05315_),
    .X(_05326_));
 sky130_fd_sc_hd__buf_1 _45518_ (.A(net313),
    .X(_05337_));
 sky130_fd_sc_hd__buf_2 _45519_ (.A(_05337_),
    .X(_05348_));
 sky130_fd_sc_hd__a21oi_2 _45520_ (.A1(_05282_),
    .A2(_05326_),
    .B1(_05348_),
    .Y(_05359_));
 sky130_fd_sc_hd__nand2_1 _45521_ (.A(_05227_),
    .B(_05271_),
    .Y(_05370_));
 sky130_fd_sc_hd__o311a_1 _45522_ (.A1(_22567_),
    .A2(_24479_),
    .A3(_05370_),
    .B1(_05348_),
    .C1(_05282_),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_2 _45523_ (.A(\delay_line[34][3] ),
    .X(_05392_));
 sky130_fd_sc_hd__clkbuf_2 _45524_ (.A(_05392_),
    .X(_05403_));
 sky130_fd_sc_hd__xor2_2 _45525_ (.A(_00601_),
    .B(_05403_),
    .X(_05414_));
 sky130_fd_sc_hd__xnor2_2 _45526_ (.A(_02271_),
    .B(_05414_),
    .Y(_05425_));
 sky130_fd_sc_hd__nor3_1 _45527_ (.A(_05359_),
    .B(_05381_),
    .C(_05425_),
    .Y(_05436_));
 sky130_fd_sc_hd__o21a_1 _45528_ (.A1(_05359_),
    .A2(_05381_),
    .B1(_05425_),
    .X(_05447_));
 sky130_fd_sc_hd__a21boi_4 _45529_ (.A1(_01040_),
    .A2(_01051_),
    .B1_N(_01084_),
    .Y(_05458_));
 sky130_fd_sc_hd__or3b_1 _45530_ (.A(_05436_),
    .B(_05447_),
    .C_N(_05458_),
    .X(_05469_));
 sky130_fd_sc_hd__nor2_1 _45531_ (.A(_05436_),
    .B(_05447_),
    .Y(_05480_));
 sky130_fd_sc_hd__or2_1 _45532_ (.A(_05458_),
    .B(_05480_),
    .X(_05491_));
 sky130_fd_sc_hd__and2_1 _45533_ (.A(_05469_),
    .B(_05491_),
    .X(_05502_));
 sky130_fd_sc_hd__a31o_1 _45534_ (.A1(_02183_),
    .A2(_02194_),
    .A3(_02139_),
    .B1(_05502_),
    .X(_05513_));
 sky130_fd_sc_hd__o21ai_1 _45535_ (.A1(_02205_),
    .A2(_02304_),
    .B1(_05502_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21a_1 _45536_ (.A1(_02304_),
    .A2(_05513_),
    .B1(_05524_),
    .X(_05535_));
 sky130_fd_sc_hd__o21ai_2 _45537_ (.A1(_05194_),
    .A2(_02359_),
    .B1(_05535_),
    .Y(_05546_));
 sky130_fd_sc_hd__or3_1 _45538_ (.A(_05194_),
    .B(_02359_),
    .C(_05535_),
    .X(_05557_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45539_ (.A(net289),
    .X(_05568_));
 sky130_fd_sc_hd__nor2_1 _45540_ (.A(_22721_),
    .B(_05568_),
    .Y(_05579_));
 sky130_fd_sc_hd__and2_1 _45541_ (.A(\delay_line[38][0] ),
    .B(net289),
    .X(_05590_));
 sky130_fd_sc_hd__buf_1 _45542_ (.A(\delay_line[39][3] ),
    .X(_05601_));
 sky130_fd_sc_hd__buf_1 _45543_ (.A(_05601_),
    .X(_05612_));
 sky130_fd_sc_hd__buf_1 _45544_ (.A(_05612_),
    .X(_05623_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45545_ (.A(_05623_),
    .X(_05634_));
 sky130_fd_sc_hd__o31a_1 _45546_ (.A1(_22754_),
    .A2(_00403_),
    .A3(_04140_),
    .B1(_05634_),
    .X(_05645_));
 sky130_fd_sc_hd__nor4_1 _45547_ (.A(_22754_),
    .B(_00414_),
    .C(_04140_),
    .D(_05634_),
    .Y(_05656_));
 sky130_fd_sc_hd__or4_1 _45548_ (.A(_05579_),
    .B(_05590_),
    .C(_05645_),
    .D(_05656_),
    .X(_05667_));
 sky130_fd_sc_hd__o22ai_2 _45549_ (.A1(_05579_),
    .A2(_05590_),
    .B1(_05645_),
    .B2(net241),
    .Y(_05678_));
 sky130_fd_sc_hd__buf_1 _45550_ (.A(\delay_line[40][3] ),
    .X(_05689_));
 sky130_fd_sc_hd__or2_1 _45551_ (.A(_04173_),
    .B(_05689_),
    .X(_05700_));
 sky130_fd_sc_hd__nand2_1 _45552_ (.A(\delay_line[40][2] ),
    .B(\delay_line[40][3] ),
    .Y(_05711_));
 sky130_fd_sc_hd__o21a_1 _45553_ (.A1(\delay_line[40][0] ),
    .A2(_04173_),
    .B1(\delay_line[40][1] ),
    .X(_05722_));
 sky130_fd_sc_hd__and3_1 _45554_ (.A(_05700_),
    .B(_05711_),
    .C(_05722_),
    .X(_05733_));
 sky130_fd_sc_hd__a21oi_1 _45555_ (.A1(_05700_),
    .A2(_05711_),
    .B1(_05722_),
    .Y(_05744_));
 sky130_fd_sc_hd__nor2_1 _45556_ (.A(_05733_),
    .B(_05744_),
    .Y(_05755_));
 sky130_fd_sc_hd__and3_1 _45557_ (.A(_05667_),
    .B(_05678_),
    .C(_05755_),
    .X(_05766_));
 sky130_fd_sc_hd__a21oi_1 _45558_ (.A1(_05667_),
    .A2(_05678_),
    .B1(_05755_),
    .Y(_05777_));
 sky130_fd_sc_hd__nor2_2 _45559_ (.A(_05766_),
    .B(_05777_),
    .Y(_05788_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45560_ (.A(\delay_line[35][3] ),
    .X(_05799_));
 sky130_fd_sc_hd__or2_1 _45561_ (.A(\delay_line[35][2] ),
    .B(_05799_),
    .X(_05810_));
 sky130_fd_sc_hd__nand2_1 _45562_ (.A(\delay_line[35][2] ),
    .B(_05799_),
    .Y(_05821_));
 sky130_fd_sc_hd__clkbuf_2 _45563_ (.A(\delay_line[35][1] ),
    .X(_05832_));
 sky130_fd_sc_hd__nand3_1 _45564_ (.A(_05810_),
    .B(_05821_),
    .C(_05832_),
    .Y(_05843_));
 sky130_fd_sc_hd__a21o_1 _45565_ (.A1(_05810_),
    .A2(_05821_),
    .B1(_05832_),
    .X(_05854_));
 sky130_fd_sc_hd__o21ba_1 _45566_ (.A1(_04327_),
    .A2(_00546_),
    .B1_N(_00535_),
    .X(_05865_));
 sky130_fd_sc_hd__a21oi_1 _45567_ (.A1(_05843_),
    .A2(_05854_),
    .B1(_05865_),
    .Y(_05876_));
 sky130_fd_sc_hd__and3_1 _45568_ (.A(_05865_),
    .B(_05843_),
    .C(_05854_),
    .X(_05887_));
 sky130_fd_sc_hd__a2bb2o_1 _45569_ (.A1_N(_05876_),
    .A2_N(_05887_),
    .B1(_04338_),
    .B2(_00546_),
    .X(_05898_));
 sky130_fd_sc_hd__clkbuf_2 _45570_ (.A(\delay_line[35][3] ),
    .X(_05909_));
 sky130_fd_sc_hd__nand3b_1 _45571_ (.A_N(_05909_),
    .B(_00546_),
    .C(_04338_),
    .Y(_05920_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45572_ (.A(\delay_line[36][0] ),
    .X(_05931_));
 sky130_fd_sc_hd__nand3_1 _45573_ (.A(_05898_),
    .B(_05920_),
    .C(_05931_),
    .Y(_05942_));
 sky130_fd_sc_hd__inv_2 _45574_ (.A(_05942_),
    .Y(_05953_));
 sky130_fd_sc_hd__a21oi_1 _45575_ (.A1(_05898_),
    .A2(_05920_),
    .B1(_05931_),
    .Y(_05964_));
 sky130_fd_sc_hd__nand2b_1 _45576_ (.A_N(\delay_line[37][3] ),
    .B(net293),
    .Y(_05975_));
 sky130_fd_sc_hd__buf_1 _45577_ (.A(\delay_line[37][3] ),
    .X(_05986_));
 sky130_fd_sc_hd__or2b_1 _45578_ (.A(net293),
    .B_N(_05986_),
    .X(_05997_));
 sky130_fd_sc_hd__buf_1 _45579_ (.A(_05997_),
    .X(_06008_));
 sky130_fd_sc_hd__nand2_1 _45580_ (.A(_05975_),
    .B(_06008_),
    .Y(_06019_));
 sky130_fd_sc_hd__xor2_1 _45581_ (.A(_04316_),
    .B(_06019_),
    .X(_06030_));
 sky130_fd_sc_hd__o21a_1 _45582_ (.A1(_05953_),
    .A2(_05964_),
    .B1(_06030_),
    .X(_06041_));
 sky130_fd_sc_hd__nor3_1 _45583_ (.A(_06030_),
    .B(_05964_),
    .C(_05953_),
    .Y(_06052_));
 sky130_fd_sc_hd__o211a_1 _45584_ (.A1(_06041_),
    .A2(_06052_),
    .B1(_04360_),
    .C1(_04382_),
    .X(_06063_));
 sky130_fd_sc_hd__a211oi_2 _45585_ (.A1(_04360_),
    .A2(_04382_),
    .B1(_06041_),
    .C1(_06052_),
    .Y(_06073_));
 sky130_fd_sc_hd__nor3_4 _45586_ (.A(_05788_),
    .B(_06063_),
    .C(_06073_),
    .Y(_06084_));
 sky130_fd_sc_hd__o21a_2 _45587_ (.A1(_06063_),
    .A2(net156),
    .B1(_05788_),
    .X(_06095_));
 sky130_fd_sc_hd__a211o_1 _45588_ (.A1(_05546_),
    .A2(_05557_),
    .B1(_06084_),
    .C1(_06095_),
    .X(_06106_));
 sky130_fd_sc_hd__o211ai_2 _45589_ (.A1(_06084_),
    .A2(_06095_),
    .B1(_05546_),
    .C1(_05557_),
    .Y(_06117_));
 sky130_fd_sc_hd__o211a_1 _45590_ (.A1(_01326_),
    .A2(_01359_),
    .B1(_06106_),
    .C1(_06117_),
    .X(_06128_));
 sky130_fd_sc_hd__a211oi_1 _45591_ (.A1(_06106_),
    .A2(_06117_),
    .B1(_01326_),
    .C1(_01359_),
    .Y(_06139_));
 sky130_fd_sc_hd__o211ai_1 _45592_ (.A1(_06128_),
    .A2(_06139_),
    .B1(_02370_),
    .C1(_04470_),
    .Y(_06150_));
 sky130_fd_sc_hd__inv_2 _45593_ (.A(_06150_),
    .Y(_06161_));
 sky130_fd_sc_hd__a211oi_1 _45594_ (.A1(_02370_),
    .A2(_04470_),
    .B1(_06128_),
    .C1(_06139_),
    .Y(_06172_));
 sky130_fd_sc_hd__buf_1 _45595_ (.A(_06172_),
    .X(_06183_));
 sky130_fd_sc_hd__o21ba_4 _45596_ (.A1(_01095_),
    .A2(_01282_),
    .B1_N(_01293_),
    .X(_06194_));
 sky130_fd_sc_hd__buf_1 _45597_ (.A(\delay_line[31][3] ),
    .X(_06205_));
 sky130_fd_sc_hd__buf_2 _45598_ (.A(_06205_),
    .X(_06216_));
 sky130_fd_sc_hd__o211a_1 _45599_ (.A1(_24589_),
    .A2(_00985_),
    .B1(_06216_),
    .C1(_22237_),
    .X(_06227_));
 sky130_fd_sc_hd__nor2_1 _45600_ (.A(_24589_),
    .B(_00985_),
    .Y(_06238_));
 sky130_fd_sc_hd__inv_2 _45601_ (.A(\delay_line[31][3] ),
    .Y(_06249_));
 sky130_fd_sc_hd__buf_1 _45602_ (.A(_06249_),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_2 _45603_ (.A(_06260_),
    .X(_06271_));
 sky130_fd_sc_hd__o21a_1 _45604_ (.A1(_24567_),
    .A2(_06238_),
    .B1(_06271_),
    .X(_06282_));
 sky130_fd_sc_hd__buf_1 _45605_ (.A(\delay_line[30][3] ),
    .X(_06293_));
 sky130_fd_sc_hd__buf_1 _45606_ (.A(_06293_),
    .X(_06304_));
 sky130_fd_sc_hd__clkbuf_2 _45607_ (.A(_06304_),
    .X(_06315_));
 sky130_fd_sc_hd__clkbuf_2 _45608_ (.A(_06315_),
    .X(_06326_));
 sky130_fd_sc_hd__clkbuf_2 _45609_ (.A(_06326_),
    .X(_06337_));
 sky130_fd_sc_hd__and2_1 _45610_ (.A(_22303_),
    .B(_06337_),
    .X(_06348_));
 sky130_fd_sc_hd__nor2_2 _45611_ (.A(_22303_),
    .B(_06337_),
    .Y(_06359_));
 sky130_fd_sc_hd__or3b_2 _45612_ (.A(_06348_),
    .B(_06359_),
    .C_N(net323),
    .X(_06370_));
 sky130_fd_sc_hd__o21bai_2 _45613_ (.A1(_06348_),
    .A2(_06359_),
    .B1_N(net323),
    .Y(_06381_));
 sky130_fd_sc_hd__and4bb_4 _45614_ (.A_N(_06227_),
    .B_N(_06282_),
    .C(_06370_),
    .D(_06381_),
    .X(_06392_));
 sky130_fd_sc_hd__a2bb2oi_4 _45615_ (.A1_N(_06227_),
    .A2_N(_06282_),
    .B1(_06370_),
    .B2(_06381_),
    .Y(_06403_));
 sky130_fd_sc_hd__buf_1 _45616_ (.A(net328),
    .X(_06414_));
 sky130_fd_sc_hd__clkbuf_2 _45617_ (.A(_06414_),
    .X(_06425_));
 sky130_fd_sc_hd__nand2_1 _45618_ (.A(_22248_),
    .B(_24369_),
    .Y(_06436_));
 sky130_fd_sc_hd__mux2_1 _45619_ (.A0(_06436_),
    .A1(_24380_),
    .S(_01128_),
    .X(_06447_));
 sky130_fd_sc_hd__xor2_2 _45620_ (.A(_06425_),
    .B(_06447_),
    .X(_06458_));
 sky130_fd_sc_hd__inv_2 _45621_ (.A(net339),
    .Y(_06469_));
 sky130_fd_sc_hd__buf_2 _45622_ (.A(_06469_),
    .X(_06480_));
 sky130_fd_sc_hd__buf_1 _45623_ (.A(\delay_line[27][3] ),
    .X(_06491_));
 sky130_fd_sc_hd__nor2_1 _45624_ (.A(_24303_),
    .B(_06491_),
    .Y(_06502_));
 sky130_fd_sc_hd__nand2_1 _45625_ (.A(_24303_),
    .B(_06491_),
    .Y(_06513_));
 sky130_fd_sc_hd__and4b_1 _45626_ (.A_N(_06502_),
    .B(_01183_),
    .C(_22468_),
    .D(_06513_),
    .X(_06524_));
 sky130_fd_sc_hd__and2_1 _45627_ (.A(\delay_line[27][1] ),
    .B(_06491_),
    .X(_06535_));
 sky130_fd_sc_hd__o2bb2ai_1 _45628_ (.A1_N(_22457_),
    .A2_N(_01183_),
    .B1(_06535_),
    .B2(_06502_),
    .Y(_06546_));
 sky130_fd_sc_hd__or3b_2 _45629_ (.A(_06480_),
    .B(_06524_),
    .C_N(_06546_),
    .X(_06557_));
 sky130_fd_sc_hd__nand4b_1 _45630_ (.A_N(_06502_),
    .B(_01183_),
    .C(_22457_),
    .D(_06513_),
    .Y(_06568_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45631_ (.A(_06568_),
    .X(_06579_));
 sky130_fd_sc_hd__buf_2 _45632_ (.A(net339),
    .X(_06590_));
 sky130_fd_sc_hd__a21o_1 _45633_ (.A1(_06579_),
    .A2(_06546_),
    .B1(_06590_),
    .X(_06601_));
 sky130_fd_sc_hd__nand3b_4 _45634_ (.A_N(_06458_),
    .B(_06557_),
    .C(_06601_),
    .Y(_06612_));
 sky130_fd_sc_hd__a21bo_1 _45635_ (.A1(_06557_),
    .A2(_06601_),
    .B1_N(_06458_),
    .X(_06623_));
 sky130_fd_sc_hd__a21o_1 _45636_ (.A1(_01172_),
    .A2(_01205_),
    .B1(_01238_),
    .X(_06634_));
 sky130_fd_sc_hd__a21oi_4 _45637_ (.A1(_06612_),
    .A2(_06623_),
    .B1(_06634_),
    .Y(_06645_));
 sky130_fd_sc_hd__and3_4 _45638_ (.A(_06634_),
    .B(_06612_),
    .C(_06623_),
    .X(_06656_));
 sky130_fd_sc_hd__o22ai_1 _45639_ (.A1(_06392_),
    .A2(_06403_),
    .B1(_06645_),
    .B2(_06656_),
    .Y(_06667_));
 sky130_fd_sc_hd__or4_1 _45640_ (.A(_06392_),
    .B(_06403_),
    .C(_06645_),
    .D(_06656_),
    .X(_06678_));
 sky130_fd_sc_hd__a211oi_1 _45641_ (.A1(_23720_),
    .A2(_23786_),
    .B1(_01545_),
    .C1(_01556_),
    .Y(_06689_));
 sky130_fd_sc_hd__a211o_1 _45642_ (.A1(_06667_),
    .A2(_06678_),
    .B1(_01545_),
    .C1(_06689_),
    .X(_06700_));
 sky130_fd_sc_hd__o211ai_1 _45643_ (.A1(_01545_),
    .A2(_06689_),
    .B1(_06667_),
    .C1(_06678_),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_1 _45644_ (.A(_06700_),
    .B(_06711_),
    .Y(_06722_));
 sky130_fd_sc_hd__xnor2_1 _45645_ (.A(_06194_),
    .B(_06722_),
    .Y(_06733_));
 sky130_fd_sc_hd__a21bo_2 _45646_ (.A1(_01424_),
    .A2(_01457_),
    .B1_N(_01523_),
    .X(_06744_));
 sky130_fd_sc_hd__inv_2 _45647_ (.A(\delay_line[25][1] ),
    .Y(_06755_));
 sky130_fd_sc_hd__buf_1 _45648_ (.A(\delay_line[25][3] ),
    .X(_06766_));
 sky130_fd_sc_hd__and2_2 _45649_ (.A(_06755_),
    .B(_06766_),
    .X(_06777_));
 sky130_fd_sc_hd__buf_1 _45650_ (.A(_06766_),
    .X(_06788_));
 sky130_fd_sc_hd__clkbuf_2 _45651_ (.A(_06788_),
    .X(_06799_));
 sky130_fd_sc_hd__buf_1 _45652_ (.A(_06755_),
    .X(_06810_));
 sky130_fd_sc_hd__buf_2 _45653_ (.A(_06810_),
    .X(_06821_));
 sky130_fd_sc_hd__nor2_2 _45654_ (.A(_06799_),
    .B(_06821_),
    .Y(_06832_));
 sky130_fd_sc_hd__or3_2 _45655_ (.A(_01512_),
    .B(_06777_),
    .C(_06832_),
    .X(_06843_));
 sky130_fd_sc_hd__o21ai_4 _45656_ (.A1(_06777_),
    .A2(_06832_),
    .B1(_01512_),
    .Y(_06854_));
 sky130_fd_sc_hd__clkbuf_2 _45657_ (.A(net355),
    .X(_06865_));
 sky130_fd_sc_hd__clkbuf_2 _45658_ (.A(_06865_),
    .X(_06876_));
 sky130_fd_sc_hd__clkbuf_2 _45659_ (.A(_06876_),
    .X(_06887_));
 sky130_fd_sc_hd__buf_1 _45660_ (.A(\delay_line[24][2] ),
    .X(_06898_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45661_ (.A(_06898_),
    .X(_06909_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45662_ (.A(_06909_),
    .X(_06920_));
 sky130_fd_sc_hd__clkbuf_4 _45663_ (.A(_06920_),
    .X(_06931_));
 sky130_fd_sc_hd__nand2_1 _45664_ (.A(_06887_),
    .B(_06931_),
    .Y(_06942_));
 sky130_fd_sc_hd__or2_1 _45665_ (.A(_06887_),
    .B(_06931_),
    .X(_06953_));
 sky130_fd_sc_hd__a22o_2 _45666_ (.A1(_06843_),
    .A2(_06854_),
    .B1(_06942_),
    .B2(_06953_),
    .X(_06964_));
 sky130_fd_sc_hd__nor2_1 _45667_ (.A(_06887_),
    .B(_06931_),
    .Y(_06975_));
 sky130_fd_sc_hd__nand2_1 _45668_ (.A(_06843_),
    .B(_06854_),
    .Y(_06986_));
 sky130_fd_sc_hd__or3b_2 _45669_ (.A(_06975_),
    .B(_06986_),
    .C_N(_06942_),
    .X(_06997_));
 sky130_fd_sc_hd__o211ai_4 _45670_ (.A1(_01699_),
    .A2(_01732_),
    .B1(_06964_),
    .C1(_06997_),
    .Y(_07008_));
 sky130_fd_sc_hd__a221o_1 _45671_ (.A1(_01710_),
    .A2(_01688_),
    .B1(_06997_),
    .B2(_06964_),
    .C1(_01732_),
    .X(_07019_));
 sky130_fd_sc_hd__and3_1 _45672_ (.A(_06744_),
    .B(_07008_),
    .C(_07019_),
    .X(_07030_));
 sky130_fd_sc_hd__a21oi_1 _45673_ (.A1(_07008_),
    .A2(_07019_),
    .B1(_06744_),
    .Y(_07041_));
 sky130_fd_sc_hd__or2_1 _45674_ (.A(_07030_),
    .B(_07041_),
    .X(_07052_));
 sky130_fd_sc_hd__inv_2 _45675_ (.A(\delay_line[15][1] ),
    .Y(_07063_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45676_ (.A(\delay_line[15][3] ),
    .X(_07074_));
 sky130_fd_sc_hd__and2_1 _45677_ (.A(_07063_),
    .B(_07074_),
    .X(_07085_));
 sky130_fd_sc_hd__buf_1 _45678_ (.A(_07074_),
    .X(_07096_));
 sky130_fd_sc_hd__buf_1 _45679_ (.A(_07096_),
    .X(_07107_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45680_ (.A(_07063_),
    .X(_07118_));
 sky130_fd_sc_hd__nor2_1 _45681_ (.A(_07107_),
    .B(_07118_),
    .Y(_07129_));
 sky130_fd_sc_hd__o21ai_1 _45682_ (.A1(_07085_),
    .A2(_07129_),
    .B1(_01809_),
    .Y(_07140_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45683_ (.A(_07140_),
    .X(_07151_));
 sky130_fd_sc_hd__or3_1 _45684_ (.A(_01809_),
    .B(_07085_),
    .C(_07129_),
    .X(_07162_));
 sky130_fd_sc_hd__buf_1 _45685_ (.A(\delay_line[14][2] ),
    .X(_07173_));
 sky130_fd_sc_hd__clkbuf_2 _45686_ (.A(_07173_),
    .X(_07184_));
 sky130_fd_sc_hd__a21oi_1 _45687_ (.A1(_07151_),
    .A2(_07162_),
    .B1(_07184_),
    .Y(_07195_));
 sky130_fd_sc_hd__clkbuf_2 _45688_ (.A(\delay_line[16][2] ),
    .X(_07206_));
 sky130_fd_sc_hd__inv_2 _45689_ (.A(_07206_),
    .Y(_07217_));
 sky130_fd_sc_hd__and3_1 _45690_ (.A(_07162_),
    .B(_07184_),
    .C(_07151_),
    .X(_07228_));
 sky130_fd_sc_hd__nor3_1 _45691_ (.A(_07195_),
    .B(_07217_),
    .C(_07228_),
    .Y(_07239_));
 sky130_fd_sc_hd__o21a_1 _45692_ (.A1(_07228_),
    .A2(_07195_),
    .B1(_07217_),
    .X(_07250_));
 sky130_fd_sc_hd__a21oi_1 _45693_ (.A1(_01776_),
    .A2(_01842_),
    .B1(_01908_),
    .Y(_07261_));
 sky130_fd_sc_hd__o21a_2 _45694_ (.A1(_07239_),
    .A2(_07250_),
    .B1(_07261_),
    .X(_07272_));
 sky130_fd_sc_hd__nor3_1 _45695_ (.A(_07261_),
    .B(_07239_),
    .C(_07250_),
    .Y(_07283_));
 sky130_fd_sc_hd__clkbuf_2 _45696_ (.A(_01600_),
    .X(_07294_));
 sky130_fd_sc_hd__buf_1 _45697_ (.A(net361),
    .X(_07305_));
 sky130_fd_sc_hd__clkbuf_2 _45698_ (.A(_07305_),
    .X(_07316_));
 sky130_fd_sc_hd__xor2_2 _45699_ (.A(_07294_),
    .B(_07316_),
    .X(_07327_));
 sky130_fd_sc_hd__clkbuf_2 _45700_ (.A(_23984_),
    .X(_07338_));
 sky130_fd_sc_hd__nand2_1 _45701_ (.A(_07338_),
    .B(_07294_),
    .Y(_07349_));
 sky130_fd_sc_hd__buf_1 _45702_ (.A(\delay_line[19][1] ),
    .X(_07360_));
 sky130_fd_sc_hd__clkbuf_2 _45703_ (.A(_07360_),
    .X(_07371_));
 sky130_fd_sc_hd__buf_1 _45704_ (.A(\delay_line[19][2] ),
    .X(_07382_));
 sky130_fd_sc_hd__buf_2 _45705_ (.A(_07382_),
    .X(_07393_));
 sky130_fd_sc_hd__xor2_2 _45706_ (.A(_07371_),
    .B(_07393_),
    .X(_07404_));
 sky130_fd_sc_hd__buf_1 _45707_ (.A(_07371_),
    .X(_07415_));
 sky130_fd_sc_hd__clkbuf_2 _45708_ (.A(_07415_),
    .X(_07426_));
 sky130_fd_sc_hd__nand2_1 _45709_ (.A(_23907_),
    .B(_07426_),
    .Y(_07437_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45710_ (.A(_07382_),
    .X(_07448_));
 sky130_fd_sc_hd__buf_1 _45711_ (.A(_07448_),
    .X(_07459_));
 sky130_fd_sc_hd__buf_1 _45712_ (.A(_07459_),
    .X(_07470_));
 sky130_fd_sc_hd__and3_1 _45713_ (.A(_23896_),
    .B(_07415_),
    .C(_07470_),
    .X(_07481_));
 sky130_fd_sc_hd__buf_1 _45714_ (.A(_07481_),
    .X(_07492_));
 sky130_fd_sc_hd__a21o_1 _45715_ (.A1(_07404_),
    .A2(_07437_),
    .B1(_07492_),
    .X(_07503_));
 sky130_fd_sc_hd__buf_2 _45716_ (.A(net374),
    .X(_07514_));
 sky130_fd_sc_hd__clkbuf_2 _45717_ (.A(_07514_),
    .X(_07525_));
 sky130_fd_sc_hd__clkbuf_2 _45718_ (.A(_07525_),
    .X(_07536_));
 sky130_fd_sc_hd__nand2_4 _45719_ (.A(_07503_),
    .B(_07536_),
    .Y(_07547_));
 sky130_fd_sc_hd__a211o_2 _45720_ (.A1(_07404_),
    .A2(_07437_),
    .B1(_07536_),
    .C1(_07492_),
    .X(_07558_));
 sky130_fd_sc_hd__buf_1 _45721_ (.A(_07294_),
    .X(_07569_));
 sky130_fd_sc_hd__buf_1 _45722_ (.A(_07316_),
    .X(_07580_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45723_ (.A(_07580_),
    .X(_07591_));
 sky130_fd_sc_hd__clkbuf_2 _45724_ (.A(_07591_),
    .X(_07602_));
 sky130_fd_sc_hd__and3_1 _45725_ (.A(_24006_),
    .B(_07569_),
    .C(_07602_),
    .X(_07613_));
 sky130_fd_sc_hd__a221o_1 _45726_ (.A1(_07327_),
    .A2(_07349_),
    .B1(_07547_),
    .B2(_07558_),
    .C1(_07613_),
    .X(_07624_));
 sky130_fd_sc_hd__a21oi_1 _45727_ (.A1(_07327_),
    .A2(_07349_),
    .B1(_07613_),
    .Y(_07635_));
 sky130_fd_sc_hd__nand3b_4 _45728_ (.A_N(_07635_),
    .B(_07558_),
    .C(_07547_),
    .Y(_07645_));
 sky130_fd_sc_hd__and2_1 _45729_ (.A(_07624_),
    .B(_07645_),
    .X(_07656_));
 sky130_fd_sc_hd__or3b_1 _45730_ (.A(_07272_),
    .B(net148),
    .C_N(_07656_),
    .X(_07667_));
 sky130_fd_sc_hd__nor2_1 _45731_ (.A(_07272_),
    .B(net148),
    .Y(_07678_));
 sky130_fd_sc_hd__or2_1 _45732_ (.A(_07656_),
    .B(_07678_),
    .X(_07689_));
 sky130_fd_sc_hd__a211oi_2 _45733_ (.A1(_24116_),
    .A2(_24160_),
    .B1(_01908_),
    .C1(_01919_),
    .Y(_07700_));
 sky130_fd_sc_hd__a211oi_2 _45734_ (.A1(_07667_),
    .A2(_07689_),
    .B1(_07700_),
    .C1(_01952_),
    .Y(_07711_));
 sky130_fd_sc_hd__o211ai_2 _45735_ (.A1(_07700_),
    .A2(_01952_),
    .B1(_07667_),
    .C1(_07689_),
    .Y(_07722_));
 sky130_fd_sc_hd__or2b_1 _45736_ (.A(_07711_),
    .B_N(_07722_),
    .X(_07733_));
 sky130_fd_sc_hd__xor2_1 _45737_ (.A(_07052_),
    .B(_07733_),
    .X(_07744_));
 sky130_fd_sc_hd__a211oi_1 _45738_ (.A1(_24171_),
    .A2(_24193_),
    .B1(_01952_),
    .C1(_01963_),
    .Y(_07755_));
 sky130_fd_sc_hd__a311o_1 _45739_ (.A1(_01567_),
    .A2(_01578_),
    .A3(_01985_),
    .B1(_07744_),
    .C1(_07755_),
    .X(_07766_));
 sky130_fd_sc_hd__o21ai_1 _45740_ (.A1(_07755_),
    .A2(_01996_),
    .B1(_07744_),
    .Y(_07777_));
 sky130_fd_sc_hd__nand2_1 _45741_ (.A(_07766_),
    .B(_07777_),
    .Y(_07788_));
 sky130_fd_sc_hd__xnor2_1 _45742_ (.A(_06733_),
    .B(_07788_),
    .Y(_07799_));
 sky130_fd_sc_hd__a21oi_1 _45743_ (.A1(_01381_),
    .A2(_02051_),
    .B1(_02040_),
    .Y(_07810_));
 sky130_fd_sc_hd__xnor2_1 _45744_ (.A(_07799_),
    .B(_07810_),
    .Y(_07821_));
 sky130_fd_sc_hd__o21ai_1 _45745_ (.A1(_06161_),
    .A2(_06183_),
    .B1(_07821_),
    .Y(_07832_));
 sky130_fd_sc_hd__or3_1 _45746_ (.A(_07821_),
    .B(_06161_),
    .C(_06172_),
    .X(_07843_));
 sky130_fd_sc_hd__and2_1 _45747_ (.A(_07832_),
    .B(_07843_),
    .X(_07854_));
 sky130_fd_sc_hd__o21a_1 _45748_ (.A1(_02084_),
    .A2(_04535_),
    .B1(_07854_),
    .X(_07865_));
 sky130_fd_sc_hd__o21ai_1 _45749_ (.A1(_02095_),
    .A2(_04514_),
    .B1(_02073_),
    .Y(_07876_));
 sky130_fd_sc_hd__nor2_1 _45750_ (.A(_07854_),
    .B(_07876_),
    .Y(_07887_));
 sky130_fd_sc_hd__or2_1 _45751_ (.A(_07865_),
    .B(_07887_),
    .X(_07898_));
 sky130_fd_sc_hd__buf_2 _45752_ (.A(_00370_),
    .X(_07909_));
 sky130_fd_sc_hd__nand2_1 _45753_ (.A(_03062_),
    .B(_03381_),
    .Y(_07920_));
 sky130_fd_sc_hd__o22a_1 _45754_ (.A1(_02744_),
    .A2(_02810_),
    .B1(_03040_),
    .B2(_03018_),
    .X(_07931_));
 sky130_fd_sc_hd__a21oi_1 _45755_ (.A1(_02612_),
    .A2(_02645_),
    .B1(_25270_),
    .Y(_07942_));
 sky130_fd_sc_hd__a21oi_2 _45756_ (.A1(_02590_),
    .A2(_02568_),
    .B1(_23150_),
    .Y(_07953_));
 sky130_fd_sc_hd__nor2_1 _45757_ (.A(_25237_),
    .B(_07953_),
    .Y(_07964_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45758_ (.A(\delay_line[4][0] ),
    .X(_07975_));
 sky130_fd_sc_hd__clkbuf_2 _45759_ (.A(\delay_line[11][1] ),
    .X(_07986_));
 sky130_fd_sc_hd__and2_1 _45760_ (.A(_07975_),
    .B(_07986_),
    .X(_07997_));
 sky130_fd_sc_hd__clkbuf_4 _45761_ (.A(_07997_),
    .X(_08008_));
 sky130_fd_sc_hd__clkbuf_2 _45762_ (.A(_07986_),
    .X(_08019_));
 sky130_fd_sc_hd__o21ai_1 _45763_ (.A1(_07975_),
    .A2(_08019_),
    .B1(\delay_line[0][3] ),
    .Y(_08030_));
 sky130_fd_sc_hd__clkbuf_2 _45764_ (.A(_08030_),
    .X(_08041_));
 sky130_fd_sc_hd__clkbuf_2 _45765_ (.A(_07975_),
    .X(_08052_));
 sky130_fd_sc_hd__nor2_1 _45766_ (.A(_08052_),
    .B(_08019_),
    .Y(_08063_));
 sky130_fd_sc_hd__clkbuf_2 _45767_ (.A(\delay_line[0][3] ),
    .X(_08074_));
 sky130_fd_sc_hd__inv_2 _45768_ (.A(_08074_),
    .Y(_08085_));
 sky130_fd_sc_hd__o21ai_4 _45769_ (.A1(_08008_),
    .A2(_08063_),
    .B1(_08085_),
    .Y(_08096_));
 sky130_fd_sc_hd__o211ai_1 _45770_ (.A1(_08008_),
    .A2(_08041_),
    .B1(_02546_),
    .C1(_08096_),
    .Y(_08107_));
 sky130_fd_sc_hd__buf_2 _45771_ (.A(_02524_),
    .X(_08118_));
 sky130_fd_sc_hd__inv_2 _45772_ (.A(\delay_line[4][0] ),
    .Y(_08129_));
 sky130_fd_sc_hd__clkbuf_2 _45773_ (.A(_08129_),
    .X(_08140_));
 sky130_fd_sc_hd__inv_2 _45774_ (.A(_07986_),
    .Y(_08151_));
 sky130_fd_sc_hd__o21ai_2 _45775_ (.A1(_08140_),
    .A2(_08151_),
    .B1(_08041_),
    .Y(_08162_));
 sky130_fd_sc_hd__o21ai_1 _45776_ (.A1(_08041_),
    .A2(_08008_),
    .B1(_08074_),
    .Y(_08173_));
 sky130_fd_sc_hd__o221ai_2 _45777_ (.A1(_08118_),
    .A2(_02579_),
    .B1(_08063_),
    .B2(_08162_),
    .C1(_08173_),
    .Y(_08184_));
 sky130_fd_sc_hd__nand3_2 _45778_ (.A(_07964_),
    .B(_08107_),
    .C(_08184_),
    .Y(_08195_));
 sky130_fd_sc_hd__nand2_1 _45779_ (.A(_08052_),
    .B(_08019_),
    .Y(_08206_));
 sky130_fd_sc_hd__nand2_1 _45780_ (.A(_08140_),
    .B(_08151_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand3_1 _45781_ (.A(_08206_),
    .B(_08217_),
    .C(_08041_),
    .Y(_08228_));
 sky130_fd_sc_hd__nand3_1 _45782_ (.A(_08173_),
    .B(_08228_),
    .C(_02546_),
    .Y(_08239_));
 sky130_fd_sc_hd__o221ai_4 _45783_ (.A1(_08118_),
    .A2(_02579_),
    .B1(_08008_),
    .B2(_08041_),
    .C1(_08096_),
    .Y(_08250_));
 sky130_fd_sc_hd__o211ai_4 _45784_ (.A1(_25237_),
    .A2(_07953_),
    .B1(_08239_),
    .C1(_08250_),
    .Y(_08261_));
 sky130_fd_sc_hd__clkbuf_2 _45785_ (.A(\delay_line[13][3] ),
    .X(_08272_));
 sky130_fd_sc_hd__a21oi_2 _45786_ (.A1(_08195_),
    .A2(_08261_),
    .B1(_08272_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand3_2 _45787_ (.A(_08195_),
    .B(_08261_),
    .C(\delay_line[13][3] ),
    .Y(_08294_));
 sky130_fd_sc_hd__and3_1 _45788_ (.A(_02623_),
    .B(_02634_),
    .C(_02480_),
    .X(_08305_));
 sky130_fd_sc_hd__nand2_1 _45789_ (.A(_08294_),
    .B(_08305_),
    .Y(_08316_));
 sky130_fd_sc_hd__nand2_1 _45790_ (.A(_02623_),
    .B(_02634_),
    .Y(_08327_));
 sky130_fd_sc_hd__a21o_1 _45791_ (.A1(_08195_),
    .A2(_08261_),
    .B1(\delay_line[13][3] ),
    .X(_08338_));
 sky130_fd_sc_hd__a2bb2o_1 _45792_ (.A1_N(_02491_),
    .A2_N(_08327_),
    .B1(_08294_),
    .B2(_08338_),
    .X(_08349_));
 sky130_fd_sc_hd__o211ai_4 _45793_ (.A1(_08283_),
    .A2(_08316_),
    .B1(_25194_),
    .C1(_08349_),
    .Y(_08360_));
 sky130_fd_sc_hd__nor2_2 _45794_ (.A(_08283_),
    .B(_08316_),
    .Y(_08371_));
 sky130_fd_sc_hd__a2bb2oi_1 _45795_ (.A1_N(_02491_),
    .A2_N(_08327_),
    .B1(_08294_),
    .B2(_08338_),
    .Y(_08382_));
 sky130_fd_sc_hd__buf_2 _45796_ (.A(_25215_),
    .X(_08393_));
 sky130_fd_sc_hd__o21ai_2 _45797_ (.A1(_08371_),
    .A2(_08382_),
    .B1(_08393_),
    .Y(_08404_));
 sky130_fd_sc_hd__a21oi_1 _45798_ (.A1(_02689_),
    .A2(_02678_),
    .B1(_02755_),
    .Y(_08415_));
 sky130_fd_sc_hd__a21o_1 _45799_ (.A1(_08360_),
    .A2(_08404_),
    .B1(_08415_),
    .X(_08426_));
 sky130_fd_sc_hd__buf_1 _45800_ (.A(_02425_),
    .X(_08437_));
 sky130_fd_sc_hd__and3b_1 _45801_ (.A_N(_08437_),
    .B(_25292_),
    .C(_23227_),
    .X(_08448_));
 sky130_fd_sc_hd__and2_1 _45802_ (.A(_02447_),
    .B(_08437_),
    .X(_08459_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45803_ (.A(net407),
    .X(_08470_));
 sky130_fd_sc_hd__clkbuf_2 _45804_ (.A(_08470_),
    .X(_08481_));
 sky130_fd_sc_hd__o21a_1 _45805_ (.A1(_08448_),
    .A2(_08459_),
    .B1(_08481_),
    .X(_08492_));
 sky130_fd_sc_hd__a211oi_2 _45806_ (.A1(_02447_),
    .A2(_08437_),
    .B1(_08481_),
    .C1(_08448_),
    .Y(_08503_));
 sky130_fd_sc_hd__nor2_1 _45807_ (.A(_08492_),
    .B(_08503_),
    .Y(_08514_));
 sky130_fd_sc_hd__clkbuf_2 _45808_ (.A(net398),
    .X(_08525_));
 sky130_fd_sc_hd__o2111ai_4 _45809_ (.A1(_08525_),
    .A2(_02766_),
    .B1(_08360_),
    .C1(_08404_),
    .D1(_02667_),
    .Y(_08536_));
 sky130_fd_sc_hd__nand3_1 _45810_ (.A(_08426_),
    .B(_08514_),
    .C(_08536_),
    .Y(_08547_));
 sky130_fd_sc_hd__a31o_1 _45811_ (.A1(_08338_),
    .A2(_08305_),
    .A3(_08294_),
    .B1(_08393_),
    .X(_08558_));
 sky130_fd_sc_hd__o211a_1 _45812_ (.A1(_08382_),
    .A2(_08558_),
    .B1(_08415_),
    .C1(_08404_),
    .X(_08569_));
 sky130_fd_sc_hd__a21oi_1 _45813_ (.A1(_08360_),
    .A2(_08404_),
    .B1(_08415_),
    .Y(_08580_));
 sky130_fd_sc_hd__o22ai_1 _45814_ (.A1(_08492_),
    .A2(_08503_),
    .B1(_08569_),
    .B2(_08580_),
    .Y(_08591_));
 sky130_fd_sc_hd__o211ai_1 _45815_ (.A1(_02744_),
    .A2(_07942_),
    .B1(_08547_),
    .C1(_08591_),
    .Y(_08602_));
 sky130_fd_sc_hd__o21ai_1 _45816_ (.A1(_08569_),
    .A2(_08580_),
    .B1(_08514_),
    .Y(_08613_));
 sky130_fd_sc_hd__o211ai_1 _45817_ (.A1(_08492_),
    .A2(_08503_),
    .B1(_08536_),
    .C1(_08426_),
    .Y(_08624_));
 sky130_fd_sc_hd__nor2_1 _45818_ (.A(_02744_),
    .B(_07942_),
    .Y(_08635_));
 sky130_fd_sc_hd__nand3_1 _45819_ (.A(_08613_),
    .B(_08624_),
    .C(_08635_),
    .Y(_08646_));
 sky130_fd_sc_hd__buf_2 _45820_ (.A(net422),
    .X(_08657_));
 sky130_fd_sc_hd__clkbuf_2 _45821_ (.A(_08657_),
    .X(_08668_));
 sky130_fd_sc_hd__nor2_1 _45822_ (.A(_23106_),
    .B(_08668_),
    .Y(_08679_));
 sky130_fd_sc_hd__and2_1 _45823_ (.A(net415),
    .B(_08657_),
    .X(_08690_));
 sky130_fd_sc_hd__buf_1 _45824_ (.A(\delay_line[10][3] ),
    .X(_08701_));
 sky130_fd_sc_hd__clkbuf_2 _45825_ (.A(_08701_),
    .X(_08712_));
 sky130_fd_sc_hd__clkbuf_2 _45826_ (.A(_08712_),
    .X(_08723_));
 sky130_fd_sc_hd__or3b_1 _45827_ (.A(_08679_),
    .B(_08690_),
    .C_N(_08723_),
    .X(_08734_));
 sky130_fd_sc_hd__nor2_1 _45828_ (.A(_08679_),
    .B(_08690_),
    .Y(_08745_));
 sky130_fd_sc_hd__or2_1 _45829_ (.A(_08723_),
    .B(_08745_),
    .X(_08756_));
 sky130_fd_sc_hd__o2111a_2 _45830_ (.A1(_02865_),
    .A2(_02887_),
    .B1(_02832_),
    .C1(_08734_),
    .D1(_08756_),
    .X(_08767_));
 sky130_fd_sc_hd__a21boi_2 _45831_ (.A1(_08734_),
    .A2(_08756_),
    .B1_N(_02909_),
    .Y(_08778_));
 sky130_fd_sc_hd__o2bb2ai_1 _45832_ (.A1_N(_08602_),
    .A2_N(_08646_),
    .B1(_08767_),
    .B2(_08778_),
    .Y(_08789_));
 sky130_fd_sc_hd__or2_1 _45833_ (.A(_08767_),
    .B(_08778_),
    .X(_08800_));
 sky130_fd_sc_hd__buf_1 _45834_ (.A(_08602_),
    .X(_08811_));
 sky130_fd_sc_hd__nand3b_1 _45835_ (.A_N(_08800_),
    .B(_08646_),
    .C(_08811_),
    .Y(_08822_));
 sky130_fd_sc_hd__nand3b_2 _45836_ (.A_N(_07931_),
    .B(_08789_),
    .C(_08822_),
    .Y(_08833_));
 sky130_fd_sc_hd__a21o_1 _45837_ (.A1(_08811_),
    .A2(_08646_),
    .B1(_08800_),
    .X(_08844_));
 sky130_fd_sc_hd__o211ai_1 _45838_ (.A1(_08767_),
    .A2(_08778_),
    .B1(_08811_),
    .C1(_08646_),
    .Y(_08855_));
 sky130_fd_sc_hd__nand3_2 _45839_ (.A(_08844_),
    .B(_07931_),
    .C(_08855_),
    .Y(_08866_));
 sky130_fd_sc_hd__clkbuf_2 _45840_ (.A(_25073_),
    .X(_08877_));
 sky130_fd_sc_hd__nor2_1 _45841_ (.A(_23084_),
    .B(_02854_),
    .Y(_08888_));
 sky130_fd_sc_hd__nor2b_2 _45842_ (.A(\delay_line[9][1] ),
    .B_N(_02843_),
    .Y(_08899_));
 sky130_fd_sc_hd__a21oi_1 _45843_ (.A1(_08877_),
    .A2(_08888_),
    .B1(_08899_),
    .Y(_08910_));
 sky130_fd_sc_hd__buf_1 _45844_ (.A(\delay_line[8][3] ),
    .X(_08921_));
 sky130_fd_sc_hd__buf_1 _45845_ (.A(_08921_),
    .X(_08932_));
 sky130_fd_sc_hd__or2_1 _45846_ (.A(_03172_),
    .B(_08932_),
    .X(_08943_));
 sky130_fd_sc_hd__clkbuf_2 _45847_ (.A(\delay_line[7][3] ),
    .X(_08954_));
 sky130_fd_sc_hd__buf_2 _45848_ (.A(_08954_),
    .X(_08965_));
 sky130_fd_sc_hd__inv_2 _45849_ (.A(_08921_),
    .Y(_08976_));
 sky130_fd_sc_hd__or2_1 _45850_ (.A(_08976_),
    .B(_03216_),
    .X(_08987_));
 sky130_fd_sc_hd__o311a_2 _45851_ (.A1(_22985_),
    .A2(_03161_),
    .A3(_08943_),
    .B1(_08965_),
    .C1(_08987_),
    .X(_08998_));
 sky130_fd_sc_hd__clkbuf_2 _45852_ (.A(_03183_),
    .X(_09009_));
 sky130_fd_sc_hd__buf_2 _45853_ (.A(_08932_),
    .X(_09020_));
 sky130_fd_sc_hd__or4_1 _45854_ (.A(_22985_),
    .B(_03161_),
    .C(_09009_),
    .D(_09020_),
    .X(_09031_));
 sky130_fd_sc_hd__a21oi_2 _45855_ (.A1(_09031_),
    .A2(_08987_),
    .B1(_08965_),
    .Y(_09042_));
 sky130_fd_sc_hd__or3_1 _45856_ (.A(_08910_),
    .B(_08998_),
    .C(_09042_),
    .X(_09053_));
 sky130_fd_sc_hd__clkbuf_2 _45857_ (.A(_09053_),
    .X(_09064_));
 sky130_fd_sc_hd__o21ai_2 _45858_ (.A1(_08998_),
    .A2(_09042_),
    .B1(_08910_),
    .Y(_09075_));
 sky130_fd_sc_hd__and3_1 _45859_ (.A(_02931_),
    .B(_09064_),
    .C(_09075_),
    .X(_09086_));
 sky130_fd_sc_hd__a21oi_1 _45860_ (.A1(_09064_),
    .A2(_09075_),
    .B1(_02931_),
    .Y(_09097_));
 sky130_fd_sc_hd__nor2_1 _45861_ (.A(_09086_),
    .B(_09097_),
    .Y(_09108_));
 sky130_fd_sc_hd__xor2_1 _45862_ (.A(_03271_),
    .B(_09108_),
    .X(_09118_));
 sky130_fd_sc_hd__a21o_1 _45863_ (.A1(_08833_),
    .A2(_08866_),
    .B1(_09118_),
    .X(_09129_));
 sky130_fd_sc_hd__nand3_1 _45864_ (.A(_08833_),
    .B(_08866_),
    .C(_09118_),
    .Y(_09140_));
 sky130_fd_sc_hd__nand3_2 _45865_ (.A(_07920_),
    .B(_09129_),
    .C(_09140_),
    .Y(_09151_));
 sky130_fd_sc_hd__xnor2_1 _45866_ (.A(_03271_),
    .B(_09108_),
    .Y(_09162_));
 sky130_fd_sc_hd__a21o_1 _45867_ (.A1(_08833_),
    .A2(_08866_),
    .B1(_09162_),
    .X(_09173_));
 sky130_fd_sc_hd__inv_2 _45868_ (.A(_07920_),
    .Y(_09184_));
 sky130_fd_sc_hd__nand3_1 _45869_ (.A(_08833_),
    .B(_08866_),
    .C(_09162_),
    .Y(_09195_));
 sky130_fd_sc_hd__nand3_2 _45870_ (.A(_09173_),
    .B(_09184_),
    .C(_09195_),
    .Y(_09206_));
 sky130_fd_sc_hd__inv_2 _45871_ (.A(\delay_line[6][3] ),
    .Y(_09217_));
 sky130_fd_sc_hd__clkbuf_4 _45872_ (.A(_09217_),
    .X(_09228_));
 sky130_fd_sc_hd__nor2_1 _45873_ (.A(_09228_),
    .B(_03227_),
    .Y(_09239_));
 sky130_fd_sc_hd__o31a_1 _45874_ (.A1(_03238_),
    .A2(_03194_),
    .A3(net280),
    .B1(_09228_),
    .X(_09250_));
 sky130_fd_sc_hd__nor2_2 _45875_ (.A(_09239_),
    .B(_09250_),
    .Y(_09261_));
 sky130_fd_sc_hd__xor2_4 _45876_ (.A(_03436_),
    .B(_09261_),
    .X(_09272_));
 sky130_fd_sc_hd__nand2_1 _45877_ (.A(_22842_),
    .B(_03502_),
    .Y(_09283_));
 sky130_fd_sc_hd__or2b_1 _45878_ (.A(net437),
    .B_N(\delay_line[2][3] ),
    .X(_09294_));
 sky130_fd_sc_hd__clkbuf_2 _45879_ (.A(\delay_line[2][3] ),
    .X(_09305_));
 sky130_fd_sc_hd__inv_2 _45880_ (.A(_09305_),
    .Y(_09316_));
 sky130_fd_sc_hd__nand2_1 _45881_ (.A(_09316_),
    .B(net437),
    .Y(_09327_));
 sky130_fd_sc_hd__and4b_1 _45882_ (.A_N(\delay_line[3][0] ),
    .B(_09294_),
    .C(_09327_),
    .D(\delay_line[2][2] ),
    .X(_09338_));
 sky130_fd_sc_hd__o2bb2a_1 _45883_ (.A1_N(_09294_),
    .A2_N(_09327_),
    .B1(\delay_line[3][0] ),
    .B2(_03678_),
    .X(_09349_));
 sky130_fd_sc_hd__or2_1 _45884_ (.A(_09338_),
    .B(_09349_),
    .X(_09360_));
 sky130_fd_sc_hd__buf_1 _45885_ (.A(_09360_),
    .X(_09371_));
 sky130_fd_sc_hd__and3_1 _45886_ (.A(_09283_),
    .B(_03623_),
    .C(_09371_),
    .X(_09382_));
 sky130_fd_sc_hd__buf_1 _45887_ (.A(_03623_),
    .X(_09393_));
 sky130_fd_sc_hd__a21oi_1 _45888_ (.A1(_09283_),
    .A2(_09393_),
    .B1(_09371_),
    .Y(_09404_));
 sky130_fd_sc_hd__nor2_2 _45889_ (.A(_09382_),
    .B(_09404_),
    .Y(_09415_));
 sky130_fd_sc_hd__nor2_1 _45890_ (.A(_22908_),
    .B(_24809_),
    .Y(_09426_));
 sky130_fd_sc_hd__clkbuf_2 _45891_ (.A(\delay_line[6][1] ),
    .X(_09437_));
 sky130_fd_sc_hd__and2_1 _45892_ (.A(_22897_),
    .B(_09437_),
    .X(_09448_));
 sky130_fd_sc_hd__clkbuf_2 _45893_ (.A(\delay_line[5][3] ),
    .X(_09459_));
 sky130_fd_sc_hd__and3_1 _45894_ (.A(_24864_),
    .B(net431),
    .C(_09459_),
    .X(_09470_));
 sky130_fd_sc_hd__clkbuf_2 _45895_ (.A(_09459_),
    .X(_09481_));
 sky130_fd_sc_hd__a21oi_1 _45896_ (.A1(_24875_),
    .A2(_03535_),
    .B1(_09481_),
    .Y(_09492_));
 sky130_fd_sc_hd__xnor2_2 _45897_ (.A(_03579_),
    .B(net436),
    .Y(_09503_));
 sky130_fd_sc_hd__nor3_2 _45898_ (.A(_09470_),
    .B(_09492_),
    .C(_09503_),
    .Y(_09514_));
 sky130_fd_sc_hd__o21a_1 _45899_ (.A1(_09470_),
    .A2(_09492_),
    .B1(_09503_),
    .X(_09525_));
 sky130_fd_sc_hd__nor4_1 _45900_ (.A(_09426_),
    .B(_09448_),
    .C(_09514_),
    .D(_09525_),
    .Y(_09536_));
 sky130_fd_sc_hd__o22a_1 _45901_ (.A1(_09426_),
    .A2(_09448_),
    .B1(_09514_),
    .B2(_09525_),
    .X(_09547_));
 sky130_fd_sc_hd__nor2_2 _45902_ (.A(net240),
    .B(_09547_),
    .Y(_09558_));
 sky130_fd_sc_hd__xor2_4 _45903_ (.A(_03645_),
    .B(_09558_),
    .X(_09569_));
 sky130_fd_sc_hd__xnor2_4 _45904_ (.A(_09415_),
    .B(_09569_),
    .Y(_09580_));
 sky130_fd_sc_hd__xor2_4 _45905_ (.A(_09272_),
    .B(_09580_),
    .X(_09591_));
 sky130_fd_sc_hd__nand2_1 _45906_ (.A(_03480_),
    .B(_03777_),
    .Y(_09602_));
 sky130_fd_sc_hd__or2_1 _45907_ (.A(_03293_),
    .B(_09602_),
    .X(_09613_));
 sky130_fd_sc_hd__nand2_1 _45908_ (.A(_09602_),
    .B(_03293_),
    .Y(_09624_));
 sky130_fd_sc_hd__nand2_1 _45909_ (.A(_09613_),
    .B(_09624_),
    .Y(_09635_));
 sky130_fd_sc_hd__xor2_1 _45910_ (.A(_09591_),
    .B(_09635_),
    .X(_09646_));
 sky130_fd_sc_hd__a21o_1 _45911_ (.A1(_09151_),
    .A2(_09206_),
    .B1(_09646_),
    .X(_09657_));
 sky130_fd_sc_hd__o2bb2a_1 _45912_ (.A1_N(_03799_),
    .A2_N(_03359_),
    .B1(_03821_),
    .B2(_03337_),
    .X(_09668_));
 sky130_fd_sc_hd__nand3_1 _45913_ (.A(_09646_),
    .B(_09151_),
    .C(_09206_),
    .Y(_09679_));
 sky130_fd_sc_hd__nand3_1 _45914_ (.A(_09657_),
    .B(_09668_),
    .C(_09679_),
    .Y(_09690_));
 sky130_fd_sc_hd__xnor2_2 _45915_ (.A(_09591_),
    .B(_09635_),
    .Y(_09701_));
 sky130_fd_sc_hd__a31oi_2 _45916_ (.A1(_09151_),
    .A2(_09206_),
    .A3(_09701_),
    .B1(_09668_),
    .Y(_09712_));
 sky130_fd_sc_hd__a21o_1 _45917_ (.A1(_09151_),
    .A2(_09206_),
    .B1(_09701_),
    .X(_09723_));
 sky130_fd_sc_hd__nand2_1 _45918_ (.A(_09712_),
    .B(_09723_),
    .Y(_09734_));
 sky130_fd_sc_hd__buf_1 _45919_ (.A(\delay_line[1][2] ),
    .X(_09745_));
 sky130_fd_sc_hd__and2b_1 _45920_ (.A_N(_09745_),
    .B(\delay_line[1][3] ),
    .X(_09756_));
 sky130_fd_sc_hd__buf_1 _45921_ (.A(\delay_line[1][3] ),
    .X(_09767_));
 sky130_fd_sc_hd__nor2b_1 _45922_ (.A(_09767_),
    .B_N(_09745_),
    .Y(_09778_));
 sky130_fd_sc_hd__or3_1 _45923_ (.A(\delay_line[2][0] ),
    .B(_09756_),
    .C(_09778_),
    .X(_09789_));
 sky130_fd_sc_hd__clkbuf_2 _45924_ (.A(_09756_),
    .X(_09800_));
 sky130_fd_sc_hd__o21ai_1 _45925_ (.A1(_09800_),
    .A2(_09778_),
    .B1(\delay_line[2][0] ),
    .Y(_09811_));
 sky130_fd_sc_hd__and2_2 _45926_ (.A(_00249_),
    .B(_03898_),
    .X(_09822_));
 sky130_fd_sc_hd__and3_1 _45927_ (.A(_23414_),
    .B(\delay_line[1][1] ),
    .C(_03898_),
    .X(_09833_));
 sky130_fd_sc_hd__o21ba_1 _45928_ (.A1(_00260_),
    .A2(_09822_),
    .B1_N(_09833_),
    .X(_09844_));
 sky130_fd_sc_hd__a21oi_1 _45929_ (.A1(_09789_),
    .A2(_09811_),
    .B1(_09844_),
    .Y(_09855_));
 sky130_fd_sc_hd__o21ai_1 _45930_ (.A1(_03887_),
    .A2(_03898_),
    .B1(_23370_),
    .Y(_09866_));
 sky130_fd_sc_hd__and3_2 _45931_ (.A(_09844_),
    .B(_09789_),
    .C(_09811_),
    .X(_09877_));
 sky130_fd_sc_hd__nor3_1 _45932_ (.A(_09855_),
    .B(_09866_),
    .C(_09877_),
    .Y(_09888_));
 sky130_fd_sc_hd__inv_2 _45933_ (.A(_09888_),
    .Y(_09899_));
 sky130_fd_sc_hd__o21ai_1 _45934_ (.A1(_09877_),
    .A2(_09855_),
    .B1(_09866_),
    .Y(_09910_));
 sky130_fd_sc_hd__and3_1 _45935_ (.A(_09899_),
    .B(_09910_),
    .C(_03711_),
    .X(_09921_));
 sky130_fd_sc_hd__a21oi_1 _45936_ (.A1(_09899_),
    .A2(_09910_),
    .B1(_03711_),
    .Y(_09932_));
 sky130_fd_sc_hd__a211o_1 _45937_ (.A1(_03656_),
    .A2(_03755_),
    .B1(_09921_),
    .C1(_09932_),
    .X(_09943_));
 sky130_fd_sc_hd__o211ai_2 _45938_ (.A1(_09921_),
    .A2(_09932_),
    .B1(_03656_),
    .C1(_03755_),
    .Y(_09954_));
 sky130_fd_sc_hd__a21o_1 _45939_ (.A1(_09943_),
    .A2(_09954_),
    .B1(_03964_),
    .X(_09965_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45940_ (.A(_09943_),
    .X(_09976_));
 sky130_fd_sc_hd__nand3_2 _45941_ (.A(_09976_),
    .B(_09954_),
    .C(_03964_),
    .Y(_09987_));
 sky130_fd_sc_hd__or4bb_4 _45942_ (.A(_24985_),
    .B(_03788_),
    .C_N(_09965_),
    .D_N(_09987_),
    .X(_09998_));
 sky130_fd_sc_hd__a2bb2o_1 _45943_ (.A1_N(_24996_),
    .A2_N(_03788_),
    .B1(_09965_),
    .B2(_09987_),
    .X(_10009_));
 sky130_fd_sc_hd__nand2_1 _45944_ (.A(_09998_),
    .B(_10009_),
    .Y(_10020_));
 sky130_fd_sc_hd__and3_1 _45945_ (.A(_10020_),
    .B(_03997_),
    .C(_03986_),
    .X(_10031_));
 sky130_fd_sc_hd__and3_1 _45946_ (.A(_03975_),
    .B(_09998_),
    .C(_10009_),
    .X(_10042_));
 sky130_fd_sc_hd__o2bb2ai_1 _45947_ (.A1_N(_09690_),
    .A2_N(_09734_),
    .B1(_10031_),
    .B2(_10042_),
    .Y(_10053_));
 sky130_fd_sc_hd__and4_1 _45948_ (.A(_09998_),
    .B(_10009_),
    .C(_03986_),
    .D(_03997_),
    .X(_10064_));
 sky130_fd_sc_hd__a22oi_4 _45949_ (.A1(_03986_),
    .A2(_03997_),
    .B1(_09998_),
    .B2(_10009_),
    .Y(_10075_));
 sky130_fd_sc_hd__buf_2 _45950_ (.A(_09690_),
    .X(_10086_));
 sky130_fd_sc_hd__buf_2 _45951_ (.A(_09734_),
    .X(_10097_));
 sky130_fd_sc_hd__o211ai_2 _45952_ (.A1(_10064_),
    .A2(_10075_),
    .B1(_10086_),
    .C1(_10097_),
    .Y(_10108_));
 sky130_fd_sc_hd__o211a_1 _45953_ (.A1(_03854_),
    .A2(_03865_),
    .B1(_00183_),
    .C1(_00216_),
    .X(_10119_));
 sky130_fd_sc_hd__o31ai_2 _45954_ (.A1(_04019_),
    .A2(_04030_),
    .A3(_10119_),
    .B1(_03843_),
    .Y(_10130_));
 sky130_fd_sc_hd__inv_2 _45955_ (.A(_10130_),
    .Y(_10141_));
 sky130_fd_sc_hd__nand3_4 _45956_ (.A(_10053_),
    .B(_10108_),
    .C(_10141_),
    .Y(_10152_));
 sky130_fd_sc_hd__o2bb2ai_4 _45957_ (.A1_N(_10086_),
    .A2_N(_10097_),
    .B1(_10064_),
    .B2(_10075_),
    .Y(_10163_));
 sky130_fd_sc_hd__o211ai_4 _45958_ (.A1(_10031_),
    .A2(_10042_),
    .B1(_10086_),
    .C1(_10097_),
    .Y(_10174_));
 sky130_fd_sc_hd__nand3_4 _45959_ (.A(net99),
    .B(_10163_),
    .C(_10174_),
    .Y(_10185_));
 sky130_fd_sc_hd__nand3_2 _45960_ (.A(_24996_),
    .B(_25007_),
    .C(_22941_),
    .Y(_10196_));
 sky130_fd_sc_hd__nand2_2 _45961_ (.A(_03975_),
    .B(_04008_),
    .Y(_10207_));
 sky130_fd_sc_hd__o2bb2ai_2 _45962_ (.A1_N(_10152_),
    .A2_N(_10185_),
    .B1(_10196_),
    .B2(_10207_),
    .Y(_10218_));
 sky130_fd_sc_hd__nor2_1 _45963_ (.A(_10031_),
    .B(_10042_),
    .Y(_10229_));
 sky130_fd_sc_hd__a21oi_2 _45964_ (.A1(_10086_),
    .A2(_10097_),
    .B1(_10229_),
    .Y(_10240_));
 sky130_fd_sc_hd__a31o_1 _45965_ (.A1(_10086_),
    .A2(_10097_),
    .A3(_10229_),
    .B1(net99),
    .X(_10251_));
 sky130_fd_sc_hd__o211ai_4 _45966_ (.A1(_10240_),
    .A2(_10251_),
    .B1(_04052_),
    .C1(_10185_),
    .Y(_10262_));
 sky130_fd_sc_hd__nand2_2 _45967_ (.A(_04085_),
    .B(_04096_),
    .Y(_10273_));
 sky130_fd_sc_hd__a21oi_2 _45968_ (.A1(_10218_),
    .A2(_10262_),
    .B1(_10273_),
    .Y(_10284_));
 sky130_fd_sc_hd__inv_2 _45969_ (.A(_10273_),
    .Y(_10295_));
 sky130_fd_sc_hd__a2bb2oi_4 _45970_ (.A1_N(_10196_),
    .A2_N(_10207_),
    .B1(_10152_),
    .B2(_10185_),
    .Y(_10306_));
 sky130_fd_sc_hd__o211a_2 _45971_ (.A1(_10240_),
    .A2(_10251_),
    .B1(_04052_),
    .C1(_10185_),
    .X(_10317_));
 sky130_fd_sc_hd__nor3_4 _45972_ (.A(_10295_),
    .B(_10306_),
    .C(_10317_),
    .Y(_10328_));
 sky130_fd_sc_hd__buf_2 _45973_ (.A(\delay_line[23][3] ),
    .X(_10339_));
 sky130_fd_sc_hd__nor2_1 _45974_ (.A(_04579_),
    .B(_10339_),
    .Y(_10350_));
 sky130_fd_sc_hd__and2_2 _45975_ (.A(\delay_line[23][2] ),
    .B(\delay_line[23][3] ),
    .X(_10361_));
 sky130_fd_sc_hd__or2_2 _45976_ (.A(_10350_),
    .B(_10361_),
    .X(_10372_));
 sky130_fd_sc_hd__o21ai_1 _45977_ (.A1(_10284_),
    .A2(_10328_),
    .B1(_10372_),
    .Y(_10383_));
 sky130_fd_sc_hd__nand3_4 _45978_ (.A(_10273_),
    .B(_10218_),
    .C(_10262_),
    .Y(_10394_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _45979_ (.A(_10394_),
    .X(_10405_));
 sky130_fd_sc_hd__o21ai_4 _45980_ (.A1(_10306_),
    .A2(_10317_),
    .B1(_10295_),
    .Y(_10416_));
 sky130_fd_sc_hd__nand3b_1 _45981_ (.A_N(_10372_),
    .B(_10405_),
    .C(_10416_),
    .Y(_10426_));
 sky130_fd_sc_hd__o211a_1 _45982_ (.A1(_04228_),
    .A2(_04261_),
    .B1(_10383_),
    .C1(_10426_),
    .X(_10437_));
 sky130_fd_sc_hd__a21o_1 _45983_ (.A1(_10416_),
    .A2(_10405_),
    .B1(_10372_),
    .X(_10448_));
 sky130_fd_sc_hd__a31o_1 _45984_ (.A1(_04107_),
    .A2(_04239_),
    .A3(_04085_),
    .B1(_04228_),
    .X(_10459_));
 sky130_fd_sc_hd__inv_2 _45985_ (.A(_10459_),
    .Y(_10470_));
 sky130_fd_sc_hd__o211ai_1 _45986_ (.A1(_10350_),
    .A2(_10361_),
    .B1(_10416_),
    .C1(_10405_),
    .Y(_10481_));
 sky130_fd_sc_hd__and3_1 _45987_ (.A(_10448_),
    .B(_10470_),
    .C(_10481_),
    .X(_10492_));
 sky130_fd_sc_hd__a21bo_1 _45988_ (.A1(_04590_),
    .A2(\delay_line[23][0] ),
    .B1_N(_04601_),
    .X(_10503_));
 sky130_fd_sc_hd__o21bai_2 _45989_ (.A1(_10437_),
    .A2(_10492_),
    .B1_N(_10503_),
    .Y(_10514_));
 sky130_fd_sc_hd__nand2_1 _45990_ (.A(_10383_),
    .B(_10426_),
    .Y(_10525_));
 sky130_fd_sc_hd__a21boi_2 _45991_ (.A1(_10525_),
    .A2(_10470_),
    .B1_N(_10503_),
    .Y(_10536_));
 sky130_fd_sc_hd__o21ai_2 _45992_ (.A1(_10470_),
    .A2(_10525_),
    .B1(_10536_),
    .Y(_10547_));
 sky130_fd_sc_hd__a31o_1 _45993_ (.A1(_04283_),
    .A2(_04382_),
    .A3(_04393_),
    .B1(_04437_),
    .X(_10558_));
 sky130_fd_sc_hd__a21oi_4 _45994_ (.A1(_10514_),
    .A2(_10547_),
    .B1(_10558_),
    .Y(_10569_));
 sky130_fd_sc_hd__o211a_4 _45995_ (.A1(_04404_),
    .A2(net91),
    .B1(_10514_),
    .C1(_10547_),
    .X(_10580_));
 sky130_fd_sc_hd__or2_1 _45996_ (.A(_10569_),
    .B(_10580_),
    .X(_10591_));
 sky130_fd_sc_hd__a41o_1 _45997_ (.A1(_00359_),
    .A2(_04678_),
    .A3(_00381_),
    .A4(_00480_),
    .B1(_04656_),
    .X(_10602_));
 sky130_fd_sc_hd__xnor2_1 _45998_ (.A(_10591_),
    .B(_10602_),
    .Y(_10613_));
 sky130_fd_sc_hd__or2_1 _45999_ (.A(_07909_),
    .B(_10613_),
    .X(_10624_));
 sky130_fd_sc_hd__buf_2 _46000_ (.A(_07909_),
    .X(_10635_));
 sky130_fd_sc_hd__nand2_1 _46001_ (.A(_10635_),
    .B(_10613_),
    .Y(_10646_));
 sky130_fd_sc_hd__a41o_1 _46002_ (.A1(_04503_),
    .A2(_00667_),
    .A3(_00678_),
    .A4(_00513_),
    .B1(_04492_),
    .X(_10657_));
 sky130_fd_sc_hd__a21oi_1 _46003_ (.A1(_10624_),
    .A2(_10646_),
    .B1(_10657_),
    .Y(_10668_));
 sky130_fd_sc_hd__nand3_2 _46004_ (.A(_10657_),
    .B(_10624_),
    .C(_10646_),
    .Y(_10679_));
 sky130_fd_sc_hd__inv_2 _46005_ (.A(_10679_),
    .Y(_10690_));
 sky130_fd_sc_hd__nor3_2 _46006_ (.A(_07898_),
    .B(_10668_),
    .C(_10690_),
    .Y(_10701_));
 sky130_fd_sc_hd__o21a_1 _46007_ (.A1(_10668_),
    .A2(_10690_),
    .B1(_07898_),
    .X(_10712_));
 sky130_fd_sc_hd__o21bai_1 _46008_ (.A1(_04733_),
    .A2(_04546_),
    .B1_N(_04755_),
    .Y(_10723_));
 sky130_fd_sc_hd__o21bai_2 _46009_ (.A1(_10701_),
    .A2(_10712_),
    .B1_N(_10723_),
    .Y(_10734_));
 sky130_fd_sc_hd__or3b_1 _46010_ (.A(_10701_),
    .B(_10712_),
    .C_N(_10723_),
    .X(_10745_));
 sky130_fd_sc_hd__nand2_1 _46011_ (.A(_04832_),
    .B(_04854_),
    .Y(_10756_));
 sky130_fd_sc_hd__buf_2 _46012_ (.A(_10756_),
    .X(_10767_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46013_ (.A(\delay_line[17][2] ),
    .X(_10778_));
 sky130_fd_sc_hd__a21o_1 _46014_ (.A1(net378),
    .A2(_10778_),
    .B1(_04876_),
    .X(_10789_));
 sky130_fd_sc_hd__o21ai_1 _46015_ (.A1(\delay_line[17][0] ),
    .A2(_04887_),
    .B1(_04876_),
    .Y(_10800_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46016_ (.A(\delay_line[17][3] ),
    .X(_10811_));
 sky130_fd_sc_hd__nor2_1 _46017_ (.A(_04887_),
    .B(_10811_),
    .Y(_10822_));
 sky130_fd_sc_hd__nand2_2 _46018_ (.A(\delay_line[17][2] ),
    .B(\delay_line[17][3] ),
    .Y(_10833_));
 sky130_fd_sc_hd__and2b_2 _46019_ (.A_N(_10822_),
    .B(_10833_),
    .X(_10844_));
 sky130_fd_sc_hd__a21o_1 _46020_ (.A1(_10789_),
    .A2(_10800_),
    .B1(_10844_),
    .X(_10855_));
 sky130_fd_sc_hd__nand2_2 _46021_ (.A(\delay_line[17][1] ),
    .B(_04887_),
    .Y(_10866_));
 sky130_fd_sc_hd__o2111ai_4 _46022_ (.A1(_04920_),
    .A2(_22139_),
    .B1(_10866_),
    .C1(_10789_),
    .D1(_10844_),
    .Y(_10877_));
 sky130_fd_sc_hd__clkbuf_2 _46023_ (.A(\delay_line[20][3] ),
    .X(_10888_));
 sky130_fd_sc_hd__and2_1 _46024_ (.A(net367),
    .B(_10888_),
    .X(_10899_));
 sky130_fd_sc_hd__clkbuf_2 _46025_ (.A(_10899_),
    .X(_10910_));
 sky130_fd_sc_hd__nor2_1 _46026_ (.A(net367),
    .B(_10888_),
    .Y(_10921_));
 sky130_fd_sc_hd__buf_2 _46027_ (.A(\delay_line[20][2] ),
    .X(_10932_));
 sky130_fd_sc_hd__a21boi_1 _46028_ (.A1(_23600_),
    .A2(_10932_),
    .B1_N(_04832_),
    .Y(_10943_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46029_ (.A(_10943_),
    .X(_10954_));
 sky130_fd_sc_hd__or3_2 _46030_ (.A(_10910_),
    .B(_10921_),
    .C(_10954_),
    .X(_10965_));
 sky130_fd_sc_hd__o21ai_1 _46031_ (.A1(_10910_),
    .A2(_10921_),
    .B1(_10954_),
    .Y(_10976_));
 sky130_fd_sc_hd__nor2_1 _46032_ (.A(\delay_line[20][0] ),
    .B(net368),
    .Y(_10987_));
 sky130_fd_sc_hd__nand2_1 _46033_ (.A(_22161_),
    .B(\delay_line[20][1] ),
    .Y(_10998_));
 sky130_fd_sc_hd__and2b_1 _46034_ (.A_N(_10987_),
    .B(_10998_),
    .X(_11009_));
 sky130_fd_sc_hd__clkbuf_2 _46035_ (.A(_11009_),
    .X(_11020_));
 sky130_fd_sc_hd__a21o_1 _46036_ (.A1(_10965_),
    .A2(_10976_),
    .B1(_11020_),
    .X(_11031_));
 sky130_fd_sc_hd__buf_2 _46037_ (.A(_10888_),
    .X(_11042_));
 sky130_fd_sc_hd__nand2_4 _46038_ (.A(_11042_),
    .B(_11020_),
    .Y(_11053_));
 sky130_fd_sc_hd__nand4_2 _46039_ (.A(_10855_),
    .B(_10877_),
    .C(_11031_),
    .D(_11053_),
    .Y(_11064_));
 sky130_fd_sc_hd__a22oi_2 _46040_ (.A1(_10855_),
    .A2(_10877_),
    .B1(_11031_),
    .B2(_11053_),
    .Y(_11075_));
 sky130_fd_sc_hd__inv_2 _46041_ (.A(_11075_),
    .Y(_11086_));
 sky130_fd_sc_hd__nand2_1 _46042_ (.A(_11064_),
    .B(_11086_),
    .Y(_11097_));
 sky130_fd_sc_hd__xnor2_1 _46043_ (.A(_04711_),
    .B(_11097_),
    .Y(_11108_));
 sky130_fd_sc_hd__or4bb_2 _46044_ (.A(_10767_),
    .B(_11108_),
    .C_N(_04964_),
    .D_N(_04942_),
    .X(_11119_));
 sky130_fd_sc_hd__or2b_1 _46045_ (.A(_04975_),
    .B_N(_11108_),
    .X(_11130_));
 sky130_fd_sc_hd__nand2_1 _46046_ (.A(_11119_),
    .B(_11130_),
    .Y(_11141_));
 sky130_fd_sc_hd__nand3_1 _46047_ (.A(_10734_),
    .B(_10745_),
    .C(_11141_),
    .Y(_11152_));
 sky130_fd_sc_hd__a21o_1 _46048_ (.A1(_10734_),
    .A2(_10745_),
    .B1(_11141_),
    .X(_11163_));
 sky130_fd_sc_hd__o2111ai_1 _46049_ (.A1(_05063_),
    .A2(_05030_),
    .B1(_11152_),
    .C1(_11163_),
    .D1(_04788_),
    .Y(_11174_));
 sky130_fd_sc_hd__a22o_1 _46050_ (.A1(_04788_),
    .A2(_05074_),
    .B1(_11152_),
    .B2(_11163_),
    .X(_11185_));
 sky130_fd_sc_hd__nand2_1 _46051_ (.A(_11174_),
    .B(_11185_),
    .Y(_11196_));
 sky130_fd_sc_hd__xor2_1 _46052_ (.A(_05183_),
    .B(_11196_),
    .X(_11207_));
 sky130_fd_sc_hd__o32a_1 _46053_ (.A1(_05107_),
    .A2(_05041_),
    .A3(_05085_),
    .B1(_00919_),
    .B2(_05118_),
    .X(_11218_));
 sky130_fd_sc_hd__nand2_1 _46054_ (.A(_05183_),
    .B(_11174_),
    .Y(_11229_));
 sky130_fd_sc_hd__or3b_1 _46055_ (.A(_11075_),
    .B(_04711_),
    .C_N(_11064_),
    .X(_11240_));
 sky130_fd_sc_hd__a21o_1 _46056_ (.A1(_11240_),
    .A2(_11119_),
    .B1(_10877_),
    .X(_11251_));
 sky130_fd_sc_hd__o211ai_1 _46057_ (.A1(_04711_),
    .A2(_11097_),
    .B1(_11119_),
    .C1(_10877_),
    .Y(_11262_));
 sky130_fd_sc_hd__nand2_1 _46058_ (.A(_11251_),
    .B(_11262_),
    .Y(_11273_));
 sky130_fd_sc_hd__nand2_1 _46059_ (.A(_10745_),
    .B(_11141_),
    .Y(_11284_));
 sky130_fd_sc_hd__clkbuf_2 _46060_ (.A(\delay_line[17][4] ),
    .X(_11295_));
 sky130_fd_sc_hd__xor2_1 _46061_ (.A(_11295_),
    .B(\delay_line[17][3] ),
    .X(_11306_));
 sky130_fd_sc_hd__nand3_1 _46062_ (.A(_11306_),
    .B(_23611_),
    .C(_22172_),
    .Y(_11317_));
 sky130_fd_sc_hd__buf_1 _46063_ (.A(_11306_),
    .X(_11328_));
 sky130_fd_sc_hd__a21o_1 _46064_ (.A1(_22183_),
    .A2(_23622_),
    .B1(_11328_),
    .X(_11339_));
 sky130_fd_sc_hd__or2b_1 _46065_ (.A(_10811_),
    .B_N(_04887_),
    .X(_11350_));
 sky130_fd_sc_hd__buf_1 _46066_ (.A(_10811_),
    .X(_11361_));
 sky130_fd_sc_hd__o2bb2a_1 _46067_ (.A1_N(_10800_),
    .A2_N(_11350_),
    .B1(_11361_),
    .B2(_10866_),
    .X(_11372_));
 sky130_fd_sc_hd__a21oi_1 _46068_ (.A1(_11317_),
    .A2(_11339_),
    .B1(_11372_),
    .Y(_11383_));
 sky130_fd_sc_hd__and3_1 _46069_ (.A(_11339_),
    .B(_11372_),
    .C(_11317_),
    .X(_11394_));
 sky130_fd_sc_hd__and2_2 _46070_ (.A(\delay_line[20][3] ),
    .B(\delay_line[20][4] ),
    .X(_11405_));
 sky130_fd_sc_hd__clkbuf_2 _46071_ (.A(\delay_line[20][4] ),
    .X(_11416_));
 sky130_fd_sc_hd__nor2_1 _46072_ (.A(_10888_),
    .B(_11416_),
    .Y(_11427_));
 sky130_fd_sc_hd__nor2_4 _46073_ (.A(_11405_),
    .B(_11427_),
    .Y(_11438_));
 sky130_fd_sc_hd__buf_1 _46074_ (.A(_11416_),
    .X(_11449_));
 sky130_fd_sc_hd__nand3b_4 _46075_ (.A_N(_11449_),
    .B(_11042_),
    .C(_10932_),
    .Y(_11460_));
 sky130_fd_sc_hd__o21a_1 _46076_ (.A1(_10910_),
    .A2(_11438_),
    .B1(_11460_),
    .X(_11471_));
 sky130_fd_sc_hd__and3_1 _46077_ (.A(_11471_),
    .B(_04865_),
    .C(_04843_),
    .X(_11482_));
 sky130_fd_sc_hd__a21oi_2 _46078_ (.A1(_04843_),
    .A2(_04865_),
    .B1(_11471_),
    .Y(_11493_));
 sky130_fd_sc_hd__a211oi_4 _46079_ (.A1(_10965_),
    .A2(_11053_),
    .B1(_11482_),
    .C1(_11493_),
    .Y(_11504_));
 sky130_fd_sc_hd__o211ai_1 _46080_ (.A1(_11482_),
    .A2(_11493_),
    .B1(_10965_),
    .C1(_11053_),
    .Y(_11515_));
 sky130_fd_sc_hd__inv_2 _46081_ (.A(_11515_),
    .Y(_11526_));
 sky130_fd_sc_hd__or4_4 _46082_ (.A(_11383_),
    .B(_11394_),
    .C(_11504_),
    .D(_11526_),
    .X(_11537_));
 sky130_fd_sc_hd__inv_2 _46083_ (.A(_11504_),
    .Y(_11548_));
 sky130_fd_sc_hd__a2bb2o_1 _46084_ (.A1_N(_11383_),
    .A2_N(_11394_),
    .B1(_11548_),
    .B2(_11515_),
    .X(_11559_));
 sky130_fd_sc_hd__nand2_1 _46085_ (.A(_11537_),
    .B(_11559_),
    .Y(_11570_));
 sky130_fd_sc_hd__xnor2_1 _46086_ (.A(_10679_),
    .B(_11570_),
    .Y(_11581_));
 sky130_fd_sc_hd__and2_1 _46087_ (.A(_11064_),
    .B(_11581_),
    .X(_11592_));
 sky130_fd_sc_hd__nor2_1 _46088_ (.A(_11064_),
    .B(_11581_),
    .Y(_11603_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46089_ (.A(_11603_),
    .X(_11614_));
 sky130_fd_sc_hd__and2_1 _46090_ (.A(_10635_),
    .B(_10613_),
    .X(_11625_));
 sky130_fd_sc_hd__inv_2 _46091_ (.A(_10569_),
    .Y(_11636_));
 sky130_fd_sc_hd__and4b_1 _46092_ (.A_N(_10580_),
    .B(_00502_),
    .C(_11636_),
    .D(_04678_),
    .X(_11647_));
 sky130_fd_sc_hd__inv_2 _46093_ (.A(_05667_),
    .Y(_11658_));
 sky130_fd_sc_hd__clkbuf_2 _46094_ (.A(_08668_),
    .X(_11669_));
 sky130_fd_sc_hd__inv_2 _46095_ (.A(net415),
    .Y(_11680_));
 sky130_fd_sc_hd__buf_2 _46096_ (.A(_11680_),
    .X(_11691_));
 sky130_fd_sc_hd__a221o_1 _46097_ (.A1(_23095_),
    .A2(_08877_),
    .B1(_11669_),
    .B2(_11691_),
    .C1(_08899_),
    .X(_11701_));
 sky130_fd_sc_hd__a21oi_1 _46098_ (.A1(_23084_),
    .A2(_08877_),
    .B1(_08899_),
    .Y(_11712_));
 sky130_fd_sc_hd__or3b_1 _46099_ (.A(_23117_),
    .B(_11712_),
    .C_N(_11669_),
    .X(_11723_));
 sky130_fd_sc_hd__nand2_1 _46100_ (.A(_03205_),
    .B(_08932_),
    .Y(_11734_));
 sky130_fd_sc_hd__nand3b_2 _46101_ (.A_N(_03150_),
    .B(_08943_),
    .C(_11734_),
    .Y(_11745_));
 sky130_fd_sc_hd__nor2_1 _46102_ (.A(_03205_),
    .B(_08932_),
    .Y(_11756_));
 sky130_fd_sc_hd__and2_1 _46103_ (.A(_03172_),
    .B(_08921_),
    .X(_11767_));
 sky130_fd_sc_hd__o21ai_2 _46104_ (.A1(_11756_),
    .A2(_11767_),
    .B1(_03150_),
    .Y(_11778_));
 sky130_fd_sc_hd__o21bai_2 _46105_ (.A1(_03205_),
    .A2(_00095_),
    .B1_N(_00084_),
    .Y(_11789_));
 sky130_fd_sc_hd__a21oi_4 _46106_ (.A1(_11745_),
    .A2(_11778_),
    .B1(_11789_),
    .Y(_11800_));
 sky130_fd_sc_hd__inv_2 _46107_ (.A(\delay_line[8][4] ),
    .Y(_11811_));
 sky130_fd_sc_hd__clkbuf_2 _46108_ (.A(_11811_),
    .X(_11822_));
 sky130_fd_sc_hd__buf_2 _46109_ (.A(_11822_),
    .X(_11833_));
 sky130_fd_sc_hd__and3_1 _46110_ (.A(_11745_),
    .B(_11778_),
    .C(_11789_),
    .X(_11844_));
 sky130_fd_sc_hd__nor3_2 _46111_ (.A(_11800_),
    .B(_11833_),
    .C(_11844_),
    .Y(_11855_));
 sky130_fd_sc_hd__buf_2 _46112_ (.A(_11833_),
    .X(_11866_));
 sky130_fd_sc_hd__o21a_1 _46113_ (.A1(_11844_),
    .A2(_11800_),
    .B1(_11866_),
    .X(_11877_));
 sky130_fd_sc_hd__nor2_1 _46114_ (.A(_11855_),
    .B(_11877_),
    .Y(_11888_));
 sky130_fd_sc_hd__buf_2 _46115_ (.A(_09009_),
    .X(_11899_));
 sky130_fd_sc_hd__a21oi_1 _46116_ (.A1(_11899_),
    .A2(_00117_),
    .B1(_08987_),
    .Y(_11910_));
 sky130_fd_sc_hd__nand2_1 _46117_ (.A(_11888_),
    .B(_11910_),
    .Y(_11921_));
 sky130_fd_sc_hd__o21bai_1 _46118_ (.A1(_11855_),
    .A2(_11877_),
    .B1_N(_11910_),
    .Y(_11932_));
 sky130_fd_sc_hd__clkbuf_2 _46119_ (.A(_03161_),
    .X(_11943_));
 sky130_fd_sc_hd__clkbuf_2 _46120_ (.A(\delay_line[7][4] ),
    .X(_11954_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46121_ (.A(_11954_),
    .X(_11965_));
 sky130_fd_sc_hd__buf_2 _46122_ (.A(_11965_),
    .X(_11976_));
 sky130_fd_sc_hd__a31o_1 _46123_ (.A1(_23051_),
    .A2(_11943_),
    .A3(_11899_),
    .B1(_11976_),
    .X(_11987_));
 sky130_fd_sc_hd__nand4_2 _46124_ (.A(_23040_),
    .B(_11943_),
    .C(_09009_),
    .D(_11976_),
    .Y(_11998_));
 sky130_fd_sc_hd__nand2_1 _46125_ (.A(_11987_),
    .B(_11998_),
    .Y(_12009_));
 sky130_fd_sc_hd__a21bo_1 _46126_ (.A1(_11921_),
    .A2(_11932_),
    .B1_N(_12009_),
    .X(_12020_));
 sky130_fd_sc_hd__nand4_2 _46127_ (.A(_11921_),
    .B(_11932_),
    .C(_11987_),
    .D(_11998_),
    .Y(_12031_));
 sky130_fd_sc_hd__a22o_1 _46128_ (.A1(_11701_),
    .A2(_11723_),
    .B1(_12020_),
    .B2(_12031_),
    .X(_12042_));
 sky130_fd_sc_hd__nand4_1 _46129_ (.A(_11701_),
    .B(_11723_),
    .C(_12020_),
    .D(_12031_),
    .Y(_12053_));
 sky130_fd_sc_hd__clkbuf_2 _46130_ (.A(_12053_),
    .X(_12064_));
 sky130_fd_sc_hd__a21oi_1 _46131_ (.A1(_12042_),
    .A2(_12064_),
    .B1(_08767_),
    .Y(_12075_));
 sky130_fd_sc_hd__and3_1 _46132_ (.A(_12042_),
    .B(_12053_),
    .C(_08767_),
    .X(_12086_));
 sky130_fd_sc_hd__or2_1 _46133_ (.A(_12075_),
    .B(_12086_),
    .X(_12097_));
 sky130_fd_sc_hd__xor2_1 _46134_ (.A(_09064_),
    .B(_12097_),
    .X(_12108_));
 sky130_fd_sc_hd__a21o_1 _46135_ (.A1(_08426_),
    .A2(_08514_),
    .B1(_08569_),
    .X(_12119_));
 sky130_fd_sc_hd__clkbuf_4 _46136_ (.A(\delay_line[12][4] ),
    .X(_12130_));
 sky130_fd_sc_hd__inv_2 _46137_ (.A(_12130_),
    .Y(_12141_));
 sky130_fd_sc_hd__buf_2 _46138_ (.A(net407),
    .X(_12152_));
 sky130_fd_sc_hd__and3_2 _46139_ (.A(_12141_),
    .B(_12152_),
    .C(_02414_),
    .X(_12163_));
 sky130_fd_sc_hd__clkbuf_2 _46140_ (.A(_12141_),
    .X(_12174_));
 sky130_fd_sc_hd__or3b_1 _46141_ (.A(_02425_),
    .B(_12174_),
    .C_N(_08481_),
    .X(_12185_));
 sky130_fd_sc_hd__o21ai_2 _46142_ (.A1(_12130_),
    .A2(_08481_),
    .B1(_12185_),
    .Y(_12196_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46143_ (.A(\delay_line[13][4] ),
    .X(_12207_));
 sky130_fd_sc_hd__nor2_1 _46144_ (.A(_23150_),
    .B(_12207_),
    .Y(_12218_));
 sky130_fd_sc_hd__and2_1 _46145_ (.A(_23150_),
    .B(\delay_line[13][4] ),
    .X(_12229_));
 sky130_fd_sc_hd__clkbuf_2 _46146_ (.A(\delay_line[4][1] ),
    .X(_12240_));
 sky130_fd_sc_hd__clkbuf_2 _46147_ (.A(_12240_),
    .X(_12251_));
 sky130_fd_sc_hd__buf_6 _46148_ (.A(\delay_line[11][2] ),
    .X(_12262_));
 sky130_fd_sc_hd__buf_6 _46149_ (.A(_12262_),
    .X(_12273_));
 sky130_fd_sc_hd__nor2_1 _46150_ (.A(_12251_),
    .B(_12273_),
    .Y(_12284_));
 sky130_fd_sc_hd__nand2_1 _46151_ (.A(_12240_),
    .B(_12273_),
    .Y(_12295_));
 sky130_fd_sc_hd__nand2_1 _46152_ (.A(_12295_),
    .B(\delay_line[0][4] ),
    .Y(_12306_));
 sky130_fd_sc_hd__o21a_1 _46153_ (.A1(_07975_),
    .A2(_08019_),
    .B1(\delay_line[0][3] ),
    .X(_12317_));
 sky130_fd_sc_hd__o22ai_4 _46154_ (.A1(_12284_),
    .A2(_12306_),
    .B1(_08008_),
    .B2(_12317_),
    .Y(_12328_));
 sky130_fd_sc_hd__inv_2 _46155_ (.A(_12240_),
    .Y(_12339_));
 sky130_fd_sc_hd__inv_2 _46156_ (.A(\delay_line[11][2] ),
    .Y(_12350_));
 sky130_fd_sc_hd__buf_2 _46157_ (.A(_12350_),
    .X(_12361_));
 sky130_fd_sc_hd__nand2_1 _46158_ (.A(_12339_),
    .B(_12361_),
    .Y(_12372_));
 sky130_fd_sc_hd__clkbuf_2 _46159_ (.A(\delay_line[0][4] ),
    .X(_12383_));
 sky130_fd_sc_hd__a21oi_2 _46160_ (.A1(_12295_),
    .A2(_12372_),
    .B1(_12383_),
    .Y(_12394_));
 sky130_fd_sc_hd__o21ai_1 _46161_ (.A1(_12284_),
    .A2(_12306_),
    .B1(_12383_),
    .Y(_12405_));
 sky130_fd_sc_hd__o21ai_2 _46162_ (.A1(_12251_),
    .A2(_12273_),
    .B1(\delay_line[0][4] ),
    .Y(_12416_));
 sky130_fd_sc_hd__nand3_1 _46163_ (.A(_12295_),
    .B(_12372_),
    .C(_12416_),
    .Y(_12427_));
 sky130_fd_sc_hd__o21a_1 _46164_ (.A1(_08129_),
    .A2(_08151_),
    .B1(_08030_),
    .X(_12438_));
 sky130_fd_sc_hd__nand3_2 _46165_ (.A(_12405_),
    .B(_12427_),
    .C(_12438_),
    .Y(_12449_));
 sky130_fd_sc_hd__o21ai_1 _46166_ (.A1(_12328_),
    .A2(_12394_),
    .B1(_12449_),
    .Y(_12460_));
 sky130_fd_sc_hd__nand2_1 _46167_ (.A(_08085_),
    .B(_12460_),
    .Y(_12471_));
 sky130_fd_sc_hd__o211ai_2 _46168_ (.A1(_12328_),
    .A2(_12394_),
    .B1(_08074_),
    .C1(_12449_),
    .Y(_12482_));
 sky130_fd_sc_hd__o21ai_1 _46169_ (.A1(_08140_),
    .A2(_08151_),
    .B1(_12317_),
    .Y(_12493_));
 sky130_fd_sc_hd__a31o_1 _46170_ (.A1(_08096_),
    .A2(_02513_),
    .A3(_12493_),
    .B1(_02524_),
    .X(_12504_));
 sky130_fd_sc_hd__a21oi_1 _46171_ (.A1(_12471_),
    .A2(_12482_),
    .B1(_12504_),
    .Y(_12515_));
 sky130_fd_sc_hd__a31oi_2 _46172_ (.A1(_08096_),
    .A2(_02513_),
    .A3(_12493_),
    .B1(_08118_),
    .Y(_12526_));
 sky130_fd_sc_hd__and2_1 _46173_ (.A(_12251_),
    .B(_12273_),
    .X(_12537_));
 sky130_fd_sc_hd__o21bai_1 _46174_ (.A1(_12537_),
    .A2(_12284_),
    .B1_N(\delay_line[0][4] ),
    .Y(_12548_));
 sky130_fd_sc_hd__o211ai_2 _46175_ (.A1(_12416_),
    .A2(_12537_),
    .B1(_08162_),
    .C1(_12548_),
    .Y(_12559_));
 sky130_fd_sc_hd__clkbuf_2 _46176_ (.A(_08074_),
    .X(_12570_));
 sky130_fd_sc_hd__a21oi_1 _46177_ (.A1(_12559_),
    .A2(_12449_),
    .B1(_12570_),
    .Y(_12581_));
 sky130_fd_sc_hd__o211a_1 _46178_ (.A1(_12328_),
    .A2(_12394_),
    .B1(_08074_),
    .C1(_12449_),
    .X(_12592_));
 sky130_fd_sc_hd__nor3_2 _46179_ (.A(_12526_),
    .B(_12581_),
    .C(_12592_),
    .Y(_12603_));
 sky130_fd_sc_hd__o22ai_1 _46180_ (.A1(_12218_),
    .A2(_12229_),
    .B1(_12515_),
    .B2(_12603_),
    .Y(_12614_));
 sky130_fd_sc_hd__o21ai_2 _46181_ (.A1(_12581_),
    .A2(_12592_),
    .B1(_12526_),
    .Y(_12625_));
 sky130_fd_sc_hd__nand3_2 _46182_ (.A(_12504_),
    .B(_12471_),
    .C(_12482_),
    .Y(_12636_));
 sky130_fd_sc_hd__nor2_1 _46183_ (.A(_12218_),
    .B(_12229_),
    .Y(_12647_));
 sky130_fd_sc_hd__nand3_1 _46184_ (.A(_12625_),
    .B(_12636_),
    .C(_12647_),
    .Y(_12658_));
 sky130_fd_sc_hd__a21bo_1 _46185_ (.A1(_08272_),
    .A2(_08261_),
    .B1_N(_08195_),
    .X(_12669_));
 sky130_fd_sc_hd__a21oi_1 _46186_ (.A1(_12614_),
    .A2(_12658_),
    .B1(_12669_),
    .Y(_12680_));
 sky130_fd_sc_hd__a21boi_2 _46187_ (.A1(_08272_),
    .A2(_08261_),
    .B1_N(_08195_),
    .Y(_12691_));
 sky130_fd_sc_hd__a21oi_2 _46188_ (.A1(_12625_),
    .A2(_12636_),
    .B1(_12647_),
    .Y(_12702_));
 sky130_fd_sc_hd__and3_1 _46189_ (.A(_12625_),
    .B(_12636_),
    .C(_12647_),
    .X(_12713_));
 sky130_fd_sc_hd__buf_2 _46190_ (.A(_12713_),
    .X(_12724_));
 sky130_fd_sc_hd__nor3_4 _46191_ (.A(_12691_),
    .B(_12702_),
    .C(_12724_),
    .Y(_12735_));
 sky130_fd_sc_hd__buf_2 _46192_ (.A(_02480_),
    .X(_12746_));
 sky130_fd_sc_hd__o21bai_4 _46193_ (.A1(_12680_),
    .A2(_12735_),
    .B1_N(_12746_),
    .Y(_12757_));
 sky130_fd_sc_hd__nand2_1 _46194_ (.A(_12669_),
    .B(_12614_),
    .Y(_12768_));
 sky130_fd_sc_hd__o21ai_1 _46195_ (.A1(_12702_),
    .A2(_12713_),
    .B1(_12691_),
    .Y(_12779_));
 sky130_fd_sc_hd__o211ai_2 _46196_ (.A1(_12724_),
    .A2(_12768_),
    .B1(_12746_),
    .C1(_12779_),
    .Y(_12790_));
 sky130_fd_sc_hd__nor2_1 _46197_ (.A(_25215_),
    .B(_08382_),
    .Y(_12801_));
 sky130_fd_sc_hd__a31o_1 _46198_ (.A1(_08305_),
    .A2(_08294_),
    .A3(_08338_),
    .B1(_12801_),
    .X(_12812_));
 sky130_fd_sc_hd__a21oi_2 _46199_ (.A1(_12757_),
    .A2(_12790_),
    .B1(_12812_),
    .Y(_12823_));
 sky130_fd_sc_hd__nand2_2 _46200_ (.A(_12779_),
    .B(_12746_),
    .Y(_12834_));
 sky130_fd_sc_hd__o221a_1 _46201_ (.A1(_08371_),
    .A2(_12801_),
    .B1(_12735_),
    .B2(_12834_),
    .C1(_12757_),
    .X(_12845_));
 sky130_fd_sc_hd__o22ai_2 _46202_ (.A1(_12163_),
    .A2(_12196_),
    .B1(_12823_),
    .B2(_12845_),
    .Y(_12856_));
 sky130_fd_sc_hd__or2_1 _46203_ (.A(_12163_),
    .B(_12196_),
    .X(_12867_));
 sky130_fd_sc_hd__a21o_1 _46204_ (.A1(_12757_),
    .A2(_12790_),
    .B1(_12812_),
    .X(_12877_));
 sky130_fd_sc_hd__o221ai_4 _46205_ (.A1(_08371_),
    .A2(_12801_),
    .B1(_12735_),
    .B2(_12834_),
    .C1(_12757_),
    .Y(_12888_));
 sky130_fd_sc_hd__nand3b_1 _46206_ (.A_N(_12867_),
    .B(_12877_),
    .C(_12888_),
    .Y(_12899_));
 sky130_fd_sc_hd__nand3_1 _46207_ (.A(_12119_),
    .B(_12856_),
    .C(_12899_),
    .Y(_12910_));
 sky130_fd_sc_hd__o21bai_1 _46208_ (.A1(_12823_),
    .A2(_12845_),
    .B1_N(_12867_),
    .Y(_12921_));
 sky130_fd_sc_hd__o31a_1 _46209_ (.A1(_08492_),
    .A2(_08503_),
    .A3(_08580_),
    .B1(_08536_),
    .X(_12932_));
 sky130_fd_sc_hd__o211ai_1 _46210_ (.A1(_12196_),
    .A2(_12163_),
    .B1(_12888_),
    .C1(_12877_),
    .Y(_12943_));
 sky130_fd_sc_hd__nand3_2 _46211_ (.A(_12921_),
    .B(_12932_),
    .C(_12943_),
    .Y(_12954_));
 sky130_fd_sc_hd__nand2_1 _46212_ (.A(_12910_),
    .B(_12954_),
    .Y(_12965_));
 sky130_fd_sc_hd__buf_1 _46213_ (.A(\delay_line[9][4] ),
    .X(_12976_));
 sky130_fd_sc_hd__buf_2 _46214_ (.A(_12976_),
    .X(_12987_));
 sky130_fd_sc_hd__nor2_1 _46215_ (.A(_25040_),
    .B(_12987_),
    .Y(_12998_));
 sky130_fd_sc_hd__and2_1 _46216_ (.A(_25040_),
    .B(_12987_),
    .X(_13009_));
 sky130_fd_sc_hd__nor2_1 _46217_ (.A(_12998_),
    .B(_13009_),
    .Y(_13020_));
 sky130_fd_sc_hd__nand2_2 _46218_ (.A(_25292_),
    .B(\delay_line[12][2] ),
    .Y(_13031_));
 sky130_fd_sc_hd__clkbuf_2 _46219_ (.A(net413),
    .X(_13042_));
 sky130_fd_sc_hd__o21ba_1 _46220_ (.A1(_08470_),
    .A2(_13031_),
    .B1_N(_13042_),
    .X(_13053_));
 sky130_fd_sc_hd__and4b_1 _46221_ (.A_N(_12152_),
    .B(_13042_),
    .C(_25292_),
    .D(_02414_),
    .X(_13064_));
 sky130_fd_sc_hd__nor2_1 _46222_ (.A(_13053_),
    .B(_13064_),
    .Y(_13075_));
 sky130_fd_sc_hd__or2_1 _46223_ (.A(_13020_),
    .B(_13075_),
    .X(_13086_));
 sky130_fd_sc_hd__or4_1 _46224_ (.A(_12998_),
    .B(_13009_),
    .C(_13053_),
    .D(_13064_),
    .X(_13097_));
 sky130_fd_sc_hd__and4b_1 _46225_ (.A_N(_08437_),
    .B(_08481_),
    .C(_23238_),
    .D(_25292_),
    .X(_13108_));
 sky130_fd_sc_hd__and3_1 _46226_ (.A(_13086_),
    .B(_13097_),
    .C(_13108_),
    .X(_13119_));
 sky130_fd_sc_hd__a21oi_1 _46227_ (.A1(_13086_),
    .A2(_13097_),
    .B1(_13108_),
    .Y(_13130_));
 sky130_fd_sc_hd__nor2_1 _46228_ (.A(_13119_),
    .B(_13130_),
    .Y(_13141_));
 sky130_fd_sc_hd__and3_1 _46229_ (.A(_08723_),
    .B(_08745_),
    .C(_13141_),
    .X(_13152_));
 sky130_fd_sc_hd__a21oi_1 _46230_ (.A1(_08723_),
    .A2(_08745_),
    .B1(_13141_),
    .Y(_13163_));
 sky130_fd_sc_hd__nor2_1 _46231_ (.A(_13152_),
    .B(_13163_),
    .Y(_13174_));
 sky130_fd_sc_hd__nand2_1 _46232_ (.A(_12965_),
    .B(_13174_),
    .Y(_13185_));
 sky130_fd_sc_hd__a31o_1 _46233_ (.A1(_08613_),
    .A2(_08624_),
    .A3(_08635_),
    .B1(_08800_),
    .X(_13196_));
 sky130_fd_sc_hd__and2_1 _46234_ (.A(_08811_),
    .B(_13196_),
    .X(_13207_));
 sky130_fd_sc_hd__o211ai_1 _46235_ (.A1(_13152_),
    .A2(_13163_),
    .B1(_12910_),
    .C1(_12954_),
    .Y(_13218_));
 sky130_fd_sc_hd__nand3_1 _46236_ (.A(_13185_),
    .B(_13207_),
    .C(_13218_),
    .Y(_13229_));
 sky130_fd_sc_hd__clkbuf_2 _46237_ (.A(_13229_),
    .X(_13240_));
 sky130_fd_sc_hd__nand2_1 _46238_ (.A(_12108_),
    .B(_13240_),
    .Y(_13251_));
 sky130_fd_sc_hd__nand2_1 _46239_ (.A(_12954_),
    .B(_13174_),
    .Y(_13262_));
 sky130_fd_sc_hd__and3_1 _46240_ (.A(_12119_),
    .B(_12856_),
    .C(_12899_),
    .X(_13273_));
 sky130_fd_sc_hd__nand2_1 _46241_ (.A(_08811_),
    .B(_13196_),
    .Y(_13284_));
 sky130_fd_sc_hd__o21ai_1 _46242_ (.A1(_13152_),
    .A2(_13163_),
    .B1(_12965_),
    .Y(_13295_));
 sky130_fd_sc_hd__o211a_2 _46243_ (.A1(_13262_),
    .A2(_13273_),
    .B1(_13284_),
    .C1(_13295_),
    .X(_13306_));
 sky130_fd_sc_hd__a21boi_1 _46244_ (.A1(_08866_),
    .A2(_09118_),
    .B1_N(_08833_),
    .Y(_13317_));
 sky130_fd_sc_hd__inv_2 _46245_ (.A(_13317_),
    .Y(_13328_));
 sky130_fd_sc_hd__o211ai_2 _46246_ (.A1(_13262_),
    .A2(_13273_),
    .B1(_13284_),
    .C1(_13295_),
    .Y(_13339_));
 sky130_fd_sc_hd__nand2_1 _46247_ (.A(_13339_),
    .B(_13229_),
    .Y(_13350_));
 sky130_fd_sc_hd__xnor2_1 _46248_ (.A(_09064_),
    .B(_12097_),
    .Y(_13361_));
 sky130_fd_sc_hd__nand2_1 _46249_ (.A(_13350_),
    .B(_13361_),
    .Y(_13372_));
 sky130_fd_sc_hd__o211ai_4 _46250_ (.A1(_13251_),
    .A2(_13306_),
    .B1(_13328_),
    .C1(_13372_),
    .Y(_13383_));
 sky130_fd_sc_hd__a21o_1 _46251_ (.A1(_13339_),
    .A2(_13240_),
    .B1(_13361_),
    .X(_13394_));
 sky130_fd_sc_hd__nand3_1 _46252_ (.A(_13339_),
    .B(_13240_),
    .C(_13361_),
    .Y(_13405_));
 sky130_fd_sc_hd__nand3_1 _46253_ (.A(_13394_),
    .B(_13317_),
    .C(_13405_),
    .Y(_13416_));
 sky130_fd_sc_hd__clkbuf_2 _46254_ (.A(_13416_),
    .X(_13427_));
 sky130_fd_sc_hd__a21oi_1 _46255_ (.A1(_03271_),
    .A2(_09108_),
    .B1(_09086_),
    .Y(_13438_));
 sky130_fd_sc_hd__clkbuf_2 _46256_ (.A(\delay_line[6][4] ),
    .X(_13449_));
 sky130_fd_sc_hd__inv_2 _46257_ (.A(_13449_),
    .Y(_13460_));
 sky130_fd_sc_hd__nand2_1 _46258_ (.A(_22974_),
    .B(_13460_),
    .Y(_13471_));
 sky130_fd_sc_hd__nand2_2 _46259_ (.A(_23018_),
    .B(_13449_),
    .Y(_13482_));
 sky130_fd_sc_hd__a31o_1 _46260_ (.A1(_11899_),
    .A2(_09020_),
    .A3(_00106_),
    .B1(_08998_),
    .X(_13493_));
 sky130_fd_sc_hd__nand3_1 _46261_ (.A(_13471_),
    .B(_13482_),
    .C(_13493_),
    .Y(_13504_));
 sky130_fd_sc_hd__a221o_1 _46262_ (.A1(_00117_),
    .A2(_11767_),
    .B1(_13471_),
    .B2(_13482_),
    .C1(_08998_),
    .X(_13515_));
 sky130_fd_sc_hd__and3_1 _46263_ (.A(_13504_),
    .B(_09239_),
    .C(_13515_),
    .X(_13526_));
 sky130_fd_sc_hd__o2bb2a_1 _46264_ (.A1_N(_13515_),
    .A2_N(_13504_),
    .B1(_09228_),
    .B2(_03227_),
    .X(_13537_));
 sky130_fd_sc_hd__and2b_1 _46265_ (.A_N(\delay_line[5][4] ),
    .B(\delay_line[5][3] ),
    .X(_13548_));
 sky130_fd_sc_hd__buf_1 _46266_ (.A(\delay_line[5][4] ),
    .X(_13559_));
 sky130_fd_sc_hd__and2b_1 _46267_ (.A_N(\delay_line[5][3] ),
    .B(_13559_),
    .X(_13570_));
 sky130_fd_sc_hd__o221ai_4 _46268_ (.A1(_03579_),
    .A2(_09459_),
    .B1(_13548_),
    .B2(_13570_),
    .C1(net431),
    .Y(_13581_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46269_ (.A(\delay_line[3][4] ),
    .X(_13592_));
 sky130_fd_sc_hd__xor2_1 _46270_ (.A(net431),
    .B(_13592_),
    .X(_13603_));
 sky130_fd_sc_hd__or2b_1 _46271_ (.A(_09459_),
    .B_N(_13559_),
    .X(_13614_));
 sky130_fd_sc_hd__o21ai_1 _46272_ (.A1(_03579_),
    .A2(_09459_),
    .B1(net431),
    .Y(_13625_));
 sky130_fd_sc_hd__nand3b_1 _46273_ (.A_N(_13548_),
    .B(_13614_),
    .C(_13625_),
    .Y(_13636_));
 sky130_fd_sc_hd__and3_1 _46274_ (.A(_13581_),
    .B(_13603_),
    .C(_13636_),
    .X(_13647_));
 sky130_fd_sc_hd__a21oi_1 _46275_ (.A1(_13636_),
    .A2(_13581_),
    .B1(_13603_),
    .Y(_13658_));
 sky130_fd_sc_hd__o21ai_1 _46276_ (.A1(_22897_),
    .A2(_24809_),
    .B1(_03414_),
    .Y(_13669_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46277_ (.A(\delay_line[6][1] ),
    .X(_13680_));
 sky130_fd_sc_hd__or3_1 _46278_ (.A(_22897_),
    .B(_13680_),
    .C(_03403_),
    .X(_13691_));
 sky130_fd_sc_hd__nand2_1 _46279_ (.A(_13669_),
    .B(_13691_),
    .Y(_13702_));
 sky130_fd_sc_hd__o21ai_1 _46280_ (.A1(_13647_),
    .A2(_13658_),
    .B1(_13702_),
    .Y(_13713_));
 sky130_fd_sc_hd__a21o_1 _46281_ (.A1(_13636_),
    .A2(_13581_),
    .B1(_13603_),
    .X(_13724_));
 sky130_fd_sc_hd__nand4b_2 _46282_ (.A_N(_13647_),
    .B(_13724_),
    .C(_13669_),
    .D(_13691_),
    .Y(_13735_));
 sky130_fd_sc_hd__and3_1 _46283_ (.A(_13713_),
    .B(_13735_),
    .C(net239),
    .X(_13746_));
 sky130_fd_sc_hd__a21oi_1 _46284_ (.A1(_13713_),
    .A2(_13735_),
    .B1(net239),
    .Y(_13757_));
 sky130_fd_sc_hd__or2b_1 _46285_ (.A(\delay_line[3][2] ),
    .B_N(net444),
    .X(_13768_));
 sky130_fd_sc_hd__inv_2 _46286_ (.A(\delay_line[2][4] ),
    .Y(_13779_));
 sky130_fd_sc_hd__nand2_1 _46287_ (.A(_13779_),
    .B(\delay_line[3][2] ),
    .Y(_13790_));
 sky130_fd_sc_hd__o2bb2ai_1 _46288_ (.A1_N(_13768_),
    .A2_N(_13790_),
    .B1(net437),
    .B2(_09316_),
    .Y(_13801_));
 sky130_fd_sc_hd__nand3b_2 _46289_ (.A_N(_09294_),
    .B(_13768_),
    .C(_13790_),
    .Y(_13812_));
 sky130_fd_sc_hd__nand4_2 _46290_ (.A(_13801_),
    .B(_03579_),
    .C(_13812_),
    .D(net436),
    .Y(_13823_));
 sky130_fd_sc_hd__inv_2 _46291_ (.A(net436),
    .Y(_13834_));
 sky130_fd_sc_hd__o2bb2ai_2 _46292_ (.A1_N(_13812_),
    .A2_N(_13801_),
    .B1(_24875_),
    .B2(_13834_),
    .Y(_13845_));
 sky130_fd_sc_hd__nand2_1 _46293_ (.A(_09294_),
    .B(_09327_),
    .Y(_13856_));
 sky130_fd_sc_hd__o2bb2ai_2 _46294_ (.A1_N(_13823_),
    .A2_N(_13845_),
    .B1(_03689_),
    .B2(_13856_),
    .Y(_13867_));
 sky130_fd_sc_hd__nand3_2 _46295_ (.A(_13845_),
    .B(_09338_),
    .C(_13823_),
    .Y(_13878_));
 sky130_fd_sc_hd__nand3_1 _46296_ (.A(_13867_),
    .B(_09514_),
    .C(_13878_),
    .Y(_13889_));
 sky130_fd_sc_hd__or2_1 _46297_ (.A(_09470_),
    .B(_09492_),
    .X(_13900_));
 sky130_fd_sc_hd__o2bb2ai_1 _46298_ (.A1_N(_13878_),
    .A2_N(_13867_),
    .B1(_09503_),
    .B2(_13900_),
    .Y(_13911_));
 sky130_fd_sc_hd__a2bb2o_1 _46299_ (.A1_N(_09283_),
    .A2_N(_09360_),
    .B1(_13889_),
    .B2(_13911_),
    .X(_13922_));
 sky130_fd_sc_hd__nor2_1 _46300_ (.A(_09283_),
    .B(_09360_),
    .Y(_13932_));
 sky130_fd_sc_hd__nand3_1 _46301_ (.A(_13911_),
    .B(_13932_),
    .C(_13889_),
    .Y(_13943_));
 sky130_fd_sc_hd__a2bb2o_1 _46302_ (.A1_N(_13746_),
    .A2_N(_13757_),
    .B1(_13922_),
    .B2(_13943_),
    .X(_13954_));
 sky130_fd_sc_hd__nor2_1 _46303_ (.A(_13746_),
    .B(_13757_),
    .Y(_13965_));
 sky130_fd_sc_hd__nand3_1 _46304_ (.A(_13965_),
    .B(_13922_),
    .C(_13943_),
    .Y(_13976_));
 sky130_fd_sc_hd__nand2_1 _46305_ (.A(_13954_),
    .B(_13976_),
    .Y(_13987_));
 sky130_fd_sc_hd__o21a_1 _46306_ (.A1(_13526_),
    .A2(_13537_),
    .B1(_13987_),
    .X(_13998_));
 sky130_fd_sc_hd__or2_1 _46307_ (.A(_13526_),
    .B(_13537_),
    .X(_14009_));
 sky130_fd_sc_hd__or2_1 _46308_ (.A(_14009_),
    .B(_13987_),
    .X(_14020_));
 sky130_fd_sc_hd__inv_2 _46309_ (.A(_14020_),
    .Y(_14031_));
 sky130_fd_sc_hd__or3_2 _46310_ (.A(_13438_),
    .B(_13998_),
    .C(_14031_),
    .X(_14042_));
 sky130_fd_sc_hd__o21ai_1 _46311_ (.A1(_13998_),
    .A2(_14031_),
    .B1(_13438_),
    .Y(_14053_));
 sky130_fd_sc_hd__nor2_1 _46312_ (.A(_09272_),
    .B(_09580_),
    .Y(_14064_));
 sky130_fd_sc_hd__a41o_1 _46313_ (.A1(_03458_),
    .A2(_03425_),
    .A3(_00117_),
    .A4(_09261_),
    .B1(_14064_),
    .X(_14075_));
 sky130_fd_sc_hd__a21oi_1 _46314_ (.A1(_14042_),
    .A2(_14053_),
    .B1(_14075_),
    .Y(_14086_));
 sky130_fd_sc_hd__and3_1 _46315_ (.A(_14075_),
    .B(_14042_),
    .C(_14053_),
    .X(_14097_));
 sky130_fd_sc_hd__nor2_1 _46316_ (.A(_14086_),
    .B(_14097_),
    .Y(_14108_));
 sky130_fd_sc_hd__a21oi_1 _46317_ (.A1(_13383_),
    .A2(_13427_),
    .B1(_14108_),
    .Y(_14119_));
 sky130_fd_sc_hd__nand2_1 _46318_ (.A(_14042_),
    .B(_14053_),
    .Y(_14130_));
 sky130_fd_sc_hd__and2_1 _46319_ (.A(_14075_),
    .B(_14130_),
    .X(_14141_));
 sky130_fd_sc_hd__nor2_1 _46320_ (.A(_14075_),
    .B(_14130_),
    .Y(_14152_));
 sky130_fd_sc_hd__o211a_1 _46321_ (.A1(_14141_),
    .A2(_14152_),
    .B1(_13383_),
    .C1(_13427_),
    .X(_14163_));
 sky130_fd_sc_hd__a32o_2 _46322_ (.A1(_07920_),
    .A2(_09129_),
    .A3(_09140_),
    .B1(_09206_),
    .B2(_09701_),
    .X(_14174_));
 sky130_fd_sc_hd__o21bai_4 _46323_ (.A1(_14119_),
    .A2(_14163_),
    .B1_N(_14174_),
    .Y(_14185_));
 sky130_fd_sc_hd__o21ai_2 _46324_ (.A1(_14141_),
    .A2(_14152_),
    .B1(_13427_),
    .Y(_14196_));
 sky130_fd_sc_hd__o211a_1 _46325_ (.A1(_13251_),
    .A2(_13306_),
    .B1(_13328_),
    .C1(_13372_),
    .X(_14207_));
 sky130_fd_sc_hd__o2bb2ai_2 _46326_ (.A1_N(_13383_),
    .A2_N(_13427_),
    .B1(_14086_),
    .B2(_14097_),
    .Y(_14218_));
 sky130_fd_sc_hd__o211ai_4 _46327_ (.A1(_14196_),
    .A2(_14207_),
    .B1(_14174_),
    .C1(_14218_),
    .Y(_14229_));
 sky130_fd_sc_hd__nand3_1 _46328_ (.A(_09899_),
    .B(_09910_),
    .C(_03711_),
    .Y(_14240_));
 sky130_fd_sc_hd__and4_1 _46329_ (.A(_03612_),
    .B(_09558_),
    .C(_09393_),
    .D(_22919_),
    .X(_14251_));
 sky130_fd_sc_hd__a21oi_2 _46330_ (.A1(_09415_),
    .A2(_09569_),
    .B1(_14251_),
    .Y(_14262_));
 sky130_fd_sc_hd__clkbuf_2 _46331_ (.A(\delay_line[1][3] ),
    .X(_14273_));
 sky130_fd_sc_hd__or2b_1 _46332_ (.A(_09745_),
    .B_N(_14273_),
    .X(_14284_));
 sky130_fd_sc_hd__or2b_1 _46333_ (.A(_14273_),
    .B_N(_09745_),
    .X(_14295_));
 sky130_fd_sc_hd__nand2_1 _46334_ (.A(_14284_),
    .B(_14295_),
    .Y(_14306_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46335_ (.A(net451),
    .X(_14317_));
 sky130_fd_sc_hd__nor2b_2 _46336_ (.A(_14317_),
    .B_N(_09767_),
    .Y(_14328_));
 sky130_fd_sc_hd__and2b_1 _46337_ (.A_N(_09767_),
    .B(net451),
    .X(_14339_));
 sky130_fd_sc_hd__o21ai_2 _46338_ (.A1(_14328_),
    .A2(_14339_),
    .B1(_24930_),
    .Y(_14350_));
 sky130_fd_sc_hd__inv_2 _46339_ (.A(\delay_line[2][1] ),
    .Y(_14361_));
 sky130_fd_sc_hd__or2b_1 _46340_ (.A(_14317_),
    .B_N(_09767_),
    .X(_14372_));
 sky130_fd_sc_hd__or2b_1 _46341_ (.A(_09767_),
    .B_N(_14317_),
    .X(_14383_));
 sky130_fd_sc_hd__nand3_2 _46342_ (.A(_14361_),
    .B(_14372_),
    .C(_14383_),
    .Y(_14394_));
 sky130_fd_sc_hd__a22oi_2 _46343_ (.A1(\delay_line[2][0] ),
    .A2(_14306_),
    .B1(_14350_),
    .B2(_14394_),
    .Y(_14405_));
 sky130_fd_sc_hd__and4bb_1 _46344_ (.A_N(\delay_line[1][0] ),
    .B_N(_14273_),
    .C(_03898_),
    .D(_00249_),
    .X(_14416_));
 sky130_fd_sc_hd__a21oi_2 _46345_ (.A1(_23414_),
    .A2(_00249_),
    .B1(_09778_),
    .Y(_14427_));
 sky130_fd_sc_hd__nor2_1 _46346_ (.A(_14416_),
    .B(_14427_),
    .Y(_14438_));
 sky130_fd_sc_hd__o2111ai_2 _46347_ (.A1(_09800_),
    .A2(_09778_),
    .B1(_14394_),
    .C1(_22875_),
    .D1(_14350_),
    .Y(_14449_));
 sky130_fd_sc_hd__nand3b_2 _46348_ (.A_N(_14405_),
    .B(_14438_),
    .C(_14449_),
    .Y(_14460_));
 sky130_fd_sc_hd__and4_1 _46349_ (.A(_14350_),
    .B(_22875_),
    .C(_14306_),
    .D(_14394_),
    .X(_14471_));
 sky130_fd_sc_hd__or2_1 _46350_ (.A(_14416_),
    .B(_14427_),
    .X(_14482_));
 sky130_fd_sc_hd__o21ai_2 _46351_ (.A1(_14471_),
    .A2(_14405_),
    .B1(_14482_),
    .Y(_14493_));
 sky130_fd_sc_hd__o211a_1 _46352_ (.A1(_09833_),
    .A2(_09877_),
    .B1(_14460_),
    .C1(_14493_),
    .X(_14504_));
 sky130_fd_sc_hd__a221oi_4 _46353_ (.A1(_09822_),
    .A2(_23414_),
    .B1(_14493_),
    .B2(_14460_),
    .C1(_09877_),
    .Y(_14515_));
 sky130_fd_sc_hd__nor4_1 _46354_ (.A(_03623_),
    .B(_09371_),
    .C(_14504_),
    .D(_14515_),
    .Y(_14526_));
 sky130_fd_sc_hd__buf_1 _46355_ (.A(_14504_),
    .X(_14537_));
 sky130_fd_sc_hd__o32a_1 _46356_ (.A1(_09393_),
    .A2(_09338_),
    .A3(_09349_),
    .B1(_14537_),
    .B2(_14515_),
    .X(_14548_));
 sky130_fd_sc_hd__o21ai_1 _46357_ (.A1(_14526_),
    .A2(_14548_),
    .B1(_09899_),
    .Y(_14559_));
 sky130_fd_sc_hd__o22ai_1 _46358_ (.A1(_09393_),
    .A2(_09371_),
    .B1(_14537_),
    .B2(_14515_),
    .Y(_14570_));
 sky130_fd_sc_hd__nand3b_1 _46359_ (.A_N(_14526_),
    .B(_14570_),
    .C(_09888_),
    .Y(_14581_));
 sky130_fd_sc_hd__nand2_1 _46360_ (.A(_14559_),
    .B(_14581_),
    .Y(_14592_));
 sky130_fd_sc_hd__xnor2_2 _46361_ (.A(_14262_),
    .B(_14592_),
    .Y(_14603_));
 sky130_fd_sc_hd__a21oi_1 _46362_ (.A1(_14240_),
    .A2(_09976_),
    .B1(_14603_),
    .Y(_14614_));
 sky130_fd_sc_hd__and3b_1 _46363_ (.A_N(_09921_),
    .B(_09976_),
    .C(_14603_),
    .X(_14625_));
 sky130_fd_sc_hd__and4bb_1 _46364_ (.A_N(_03271_),
    .B_N(_03282_),
    .C(_25139_),
    .D(_09602_),
    .X(_14636_));
 sky130_fd_sc_hd__o21ai_1 _46365_ (.A1(_09591_),
    .A2(_14636_),
    .B1(_09613_),
    .Y(_14647_));
 sky130_fd_sc_hd__o21ai_1 _46366_ (.A1(_14614_),
    .A2(_14625_),
    .B1(_14647_),
    .Y(_14658_));
 sky130_fd_sc_hd__or3_1 _46367_ (.A(_14647_),
    .B(_14614_),
    .C(_14625_),
    .X(_14669_));
 sky130_fd_sc_hd__nand2_1 _46368_ (.A(_14658_),
    .B(_14669_),
    .Y(_14680_));
 sky130_fd_sc_hd__xor2_2 _46369_ (.A(_09987_),
    .B(_14680_),
    .X(_14691_));
 sky130_fd_sc_hd__a21oi_2 _46370_ (.A1(_14185_),
    .A2(_14229_),
    .B1(_14691_),
    .Y(_14702_));
 sky130_fd_sc_hd__a31oi_1 _46371_ (.A1(_09657_),
    .A2(_09668_),
    .A3(_09679_),
    .B1(_10229_),
    .Y(_14713_));
 sky130_fd_sc_hd__a21oi_2 _46372_ (.A1(_09723_),
    .A2(_09712_),
    .B1(_14713_),
    .Y(_14724_));
 sky130_fd_sc_hd__a31o_1 _46373_ (.A1(_14185_),
    .A2(_14229_),
    .A3(_14691_),
    .B1(_14724_),
    .X(_14735_));
 sky130_fd_sc_hd__o211ai_1 _46374_ (.A1(_14141_),
    .A2(_14152_),
    .B1(_13383_),
    .C1(_13427_),
    .Y(_14746_));
 sky130_fd_sc_hd__a21oi_2 _46375_ (.A1(_14218_),
    .A2(_14746_),
    .B1(_14174_),
    .Y(_14757_));
 sky130_fd_sc_hd__o211a_2 _46376_ (.A1(_14196_),
    .A2(_14207_),
    .B1(_14174_),
    .C1(_14218_),
    .X(_14768_));
 sky130_fd_sc_hd__inv_2 _46377_ (.A(_09987_),
    .Y(_14779_));
 sky130_fd_sc_hd__xor2_1 _46378_ (.A(_14779_),
    .B(_14680_),
    .X(_14789_));
 sky130_fd_sc_hd__o21bai_1 _46379_ (.A1(_14757_),
    .A2(_14768_),
    .B1_N(_14789_),
    .Y(_14800_));
 sky130_fd_sc_hd__nand3_1 _46380_ (.A(_14185_),
    .B(_14229_),
    .C(_14789_),
    .Y(_14811_));
 sky130_fd_sc_hd__nand3_2 _46381_ (.A(_14800_),
    .B(_14724_),
    .C(_14811_),
    .Y(_14822_));
 sky130_fd_sc_hd__o21ai_1 _46382_ (.A1(_14702_),
    .A2(_14735_),
    .B1(_14822_),
    .Y(_14833_));
 sky130_fd_sc_hd__o21ai_4 _46383_ (.A1(_03975_),
    .A2(_10020_),
    .B1(_09998_),
    .Y(_14844_));
 sky130_fd_sc_hd__inv_2 _46384_ (.A(_14844_),
    .Y(_14855_));
 sky130_fd_sc_hd__nand2_1 _46385_ (.A(_14833_),
    .B(_14855_),
    .Y(_14866_));
 sky130_fd_sc_hd__o211ai_2 _46386_ (.A1(_14702_),
    .A2(_14735_),
    .B1(_14822_),
    .C1(_14844_),
    .Y(_14877_));
 sky130_fd_sc_hd__a32o_1 _46387_ (.A1(net99),
    .A2(_10163_),
    .A3(_10174_),
    .B1(_10152_),
    .B2(_04052_),
    .X(_14888_));
 sky130_fd_sc_hd__a21oi_4 _46388_ (.A1(_14866_),
    .A2(_14877_),
    .B1(_14888_),
    .Y(_14899_));
 sky130_fd_sc_hd__a32oi_4 _46389_ (.A1(net99),
    .A2(_10163_),
    .A3(_10174_),
    .B1(_10152_),
    .B2(_04052_),
    .Y(_14910_));
 sky130_fd_sc_hd__a31oi_1 _46390_ (.A1(_14185_),
    .A2(_14229_),
    .A3(_14691_),
    .B1(_14724_),
    .Y(_14921_));
 sky130_fd_sc_hd__o21ai_1 _46391_ (.A1(_14757_),
    .A2(_14768_),
    .B1(_14789_),
    .Y(_14932_));
 sky130_fd_sc_hd__nand2_1 _46392_ (.A(_14921_),
    .B(_14932_),
    .Y(_14943_));
 sky130_fd_sc_hd__a21oi_2 _46393_ (.A1(_14822_),
    .A2(_14943_),
    .B1(_14844_),
    .Y(_14954_));
 sky130_fd_sc_hd__o211a_2 _46394_ (.A1(_14702_),
    .A2(_14735_),
    .B1(_14822_),
    .C1(_14844_),
    .X(_14965_));
 sky130_fd_sc_hd__nor3_2 _46395_ (.A(_14910_),
    .B(_14954_),
    .C(_14965_),
    .Y(_14976_));
 sky130_fd_sc_hd__o21ai_1 _46396_ (.A1(_14899_),
    .A2(_14976_),
    .B1(_10394_),
    .Y(_14987_));
 sky130_fd_sc_hd__o21ai_2 _46397_ (.A1(_14954_),
    .A2(_14965_),
    .B1(_14910_),
    .Y(_14998_));
 sky130_fd_sc_hd__nand2_2 _46398_ (.A(_14998_),
    .B(_10328_),
    .Y(_15009_));
 sky130_fd_sc_hd__and2_4 _46399_ (.A(\delay_line[23][4] ),
    .B(_10339_),
    .X(_15020_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46400_ (.A(\delay_line[23][4] ),
    .X(_15031_));
 sky130_fd_sc_hd__nor2_1 _46401_ (.A(_15031_),
    .B(_10339_),
    .Y(_15042_));
 sky130_fd_sc_hd__nor2_2 _46402_ (.A(_15020_),
    .B(_15042_),
    .Y(_15053_));
 sky130_fd_sc_hd__nand3_2 _46403_ (.A(_14987_),
    .B(_15009_),
    .C(_15053_),
    .Y(_15064_));
 sky130_fd_sc_hd__a21o_1 _46404_ (.A1(_14833_),
    .A2(_14855_),
    .B1(_14910_),
    .X(_15075_));
 sky130_fd_sc_hd__o211ai_4 _46405_ (.A1(_14965_),
    .A2(_15075_),
    .B1(_14998_),
    .C1(_10394_),
    .Y(_15086_));
 sky130_fd_sc_hd__o21ai_1 _46406_ (.A1(_14899_),
    .A2(_14976_),
    .B1(_10328_),
    .Y(_15097_));
 sky130_fd_sc_hd__o211ai_4 _46407_ (.A1(_15020_),
    .A2(_15042_),
    .B1(_15086_),
    .C1(_15097_),
    .Y(_15108_));
 sky130_fd_sc_hd__o211a_2 _46408_ (.A1(_11658_),
    .A2(_05766_),
    .B1(_15064_),
    .C1(_15108_),
    .X(_15119_));
 sky130_fd_sc_hd__a21o_1 _46409_ (.A1(_05755_),
    .A2(_05678_),
    .B1(_11658_),
    .X(_15130_));
 sky130_fd_sc_hd__a21oi_1 _46410_ (.A1(_15064_),
    .A2(_15108_),
    .B1(_15130_),
    .Y(_15141_));
 sky130_fd_sc_hd__nand2_1 _46411_ (.A(_10416_),
    .B(_10405_),
    .Y(_15152_));
 sky130_fd_sc_hd__nand2_2 _46412_ (.A(_04579_),
    .B(_10339_),
    .Y(_15163_));
 sky130_fd_sc_hd__a21oi_1 _46413_ (.A1(_15152_),
    .A2(_15163_),
    .B1(_10350_),
    .Y(_15174_));
 sky130_fd_sc_hd__o21bai_4 _46414_ (.A1(_15119_),
    .A2(_15141_),
    .B1_N(_15174_),
    .Y(_15185_));
 sky130_fd_sc_hd__o211ai_4 _46415_ (.A1(_11658_),
    .A2(_05766_),
    .B1(_15064_),
    .C1(_15108_),
    .Y(_15196_));
 sky130_fd_sc_hd__a21o_1 _46416_ (.A1(_15064_),
    .A2(_15108_),
    .B1(_15130_),
    .X(_15207_));
 sky130_fd_sc_hd__nand3_1 _46417_ (.A(_15196_),
    .B(_15207_),
    .C(_15174_),
    .Y(_15218_));
 sky130_fd_sc_hd__buf_2 _46418_ (.A(_15218_),
    .X(_15229_));
 sky130_fd_sc_hd__and2b_1 _46419_ (.A_N(_06063_),
    .B(_05788_),
    .X(_15240_));
 sky130_fd_sc_hd__nor2_1 _46420_ (.A(net156),
    .B(_15240_),
    .Y(_15251_));
 sky130_fd_sc_hd__a21boi_1 _46421_ (.A1(_15185_),
    .A2(_15229_),
    .B1_N(_15251_),
    .Y(_15262_));
 sky130_fd_sc_hd__o211a_2 _46422_ (.A1(net156),
    .A2(_15240_),
    .B1(_15185_),
    .C1(_15229_),
    .X(_15273_));
 sky130_fd_sc_hd__a31o_1 _46423_ (.A1(_10459_),
    .A2(_10383_),
    .A3(_10426_),
    .B1(_10536_),
    .X(_15284_));
 sky130_fd_sc_hd__o21bai_4 _46424_ (.A1(_15262_),
    .A2(_15273_),
    .B1_N(_15284_),
    .Y(_15295_));
 sky130_fd_sc_hd__nand2_1 _46425_ (.A(_15185_),
    .B(_15218_),
    .Y(_15306_));
 sky130_fd_sc_hd__nand2_2 _46426_ (.A(_15306_),
    .B(_15251_),
    .Y(_15317_));
 sky130_fd_sc_hd__o211ai_4 _46427_ (.A1(net156),
    .A2(_15240_),
    .B1(_15185_),
    .C1(_15229_),
    .Y(_15328_));
 sky130_fd_sc_hd__o211ai_4 _46428_ (.A1(_10437_),
    .A2(_10536_),
    .B1(_15317_),
    .C1(_15328_),
    .Y(_15339_));
 sky130_fd_sc_hd__o21a_1 _46429_ (.A1(_04656_),
    .A2(_10580_),
    .B1(_11636_),
    .X(_15350_));
 sky130_fd_sc_hd__a21oi_2 _46430_ (.A1(_15295_),
    .A2(_15339_),
    .B1(_15350_),
    .Y(_15361_));
 sky130_fd_sc_hd__and3_1 _46431_ (.A(_15295_),
    .B(_15339_),
    .C(_15350_),
    .X(_15372_));
 sky130_fd_sc_hd__buf_1 _46432_ (.A(_04579_),
    .X(_15383_));
 sky130_fd_sc_hd__inv_2 _46433_ (.A(_15383_),
    .Y(_15394_));
 sky130_fd_sc_hd__o21ai_2 _46434_ (.A1(_15361_),
    .A2(_15372_),
    .B1(_15394_),
    .Y(_15405_));
 sky130_fd_sc_hd__o2111ai_4 _46435_ (.A1(_04656_),
    .A2(_10580_),
    .B1(_15295_),
    .C1(_15339_),
    .D1(_11636_),
    .Y(_15416_));
 sky130_fd_sc_hd__buf_2 _46436_ (.A(_15383_),
    .X(_15427_));
 sky130_fd_sc_hd__nand3b_2 _46437_ (.A_N(_15361_),
    .B(_15416_),
    .C(_15427_),
    .Y(_15438_));
 sky130_fd_sc_hd__nor2_1 _46438_ (.A(_06128_),
    .B(_06183_),
    .Y(_15449_));
 sky130_fd_sc_hd__a21boi_2 _46439_ (.A1(_15405_),
    .A2(_15438_),
    .B1_N(_15449_),
    .Y(_15460_));
 sky130_fd_sc_hd__o211a_1 _46440_ (.A1(_06128_),
    .A2(_06183_),
    .B1(_15405_),
    .C1(_15438_),
    .X(_15471_));
 sky130_fd_sc_hd__o22ai_2 _46441_ (.A1(_11625_),
    .A2(_11647_),
    .B1(_15460_),
    .B2(_15471_),
    .Y(_15482_));
 sky130_fd_sc_hd__nand2_1 _46442_ (.A(_15405_),
    .B(_15438_),
    .Y(_15493_));
 sky130_fd_sc_hd__nand2_1 _46443_ (.A(_15493_),
    .B(_15449_),
    .Y(_15504_));
 sky130_fd_sc_hd__o211ai_1 _46444_ (.A1(_06128_),
    .A2(_06183_),
    .B1(_15405_),
    .C1(_15438_),
    .Y(_15515_));
 sky130_fd_sc_hd__o31a_1 _46445_ (.A1(_04667_),
    .A2(_10569_),
    .A3(_10580_),
    .B1(_10646_),
    .X(_15526_));
 sky130_fd_sc_hd__nand3_1 _46446_ (.A(_15504_),
    .B(_15515_),
    .C(_15526_),
    .Y(_15537_));
 sky130_fd_sc_hd__or2_1 _46447_ (.A(_07810_),
    .B(_07799_),
    .X(_15548_));
 sky130_fd_sc_hd__nand3_1 _46448_ (.A(_06744_),
    .B(_07008_),
    .C(_07019_),
    .Y(_15559_));
 sky130_fd_sc_hd__clkbuf_2 _46449_ (.A(\delay_line[30][4] ),
    .X(_15569_));
 sky130_fd_sc_hd__clkbuf_2 _46450_ (.A(_15569_),
    .X(_15580_));
 sky130_fd_sc_hd__nor2_1 _46451_ (.A(_24622_),
    .B(_15580_),
    .Y(_15591_));
 sky130_fd_sc_hd__and2_2 _46452_ (.A(_24611_),
    .B(_15569_),
    .X(_15602_));
 sky130_fd_sc_hd__and4bb_1 _46453_ (.A_N(_15591_),
    .B_N(_15602_),
    .C(_22281_),
    .D(_06337_),
    .X(_15613_));
 sky130_fd_sc_hd__clkbuf_2 _46454_ (.A(_15613_),
    .X(_15624_));
 sky130_fd_sc_hd__o2bb2a_1 _46455_ (.A1_N(_22292_),
    .A2_N(_06337_),
    .B1(_15591_),
    .B2(_15602_),
    .X(_15635_));
 sky130_fd_sc_hd__buf_1 _46456_ (.A(\delay_line[29][2] ),
    .X(_15646_));
 sky130_fd_sc_hd__nor3b_2 _46457_ (.A(_15624_),
    .B(_15635_),
    .C_N(_15646_),
    .Y(_15657_));
 sky130_fd_sc_hd__o21ba_1 _46458_ (.A1(_15624_),
    .A2(_15635_),
    .B1_N(_15646_),
    .X(_15668_));
 sky130_fd_sc_hd__o21ai_1 _46459_ (.A1(\delay_line[31][2] ),
    .A2(_06205_),
    .B1(\delay_line[31][1] ),
    .Y(_15679_));
 sky130_fd_sc_hd__a21oi_2 _46460_ (.A1(_00952_),
    .A2(_06216_),
    .B1(_15679_),
    .Y(_15690_));
 sky130_fd_sc_hd__inv_2 _46461_ (.A(\delay_line[31][2] ),
    .Y(_15701_));
 sky130_fd_sc_hd__clkbuf_2 _46462_ (.A(_15701_),
    .X(_15712_));
 sky130_fd_sc_hd__nor2_1 _46463_ (.A(_15712_),
    .B(_06260_),
    .Y(_15723_));
 sky130_fd_sc_hd__nor2_1 _46464_ (.A(_00952_),
    .B(_06216_),
    .Y(_15734_));
 sky130_fd_sc_hd__o21ba_1 _46465_ (.A1(_15723_),
    .A2(_15734_),
    .B1_N(_24578_),
    .X(_15745_));
 sky130_fd_sc_hd__a211oi_2 _46466_ (.A1(_24633_),
    .A2(_00974_),
    .B1(_15690_),
    .C1(_15745_),
    .Y(_15756_));
 sky130_fd_sc_hd__and4_1 _46467_ (.A(_06271_),
    .B(_00963_),
    .C(_24589_),
    .D(_22215_),
    .X(_15767_));
 sky130_fd_sc_hd__nor2_1 _46468_ (.A(net318),
    .B(\delay_line[31][3] ),
    .Y(_15778_));
 sky130_fd_sc_hd__buf_1 _46469_ (.A(net318),
    .X(_15789_));
 sky130_fd_sc_hd__nand2_1 _46470_ (.A(_15789_),
    .B(_06205_),
    .Y(_15800_));
 sky130_fd_sc_hd__nand3b_2 _46471_ (.A_N(_15778_),
    .B(_15800_),
    .C(\delay_line[31][2] ),
    .Y(_15811_));
 sky130_fd_sc_hd__and2_1 _46472_ (.A(_15789_),
    .B(_06205_),
    .X(_15822_));
 sky130_fd_sc_hd__o21ai_2 _46473_ (.A1(_15778_),
    .A2(_15822_),
    .B1(_15712_),
    .Y(_15833_));
 sky130_fd_sc_hd__a221oi_4 _46474_ (.A1(_00963_),
    .A2(_06216_),
    .B1(_15811_),
    .B2(_15833_),
    .C1(_15690_),
    .Y(_15844_));
 sky130_fd_sc_hd__o211a_1 _46475_ (.A1(_15723_),
    .A2(_15690_),
    .B1(_15811_),
    .C1(_15833_),
    .X(_15855_));
 sky130_fd_sc_hd__buf_1 _46476_ (.A(_15855_),
    .X(_15866_));
 sky130_fd_sc_hd__or4_1 _46477_ (.A(_15756_),
    .B(_15767_),
    .C(_15844_),
    .D(_15866_),
    .X(_15877_));
 sky130_fd_sc_hd__o22ai_2 _46478_ (.A1(_15756_),
    .A2(_15767_),
    .B1(_15844_),
    .B2(_15866_),
    .Y(_15888_));
 sky130_fd_sc_hd__o211a_1 _46479_ (.A1(_15657_),
    .A2(_15668_),
    .B1(_15877_),
    .C1(_15888_),
    .X(_15899_));
 sky130_fd_sc_hd__a211oi_2 _46480_ (.A1(_15877_),
    .A2(_15888_),
    .B1(_15657_),
    .C1(_15668_),
    .Y(_15910_));
 sky130_fd_sc_hd__inv_2 _46481_ (.A(\delay_line[28][2] ),
    .Y(_15921_));
 sky130_fd_sc_hd__and3b_1 _46482_ (.A_N(_06414_),
    .B(_01117_),
    .C(_24369_),
    .X(_15932_));
 sky130_fd_sc_hd__a21o_1 _46483_ (.A1(_15921_),
    .A2(_06425_),
    .B1(_15932_),
    .X(_15943_));
 sky130_fd_sc_hd__or3b_2 _46484_ (.A(_06436_),
    .B(_01117_),
    .C_N(_06414_),
    .X(_15954_));
 sky130_fd_sc_hd__clkbuf_2 _46485_ (.A(net327),
    .X(_15965_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46486_ (.A(_15965_),
    .X(_15976_));
 sky130_fd_sc_hd__nand3_2 _46487_ (.A(_15943_),
    .B(_15954_),
    .C(_15976_),
    .Y(_15987_));
 sky130_fd_sc_hd__a21o_1 _46488_ (.A1(_15943_),
    .A2(_15954_),
    .B1(_15976_),
    .X(_15998_));
 sky130_fd_sc_hd__buf_1 _46489_ (.A(\delay_line[26][3] ),
    .X(_16009_));
 sky130_fd_sc_hd__buf_2 _46490_ (.A(_16009_),
    .X(_16020_));
 sky130_fd_sc_hd__clkbuf_2 _46491_ (.A(_16020_),
    .X(_16031_));
 sky130_fd_sc_hd__buf_1 _46492_ (.A(\delay_line[27][4] ),
    .X(_16042_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46493_ (.A(_16042_),
    .X(_16053_));
 sky130_fd_sc_hd__nor2_1 _46494_ (.A(_01183_),
    .B(_16053_),
    .Y(_16064_));
 sky130_fd_sc_hd__and2_1 _46495_ (.A(\delay_line[27][2] ),
    .B(_16042_),
    .X(_16075_));
 sky130_fd_sc_hd__or3_1 _46496_ (.A(_06513_),
    .B(_16064_),
    .C(_16075_),
    .X(_16086_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46497_ (.A(_16086_),
    .X(_16097_));
 sky130_fd_sc_hd__buf_1 _46498_ (.A(_16097_),
    .X(_16108_));
 sky130_fd_sc_hd__a2bb2o_1 _46499_ (.A1_N(_16064_),
    .A2_N(_16075_),
    .B1(_24303_),
    .B2(_06491_),
    .X(_16119_));
 sky130_fd_sc_hd__a21oi_1 _46500_ (.A1(_16108_),
    .A2(_16119_),
    .B1(_06524_),
    .Y(_16130_));
 sky130_fd_sc_hd__o21ba_1 _46501_ (.A1(_16053_),
    .A2(_06579_),
    .B1_N(_16130_),
    .X(_16141_));
 sky130_fd_sc_hd__nand2_1 _46502_ (.A(_16031_),
    .B(_16141_),
    .Y(_16151_));
 sky130_fd_sc_hd__or2_1 _46503_ (.A(_16031_),
    .B(_16141_),
    .X(_16162_));
 sky130_fd_sc_hd__a22oi_4 _46504_ (.A1(_15987_),
    .A2(_15998_),
    .B1(_16151_),
    .B2(_16162_),
    .Y(_16173_));
 sky130_fd_sc_hd__and4_1 _46505_ (.A(_15987_),
    .B(_15998_),
    .C(_16151_),
    .D(_16162_),
    .X(_16184_));
 sky130_fd_sc_hd__a211o_2 _46506_ (.A1(_06557_),
    .A2(_06612_),
    .B1(_16173_),
    .C1(_16184_),
    .X(_16195_));
 sky130_fd_sc_hd__nand2_2 _46507_ (.A(_06568_),
    .B(_06546_),
    .Y(_16206_));
 sky130_fd_sc_hd__o221ai_4 _46508_ (.A1(_06480_),
    .A2(_16206_),
    .B1(_16173_),
    .B2(_16184_),
    .C1(_06612_),
    .Y(_16217_));
 sky130_fd_sc_hd__nand2_1 _46509_ (.A(_16195_),
    .B(_16217_),
    .Y(_16228_));
 sky130_fd_sc_hd__o21a_2 _46510_ (.A1(_15899_),
    .A2(_15910_),
    .B1(_16228_),
    .X(_16239_));
 sky130_fd_sc_hd__and4bb_4 _46511_ (.A_N(_15899_),
    .B_N(_15910_),
    .C(_16195_),
    .D(_16217_),
    .X(_16250_));
 sky130_fd_sc_hd__a211o_2 _46512_ (.A1(_07008_),
    .A2(_15559_),
    .B1(_16239_),
    .C1(_16250_),
    .X(_16261_));
 sky130_fd_sc_hd__o211ai_2 _46513_ (.A1(_16239_),
    .A2(_16250_),
    .B1(_07008_),
    .C1(_15559_),
    .Y(_16272_));
 sky130_fd_sc_hd__and2b_1 _46514_ (.A_N(_06656_),
    .B(_06678_),
    .X(_16283_));
 sky130_fd_sc_hd__a21boi_1 _46515_ (.A1(_16261_),
    .A2(_16272_),
    .B1_N(_16283_),
    .Y(_16294_));
 sky130_fd_sc_hd__nand3b_2 _46516_ (.A_N(_16283_),
    .B(_16261_),
    .C(_16272_),
    .Y(_16305_));
 sky130_fd_sc_hd__and2b_1 _46517_ (.A_N(_16294_),
    .B(_16305_),
    .X(_16316_));
 sky130_fd_sc_hd__inv_2 _46518_ (.A(\delay_line[18][3] ),
    .Y(_16327_));
 sky130_fd_sc_hd__buf_2 _46519_ (.A(_16327_),
    .X(_16338_));
 sky130_fd_sc_hd__clkbuf_2 _46520_ (.A(_16338_),
    .X(_16349_));
 sky130_fd_sc_hd__inv_2 _46521_ (.A(\delay_line[19][2] ),
    .Y(_16360_));
 sky130_fd_sc_hd__clkbuf_2 _46522_ (.A(_16360_),
    .X(_16371_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46523_ (.A(\delay_line[19][3] ),
    .X(_16382_));
 sky130_fd_sc_hd__and2b_1 _46524_ (.A_N(_07382_),
    .B(_16382_),
    .X(_16393_));
 sky130_fd_sc_hd__clkbuf_2 _46525_ (.A(_16393_),
    .X(_16404_));
 sky130_fd_sc_hd__nor2_1 _46526_ (.A(_16382_),
    .B(_16360_),
    .Y(_16415_));
 sky130_fd_sc_hd__or2_1 _46527_ (.A(_16404_),
    .B(_16415_),
    .X(_16426_));
 sky130_fd_sc_hd__a211o_2 _46528_ (.A1(_23962_),
    .A2(_16371_),
    .B1(_16426_),
    .C1(_01644_),
    .X(_16437_));
 sky130_fd_sc_hd__nand2_1 _46529_ (.A(_23962_),
    .B(_16371_),
    .Y(_16448_));
 sky130_fd_sc_hd__a2bb2o_1 _46530_ (.A1_N(_16404_),
    .A2_N(_16415_),
    .B1(_07426_),
    .B2(_16448_),
    .X(_16459_));
 sky130_fd_sc_hd__and3_1 _46531_ (.A(_16349_),
    .B(_16437_),
    .C(_16459_),
    .X(_16470_));
 sky130_fd_sc_hd__a21oi_4 _46532_ (.A1(_16437_),
    .A2(_16459_),
    .B1(_16349_),
    .Y(_16481_));
 sky130_fd_sc_hd__clkbuf_2 _46533_ (.A(_07569_),
    .X(_16492_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46534_ (.A(\delay_line[21][3] ),
    .X(_16503_));
 sky130_fd_sc_hd__nand2b_2 _46535_ (.A_N(_16503_),
    .B(net361),
    .Y(_16514_));
 sky130_fd_sc_hd__nand2b_2 _46536_ (.A_N(net361),
    .B(_16503_),
    .Y(_16525_));
 sky130_fd_sc_hd__o2111ai_4 _46537_ (.A1(_24006_),
    .A2(_07602_),
    .B1(_16492_),
    .C1(_16514_),
    .D1(_16525_),
    .Y(_16536_));
 sky130_fd_sc_hd__o21a_1 _46538_ (.A1(_24017_),
    .A2(_07602_),
    .B1(_16492_),
    .X(_16547_));
 sky130_fd_sc_hd__a21o_1 _46539_ (.A1(_16525_),
    .A2(_16514_),
    .B1(_16547_),
    .X(_16558_));
 sky130_fd_sc_hd__o211a_1 _46540_ (.A1(_16470_),
    .A2(_16481_),
    .B1(_16536_),
    .C1(_16558_),
    .X(_16568_));
 sky130_fd_sc_hd__a211oi_4 _46541_ (.A1(_16536_),
    .A2(_16558_),
    .B1(_16470_),
    .C1(_16481_),
    .Y(_16579_));
 sky130_fd_sc_hd__clkbuf_2 _46542_ (.A(\delay_line[16][3] ),
    .X(_16590_));
 sky130_fd_sc_hd__clkbuf_2 _46543_ (.A(_16590_),
    .X(_16601_));
 sky130_fd_sc_hd__clkbuf_2 _46544_ (.A(_16601_),
    .X(_16612_));
 sky130_fd_sc_hd__nor2_1 _46545_ (.A(_24138_),
    .B(_16612_),
    .Y(_16623_));
 sky130_fd_sc_hd__inv_2 _46546_ (.A(\delay_line[16][0] ),
    .Y(_16634_));
 sky130_fd_sc_hd__clkbuf_2 _46547_ (.A(_16634_),
    .X(_16645_));
 sky130_fd_sc_hd__buf_2 _46548_ (.A(\delay_line[16][3] ),
    .X(_16656_));
 sky130_fd_sc_hd__inv_2 _46549_ (.A(_16656_),
    .Y(_16667_));
 sky130_fd_sc_hd__nor2_1 _46550_ (.A(_16645_),
    .B(_16667_),
    .Y(_16678_));
 sky130_fd_sc_hd__inv_2 _46551_ (.A(net387),
    .Y(_16689_));
 sky130_fd_sc_hd__nand2_1 _46552_ (.A(_16689_),
    .B(_01787_),
    .Y(_16700_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46553_ (.A(_16700_),
    .X(_16711_));
 sky130_fd_sc_hd__inv_2 _46554_ (.A(\delay_line[15][2] ),
    .Y(_16722_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46555_ (.A(net387),
    .X(_16733_));
 sky130_fd_sc_hd__nand2_1 _46556_ (.A(_16722_),
    .B(_16733_),
    .Y(_16744_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46557_ (.A(_16744_),
    .X(_16755_));
 sky130_fd_sc_hd__nand2_1 _46558_ (.A(_16711_),
    .B(_16755_),
    .Y(_16766_));
 sky130_fd_sc_hd__buf_1 _46559_ (.A(_07074_),
    .X(_16777_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46560_ (.A(_16777_),
    .X(_16788_));
 sky130_fd_sc_hd__and2_1 _46561_ (.A(_24083_),
    .B(_16788_),
    .X(_16799_));
 sky130_fd_sc_hd__or3b_2 _46562_ (.A(_16766_),
    .B(_16799_),
    .C_N(_07140_),
    .X(_16810_));
 sky130_fd_sc_hd__buf_1 _46563_ (.A(net392),
    .X(_16821_));
 sky130_fd_sc_hd__buf_1 _46564_ (.A(_16821_),
    .X(_16832_));
 sky130_fd_sc_hd__buf_2 _46565_ (.A(_16832_),
    .X(_16843_));
 sky130_fd_sc_hd__nand2_1 _46566_ (.A(_24083_),
    .B(_16788_),
    .Y(_16854_));
 sky130_fd_sc_hd__a22o_1 _46567_ (.A1(_16711_),
    .A2(_16755_),
    .B1(_16854_),
    .B2(_07140_),
    .X(_16865_));
 sky130_fd_sc_hd__and3_1 _46568_ (.A(_16810_),
    .B(_16843_),
    .C(_16865_),
    .X(_16876_));
 sky130_fd_sc_hd__a21oi_2 _46569_ (.A1(_16865_),
    .A2(_16810_),
    .B1(_16843_),
    .Y(_16887_));
 sky130_fd_sc_hd__or4_4 _46570_ (.A(_16623_),
    .B(_16678_),
    .C(_16876_),
    .D(_16887_),
    .X(_16898_));
 sky130_fd_sc_hd__o22ai_4 _46571_ (.A1(_16623_),
    .A2(_16678_),
    .B1(_16876_),
    .B2(_16887_),
    .Y(_16908_));
 sky130_fd_sc_hd__a31o_1 _46572_ (.A1(_07184_),
    .A2(_07151_),
    .A3(_07162_),
    .B1(_07239_),
    .X(_16919_));
 sky130_fd_sc_hd__a21oi_4 _46573_ (.A1(_16898_),
    .A2(_16908_),
    .B1(_16919_),
    .Y(_16930_));
 sky130_fd_sc_hd__and3_4 _46574_ (.A(_16919_),
    .B(_16898_),
    .C(_16908_),
    .X(_16941_));
 sky130_fd_sc_hd__or4_2 _46575_ (.A(_16568_),
    .B(_16579_),
    .C(_16930_),
    .D(_16941_),
    .X(_16952_));
 sky130_fd_sc_hd__o22ai_2 _46576_ (.A1(_16568_),
    .A2(_16579_),
    .B1(_16930_),
    .B2(_16941_),
    .Y(_16963_));
 sky130_fd_sc_hd__a21o_1 _46577_ (.A1(_07656_),
    .A2(_07678_),
    .B1(net148),
    .X(_16974_));
 sky130_fd_sc_hd__a21oi_2 _46578_ (.A1(_16952_),
    .A2(_16963_),
    .B1(_16974_),
    .Y(_16985_));
 sky130_fd_sc_hd__and3_2 _46579_ (.A(_16974_),
    .B(_16952_),
    .C(_16963_),
    .X(_16996_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46580_ (.A(\delay_line[24][3] ),
    .X(_17007_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46581_ (.A(_17007_),
    .X(_17018_));
 sky130_fd_sc_hd__clkbuf_2 _46582_ (.A(_17018_),
    .X(_17029_));
 sky130_fd_sc_hd__clkbuf_2 _46583_ (.A(_17029_),
    .X(_17040_));
 sky130_fd_sc_hd__nor2_1 _46584_ (.A(_23698_),
    .B(_17040_),
    .Y(_17051_));
 sky130_fd_sc_hd__and2_1 _46585_ (.A(_23698_),
    .B(_17040_),
    .X(_17062_));
 sky130_fd_sc_hd__inv_2 _46586_ (.A(net354),
    .Y(_17073_));
 sky130_fd_sc_hd__buf_1 _46587_ (.A(_17073_),
    .X(_17084_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46588_ (.A(_17084_),
    .X(_17095_));
 sky130_fd_sc_hd__clkbuf_2 _46589_ (.A(_17095_),
    .X(_17106_));
 sky130_fd_sc_hd__o21ai_2 _46590_ (.A1(_17051_),
    .A2(_17062_),
    .B1(_17106_),
    .Y(_17117_));
 sky130_fd_sc_hd__or3_2 _46591_ (.A(_17106_),
    .B(_17051_),
    .C(_17062_),
    .X(_17128_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46592_ (.A(\delay_line[25][2] ),
    .X(_17139_));
 sky130_fd_sc_hd__buf_1 _46593_ (.A(_17139_),
    .X(_17150_));
 sky130_fd_sc_hd__o211a_1 _46594_ (.A1(_06777_),
    .A2(_06832_),
    .B1(_22369_),
    .C1(_17150_),
    .X(_17161_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46595_ (.A(_06766_),
    .X(_17171_));
 sky130_fd_sc_hd__buf_1 _46596_ (.A(_17171_),
    .X(_17182_));
 sky130_fd_sc_hd__and2_2 _46597_ (.A(_23731_),
    .B(_17182_),
    .X(_17193_));
 sky130_fd_sc_hd__buf_1 _46598_ (.A(\delay_line[25][4] ),
    .X(_17204_));
 sky130_fd_sc_hd__buf_2 _46599_ (.A(_17204_),
    .X(_17215_));
 sky130_fd_sc_hd__buf_1 _46600_ (.A(_01490_),
    .X(_17226_));
 sky130_fd_sc_hd__or2b_1 _46601_ (.A(_17215_),
    .B_N(_17226_),
    .X(_17237_));
 sky130_fd_sc_hd__buf_1 _46602_ (.A(_17204_),
    .X(_17248_));
 sky130_fd_sc_hd__or2b_1 _46603_ (.A(_01490_),
    .B_N(_17248_),
    .X(_17259_));
 sky130_fd_sc_hd__nand2_2 _46604_ (.A(_17237_),
    .B(_17259_),
    .Y(_17270_));
 sky130_fd_sc_hd__o21ai_4 _46605_ (.A1(_17161_),
    .A2(_17193_),
    .B1(_17270_),
    .Y(_17281_));
 sky130_fd_sc_hd__or3_4 _46606_ (.A(_17270_),
    .B(_17193_),
    .C(_17161_),
    .X(_17292_));
 sky130_fd_sc_hd__and4_1 _46607_ (.A(_17117_),
    .B(_17128_),
    .C(_17281_),
    .D(_17292_),
    .X(_17303_));
 sky130_fd_sc_hd__a22oi_4 _46608_ (.A1(_17117_),
    .A2(_17128_),
    .B1(_17281_),
    .B2(_17292_),
    .Y(_17314_));
 sky130_fd_sc_hd__o211a_1 _46609_ (.A1(_17303_),
    .A2(_17314_),
    .B1(_07547_),
    .C1(_07645_),
    .X(_17325_));
 sky130_fd_sc_hd__a211oi_2 _46610_ (.A1(_07547_),
    .A2(_07645_),
    .B1(_17303_),
    .C1(_17314_),
    .Y(_17336_));
 sky130_fd_sc_hd__a211oi_1 _46611_ (.A1(_06942_),
    .A2(_06997_),
    .B1(_17325_),
    .C1(_17336_),
    .Y(_17346_));
 sky130_fd_sc_hd__o221a_1 _46612_ (.A1(_06975_),
    .A2(_06986_),
    .B1(_17336_),
    .B2(_17325_),
    .C1(_06942_),
    .X(_17357_));
 sky130_fd_sc_hd__or2_1 _46613_ (.A(_17346_),
    .B(_17357_),
    .X(_17368_));
 sky130_fd_sc_hd__o21ai_1 _46614_ (.A1(_16985_),
    .A2(_16996_),
    .B1(_17368_),
    .Y(_17379_));
 sky130_fd_sc_hd__o21ai_1 _46615_ (.A1(_07052_),
    .A2(_07711_),
    .B1(_07722_),
    .Y(_17390_));
 sky130_fd_sc_hd__o31a_1 _46616_ (.A1(_17368_),
    .A2(_16985_),
    .A3(_16996_),
    .B1(_17390_),
    .X(_17401_));
 sky130_fd_sc_hd__or3_1 _46617_ (.A(_17368_),
    .B(_16985_),
    .C(_16996_),
    .X(_17412_));
 sky130_fd_sc_hd__a21oi_1 _46618_ (.A1(_17412_),
    .A2(_17379_),
    .B1(_17390_),
    .Y(_17423_));
 sky130_fd_sc_hd__a21oi_1 _46619_ (.A1(_17379_),
    .A2(_17401_),
    .B1(_17423_),
    .Y(_17434_));
 sky130_fd_sc_hd__xnor2_1 _46620_ (.A(_16316_),
    .B(_17434_),
    .Y(_17445_));
 sky130_fd_sc_hd__o21ai_1 _46621_ (.A1(_06733_),
    .A2(_07788_),
    .B1(_07777_),
    .Y(_17456_));
 sky130_fd_sc_hd__xnor2_1 _46622_ (.A(_17445_),
    .B(_17456_),
    .Y(_17467_));
 sky130_fd_sc_hd__o21ai_1 _46623_ (.A1(_06194_),
    .A2(_06722_),
    .B1(_06711_),
    .Y(_17477_));
 sky130_fd_sc_hd__o21ai_2 _46624_ (.A1(_06030_),
    .A2(_05964_),
    .B1(_05942_),
    .Y(_17488_));
 sky130_fd_sc_hd__nor2_1 _46625_ (.A(\delay_line[37][0] ),
    .B(\delay_line[37][2] ),
    .Y(_17499_));
 sky130_fd_sc_hd__nand2_1 _46626_ (.A(_05975_),
    .B(_04294_),
    .Y(_17510_));
 sky130_fd_sc_hd__nor2b_1 _46627_ (.A(\delay_line[37][2] ),
    .B_N(\delay_line[37][4] ),
    .Y(_17521_));
 sky130_fd_sc_hd__and2b_1 _46628_ (.A_N(\delay_line[37][4] ),
    .B(\delay_line[37][2] ),
    .X(_17532_));
 sky130_fd_sc_hd__nor2_1 _46629_ (.A(_17521_),
    .B(_17532_),
    .Y(_17543_));
 sky130_fd_sc_hd__a21oi_1 _46630_ (.A1(_06008_),
    .A2(_17510_),
    .B1(_17543_),
    .Y(_17554_));
 sky130_fd_sc_hd__and3_1 _46631_ (.A(_17543_),
    .B(_17510_),
    .C(_06008_),
    .X(_17564_));
 sky130_fd_sc_hd__a311oi_2 _46632_ (.A1(_05975_),
    .A2(_17499_),
    .A3(_06008_),
    .B1(_17554_),
    .C1(_17564_),
    .Y(_17575_));
 sky130_fd_sc_hd__and4b_1 _46633_ (.A_N(\delay_line[37][4] ),
    .B(_05975_),
    .C(_05997_),
    .D(_17499_),
    .X(_17586_));
 sky130_fd_sc_hd__clkbuf_2 _46634_ (.A(\delay_line[35][4] ),
    .X(_17597_));
 sky130_fd_sc_hd__nor2_1 _46635_ (.A(_17597_),
    .B(_05799_),
    .Y(_17608_));
 sky130_fd_sc_hd__nand2_1 _46636_ (.A(_17597_),
    .B(_05799_),
    .Y(_17619_));
 sky130_fd_sc_hd__nand3b_1 _46637_ (.A_N(_17608_),
    .B(_17619_),
    .C(_04327_),
    .Y(_17630_));
 sky130_fd_sc_hd__and2_1 _46638_ (.A(_17597_),
    .B(\delay_line[35][3] ),
    .X(_17641_));
 sky130_fd_sc_hd__o21bai_1 _46639_ (.A1(_17608_),
    .A2(_17641_),
    .B1_N(\delay_line[35][2] ),
    .Y(_17652_));
 sky130_fd_sc_hd__nand2_1 _46640_ (.A(_17630_),
    .B(_17652_),
    .Y(_17662_));
 sky130_fd_sc_hd__a21o_1 _46641_ (.A1(_05821_),
    .A2(_05843_),
    .B1(_17662_),
    .X(_17673_));
 sky130_fd_sc_hd__nand3_1 _46642_ (.A(_05821_),
    .B(_05843_),
    .C(_17662_),
    .Y(_17684_));
 sky130_fd_sc_hd__and2_2 _46643_ (.A(_17673_),
    .B(_17684_),
    .X(_17695_));
 sky130_fd_sc_hd__and3b_1 _46644_ (.A_N(_05887_),
    .B(_17695_),
    .C(_05920_),
    .X(_17705_));
 sky130_fd_sc_hd__and4b_2 _46645_ (.A_N(_05909_),
    .B(_04327_),
    .C(_05832_),
    .D(_22677_),
    .X(_17716_));
 sky130_fd_sc_hd__o21ba_1 _46646_ (.A1(_05887_),
    .A2(_17716_),
    .B1_N(_17695_),
    .X(_17727_));
 sky130_fd_sc_hd__or3_1 _46647_ (.A(net298),
    .B(_17705_),
    .C(_17727_),
    .X(_17737_));
 sky130_fd_sc_hd__o21ai_2 _46648_ (.A1(_17705_),
    .A2(_17727_),
    .B1(net298),
    .Y(_17748_));
 sky130_fd_sc_hd__a2bb2o_1 _46649_ (.A1_N(_17575_),
    .A2_N(_17586_),
    .B1(_17737_),
    .B2(_17748_),
    .X(_17758_));
 sky130_fd_sc_hd__or4bb_4 _46650_ (.A(_17575_),
    .B(_17586_),
    .C_N(_17737_),
    .D_N(_17748_),
    .X(_17765_));
 sky130_fd_sc_hd__and3_4 _46651_ (.A(_17488_),
    .B(_17758_),
    .C(_17765_),
    .X(_17767_));
 sky130_fd_sc_hd__a21oi_2 _46652_ (.A1(_17758_),
    .A2(_17765_),
    .B1(_17488_),
    .Y(_17768_));
 sky130_fd_sc_hd__buf_1 _46653_ (.A(\delay_line[40][4] ),
    .X(_17769_));
 sky130_fd_sc_hd__nor2_1 _46654_ (.A(_17769_),
    .B(_05711_),
    .Y(_17770_));
 sky130_fd_sc_hd__or2b_1 _46655_ (.A(\delay_line[40][2] ),
    .B_N(\delay_line[40][4] ),
    .X(_17771_));
 sky130_fd_sc_hd__and2b_1 _46656_ (.A_N(\delay_line[40][3] ),
    .B(\delay_line[40][4] ),
    .X(_17772_));
 sky130_fd_sc_hd__a21oi_1 _46657_ (.A1(_17771_),
    .A2(_05689_),
    .B1(_17772_),
    .Y(_17773_));
 sky130_fd_sc_hd__o21a_1 _46658_ (.A1(_17770_),
    .A2(_17773_),
    .B1(_22776_),
    .X(_17774_));
 sky130_fd_sc_hd__nor3_1 _46659_ (.A(_22776_),
    .B(_17770_),
    .C(_17773_),
    .Y(_17775_));
 sky130_fd_sc_hd__a311o_1 _46660_ (.A1(_05722_),
    .A2(_05700_),
    .A3(_05711_),
    .B1(_17774_),
    .C1(_17775_),
    .X(_17776_));
 sky130_fd_sc_hd__o21ai_1 _46661_ (.A1(_17774_),
    .A2(_17775_),
    .B1(_05733_),
    .Y(_17777_));
 sky130_fd_sc_hd__nor2_1 _46662_ (.A(_00458_),
    .B(net288),
    .Y(_17778_));
 sky130_fd_sc_hd__and2_1 _46663_ (.A(\delay_line[38][1] ),
    .B(net288),
    .X(_17779_));
 sky130_fd_sc_hd__buf_1 _46664_ (.A(_17779_),
    .X(_17780_));
 sky130_fd_sc_hd__and4bb_1 _46665_ (.A_N(_17778_),
    .B_N(_17780_),
    .C(\delay_line[38][0] ),
    .D(_05568_),
    .X(_17781_));
 sky130_fd_sc_hd__o2bb2a_1 _46666_ (.A1_N(_22721_),
    .A2_N(_05568_),
    .B1(_17778_),
    .B2(_17780_),
    .X(_17782_));
 sky130_fd_sc_hd__nor2_1 _46667_ (.A(_17781_),
    .B(_17782_),
    .Y(_17783_));
 sky130_fd_sc_hd__nand4_1 _46668_ (.A(\delay_line[39][0] ),
    .B(_00403_),
    .C(_04129_),
    .D(_05623_),
    .Y(_17784_));
 sky130_fd_sc_hd__a31o_1 _46669_ (.A1(_00392_),
    .A2(_04129_),
    .A3(_05623_),
    .B1(\delay_line[39][0] ),
    .X(_17785_));
 sky130_fd_sc_hd__o311a_1 _46670_ (.A1(_00403_),
    .A2(_04140_),
    .A3(_05634_),
    .B1(_17784_),
    .C1(_17785_),
    .X(_17786_));
 sky130_fd_sc_hd__and2_1 _46671_ (.A(\delay_line[39][4] ),
    .B(\delay_line[39][3] ),
    .X(_17787_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46672_ (.A(\delay_line[39][4] ),
    .X(_17788_));
 sky130_fd_sc_hd__nor2_1 _46673_ (.A(_17788_),
    .B(_05601_),
    .Y(_17789_));
 sky130_fd_sc_hd__or3b_1 _46674_ (.A(_17787_),
    .B(_17789_),
    .C_N(\delay_line[39][2] ),
    .X(_17790_));
 sky130_fd_sc_hd__o21bai_1 _46675_ (.A1(_17787_),
    .A2(_17789_),
    .B1_N(\delay_line[39][2] ),
    .Y(_17791_));
 sky130_fd_sc_hd__o21a_1 _46676_ (.A1(\delay_line[39][2] ),
    .A2(_05601_),
    .B1(\delay_line[39][1] ),
    .X(_17792_));
 sky130_fd_sc_hd__a21o_1 _46677_ (.A1(_04118_),
    .A2(_05601_),
    .B1(_17792_),
    .X(_17793_));
 sky130_fd_sc_hd__a21oi_1 _46678_ (.A1(_17790_),
    .A2(_17791_),
    .B1(_17793_),
    .Y(_17794_));
 sky130_fd_sc_hd__and3_2 _46679_ (.A(_17793_),
    .B(_17790_),
    .C(_17791_),
    .X(_17795_));
 sky130_fd_sc_hd__o21ba_1 _46680_ (.A1(_17794_),
    .A2(_17795_),
    .B1_N(_00392_),
    .X(_17796_));
 sky130_fd_sc_hd__nor3b_1 _46681_ (.A(_17794_),
    .B(_17795_),
    .C_N(_00392_),
    .Y(_17797_));
 sky130_fd_sc_hd__or2_1 _46682_ (.A(_17796_),
    .B(_17797_),
    .X(_17798_));
 sky130_fd_sc_hd__xnor2_1 _46683_ (.A(_17786_),
    .B(_17798_),
    .Y(_17799_));
 sky130_fd_sc_hd__and2_2 _46684_ (.A(_17783_),
    .B(_17799_),
    .X(_17800_));
 sky130_fd_sc_hd__nor2_1 _46685_ (.A(_17783_),
    .B(_17799_),
    .Y(_17801_));
 sky130_fd_sc_hd__nor2_1 _46686_ (.A(_17800_),
    .B(_17801_),
    .Y(_17802_));
 sky130_fd_sc_hd__a21oi_1 _46687_ (.A1(_17776_),
    .A2(_17777_),
    .B1(_17802_),
    .Y(_17803_));
 sky130_fd_sc_hd__and3_2 _46688_ (.A(_17802_),
    .B(_17777_),
    .C(_17776_),
    .X(_17804_));
 sky130_fd_sc_hd__nor2_1 _46689_ (.A(_17803_),
    .B(_17804_),
    .Y(_17805_));
 sky130_fd_sc_hd__o21ba_2 _46690_ (.A1(_17767_),
    .A2(_17768_),
    .B1_N(_17805_),
    .X(_17806_));
 sky130_fd_sc_hd__nor3b_4 _46691_ (.A(_17767_),
    .B(_17768_),
    .C_N(_17805_),
    .Y(_17807_));
 sky130_fd_sc_hd__inv_2 _46692_ (.A(_05359_),
    .Y(_17808_));
 sky130_fd_sc_hd__xor2_1 _46693_ (.A(\delay_line[34][0] ),
    .B(net308),
    .X(_17809_));
 sky130_fd_sc_hd__buf_1 _46694_ (.A(\delay_line[34][4] ),
    .X(_17810_));
 sky130_fd_sc_hd__nand2_1 _46695_ (.A(_02238_),
    .B(_17810_),
    .Y(_17811_));
 sky130_fd_sc_hd__clkbuf_2 _46696_ (.A(_17810_),
    .X(_17812_));
 sky130_fd_sc_hd__o211a_1 _46697_ (.A1(_02238_),
    .A2(_17812_),
    .B1(_05392_),
    .C1(net308),
    .X(_17813_));
 sky130_fd_sc_hd__and2_1 _46698_ (.A(net307),
    .B(_17810_),
    .X(_17814_));
 sky130_fd_sc_hd__nor2_1 _46699_ (.A(_02238_),
    .B(_17812_),
    .Y(_17815_));
 sky130_fd_sc_hd__o2bb2ai_1 _46700_ (.A1_N(_00601_),
    .A2_N(_05392_),
    .B1(_17814_),
    .B2(_17815_),
    .Y(_17816_));
 sky130_fd_sc_hd__a21boi_1 _46701_ (.A1(_17811_),
    .A2(_17813_),
    .B1_N(_17816_),
    .Y(_17817_));
 sky130_fd_sc_hd__xor2_1 _46702_ (.A(_17809_),
    .B(_17817_),
    .X(_17818_));
 sky130_fd_sc_hd__o211a_1 _46703_ (.A1(_02249_),
    .A2(_05414_),
    .B1(_17818_),
    .C1(_22611_),
    .X(_17819_));
 sky130_fd_sc_hd__o21a_1 _46704_ (.A1(_02260_),
    .A2(_05414_),
    .B1(_22622_),
    .X(_17820_));
 sky130_fd_sc_hd__nor2_1 _46705_ (.A(_17820_),
    .B(_17818_),
    .Y(_17821_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46706_ (.A(\delay_line[33][4] ),
    .X(_17822_));
 sky130_fd_sc_hd__clkbuf_2 _46707_ (.A(_17822_),
    .X(_17823_));
 sky130_fd_sc_hd__clkbuf_2 _46708_ (.A(_17823_),
    .X(_17824_));
 sky130_fd_sc_hd__clkbuf_2 _46709_ (.A(_17824_),
    .X(_17825_));
 sky130_fd_sc_hd__nor2_1 _46710_ (.A(_22545_),
    .B(_17825_),
    .Y(_17826_));
 sky130_fd_sc_hd__and2_1 _46711_ (.A(_22534_),
    .B(_17825_),
    .X(_17827_));
 sky130_fd_sc_hd__a21oi_1 _46712_ (.A1(_02106_),
    .A2(_05315_),
    .B1(\delay_line[32][0] ),
    .Y(_17828_));
 sky130_fd_sc_hd__o2bb2a_1 _46713_ (.A1_N(\delay_line[32][0] ),
    .A2_N(_05370_),
    .B1(_17828_),
    .B2(_24534_),
    .X(_17829_));
 sky130_fd_sc_hd__a31o_1 _46714_ (.A1(_02128_),
    .A2(_05315_),
    .A3(_24556_),
    .B1(_17829_),
    .X(_17830_));
 sky130_fd_sc_hd__clkbuf_2 _46715_ (.A(\delay_line[32][4] ),
    .X(_17831_));
 sky130_fd_sc_hd__buf_1 _46716_ (.A(\delay_line[32][4] ),
    .X(_17832_));
 sky130_fd_sc_hd__o21ai_1 _46717_ (.A1(_17832_),
    .A2(_05293_),
    .B1(\delay_line[32][2] ),
    .Y(_17833_));
 sky130_fd_sc_hd__a21o_1 _46718_ (.A1(_17831_),
    .A2(_05293_),
    .B1(_17833_),
    .X(_17834_));
 sky130_fd_sc_hd__and2_1 _46719_ (.A(_17832_),
    .B(\delay_line[32][3] ),
    .X(_17835_));
 sky130_fd_sc_hd__nor2_1 _46720_ (.A(_17831_),
    .B(_05293_),
    .Y(_17836_));
 sky130_fd_sc_hd__o21ai_1 _46721_ (.A1(_17835_),
    .A2(_17836_),
    .B1(_05216_),
    .Y(_17837_));
 sky130_fd_sc_hd__o21ai_1 _46722_ (.A1(\delay_line[32][2] ),
    .A2(_05293_),
    .B1(_24457_),
    .Y(_17838_));
 sky130_fd_sc_hd__o21ai_1 _46723_ (.A1(_05205_),
    .A2(_05249_),
    .B1(_17838_),
    .Y(_17839_));
 sky130_fd_sc_hd__a21oi_1 _46724_ (.A1(_17834_),
    .A2(_17837_),
    .B1(_17839_),
    .Y(_17840_));
 sky130_fd_sc_hd__and3_1 _46725_ (.A(_17839_),
    .B(_17834_),
    .C(_17837_),
    .X(_17841_));
 sky130_fd_sc_hd__or3_1 _46726_ (.A(_24534_),
    .B(_17840_),
    .C(_17841_),
    .X(_17842_));
 sky130_fd_sc_hd__o21ai_1 _46727_ (.A1(_17840_),
    .A2(_17841_),
    .B1(_24534_),
    .Y(_17843_));
 sky130_fd_sc_hd__nand2_1 _46728_ (.A(_17842_),
    .B(_17843_),
    .Y(_17844_));
 sky130_fd_sc_hd__xor2_1 _46729_ (.A(_17830_),
    .B(_17844_),
    .X(_17845_));
 sky130_fd_sc_hd__nor3b_1 _46730_ (.A(_17826_),
    .B(_17827_),
    .C_N(_17845_),
    .Y(_17846_));
 sky130_fd_sc_hd__inv_2 _46731_ (.A(_17846_),
    .Y(_17847_));
 sky130_fd_sc_hd__o21bai_1 _46732_ (.A1(_17826_),
    .A2(_17827_),
    .B1_N(_17845_),
    .Y(_17848_));
 sky130_fd_sc_hd__a2bb2o_1 _46733_ (.A1_N(_17819_),
    .A2_N(_17821_),
    .B1(_17847_),
    .B2(_17848_),
    .X(_17849_));
 sky130_fd_sc_hd__or4b_2 _46734_ (.A(_17819_),
    .B(_17821_),
    .C(_17846_),
    .D_N(_17848_),
    .X(_17850_));
 sky130_fd_sc_hd__nor3b_4 _46735_ (.A(_06348_),
    .B(_06359_),
    .C_N(net323),
    .Y(_17851_));
 sky130_fd_sc_hd__a211oi_2 _46736_ (.A1(_17849_),
    .A2(_17850_),
    .B1(_17851_),
    .C1(_06392_),
    .Y(_17852_));
 sky130_fd_sc_hd__o211a_1 _46737_ (.A1(_17851_),
    .A2(_06392_),
    .B1(_17849_),
    .C1(_17850_),
    .X(_17853_));
 sky130_fd_sc_hd__a2111oi_1 _46738_ (.A1(_05425_),
    .A2(_17808_),
    .B1(_05381_),
    .C1(_17852_),
    .D1(_17853_),
    .Y(_17854_));
 sky130_fd_sc_hd__a21oi_1 _46739_ (.A1(_17808_),
    .A2(_05425_),
    .B1(_05381_),
    .Y(_17855_));
 sky130_fd_sc_hd__o21ba_1 _46740_ (.A1(_17852_),
    .A2(_17853_),
    .B1_N(_17855_),
    .X(_17856_));
 sky130_fd_sc_hd__nor2_1 _46741_ (.A(net122),
    .B(_17856_),
    .Y(_17857_));
 sky130_fd_sc_hd__and3_1 _46742_ (.A(_17857_),
    .B(_05524_),
    .C(_05491_),
    .X(_17858_));
 sky130_fd_sc_hd__o2bb2a_1 _46743_ (.A1_N(_05491_),
    .A2_N(_05524_),
    .B1(net123),
    .B2(_17856_),
    .X(_17859_));
 sky130_fd_sc_hd__nor4_1 _46744_ (.A(_17806_),
    .B(net139),
    .C(_17858_),
    .D(_17859_),
    .Y(_17860_));
 sky130_fd_sc_hd__o22a_1 _46745_ (.A1(_17806_),
    .A2(net139),
    .B1(_17858_),
    .B2(_17859_),
    .X(_17861_));
 sky130_fd_sc_hd__nor2_1 _46746_ (.A(_17860_),
    .B(_17861_),
    .Y(_17862_));
 sky130_fd_sc_hd__xnor2_1 _46747_ (.A(_17477_),
    .B(_17862_),
    .Y(_17863_));
 sky130_fd_sc_hd__a21oi_1 _46748_ (.A1(_05546_),
    .A2(_06117_),
    .B1(_17863_),
    .Y(_17864_));
 sky130_fd_sc_hd__and3_1 _46749_ (.A(_05546_),
    .B(_06117_),
    .C(_17863_),
    .X(_17865_));
 sky130_fd_sc_hd__nor2_1 _46750_ (.A(_17864_),
    .B(_17865_),
    .Y(_17866_));
 sky130_fd_sc_hd__xnor2_1 _46751_ (.A(_17467_),
    .B(_17866_),
    .Y(_17867_));
 sky130_fd_sc_hd__a21oi_2 _46752_ (.A1(_15548_),
    .A2(_07843_),
    .B1(_17867_),
    .Y(_17868_));
 sky130_fd_sc_hd__o311a_1 _46753_ (.A1(_07821_),
    .A2(_06161_),
    .A3(_06183_),
    .B1(_17867_),
    .C1(_15548_),
    .X(_17869_));
 sky130_fd_sc_hd__or2_1 _46754_ (.A(_17868_),
    .B(_17869_),
    .X(_17870_));
 sky130_fd_sc_hd__nand3_2 _46755_ (.A(_15482_),
    .B(_15537_),
    .C(_17870_),
    .Y(_17871_));
 sky130_fd_sc_hd__o21ai_1 _46756_ (.A1(_15460_),
    .A2(_15471_),
    .B1(_15526_),
    .Y(_17872_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46757_ (.A(_15515_),
    .X(_17873_));
 sky130_fd_sc_hd__o211ai_1 _46758_ (.A1(_11625_),
    .A2(_11647_),
    .B1(_15504_),
    .C1(_17873_),
    .Y(_17874_));
 sky130_fd_sc_hd__nor2_1 _46759_ (.A(_17868_),
    .B(_17869_),
    .Y(_17875_));
 sky130_fd_sc_hd__nand3_1 _46760_ (.A(_17872_),
    .B(_17874_),
    .C(_17875_),
    .Y(_17876_));
 sky130_fd_sc_hd__o211a_1 _46761_ (.A1(_07865_),
    .A2(_10701_),
    .B1(_17871_),
    .C1(_17876_),
    .X(_17877_));
 sky130_fd_sc_hd__a21o_1 _46762_ (.A1(_07854_),
    .A2(_07876_),
    .B1(_10701_),
    .X(_17878_));
 sky130_fd_sc_hd__a21oi_1 _46763_ (.A1(_17871_),
    .A2(_17876_),
    .B1(_17878_),
    .Y(_17879_));
 sky130_fd_sc_hd__o22ai_1 _46764_ (.A1(_11592_),
    .A2(_11614_),
    .B1(_17877_),
    .B2(_17879_),
    .Y(_17880_));
 sky130_fd_sc_hd__a21o_1 _46765_ (.A1(_17871_),
    .A2(_17876_),
    .B1(_17878_),
    .X(_17881_));
 sky130_fd_sc_hd__nor2_1 _46766_ (.A(_11592_),
    .B(_11603_),
    .Y(_17882_));
 sky130_fd_sc_hd__o211ai_1 _46767_ (.A1(_07865_),
    .A2(_10701_),
    .B1(_17871_),
    .C1(_17876_),
    .Y(_17883_));
 sky130_fd_sc_hd__nand3_1 _46768_ (.A(_17881_),
    .B(_17882_),
    .C(_17883_),
    .Y(_17884_));
 sky130_fd_sc_hd__a22oi_1 _46769_ (.A1(_10734_),
    .A2(_11284_),
    .B1(_17880_),
    .B2(_17884_),
    .Y(_17885_));
 sky130_fd_sc_hd__nand4_1 _46770_ (.A(_10734_),
    .B(_11284_),
    .C(_17880_),
    .D(_17884_),
    .Y(_17886_));
 sky130_fd_sc_hd__or2b_1 _46771_ (.A(_17885_),
    .B_N(_17886_),
    .X(_17887_));
 sky130_fd_sc_hd__xnor2_1 _46772_ (.A(_11273_),
    .B(_17887_),
    .Y(_17888_));
 sky130_fd_sc_hd__nand3_1 _46773_ (.A(_11185_),
    .B(_11229_),
    .C(_17888_),
    .Y(_17889_));
 sky130_fd_sc_hd__a21o_1 _46774_ (.A1(_11185_),
    .A2(_11229_),
    .B1(_17888_),
    .X(_17890_));
 sky130_fd_sc_hd__a2bb2o_1 _46775_ (.A1_N(_11207_),
    .A2_N(_11218_),
    .B1(_17889_),
    .B2(_17890_),
    .X(_17891_));
 sky130_fd_sc_hd__nor2_1 _46776_ (.A(_11218_),
    .B(_11207_),
    .Y(_17892_));
 sky130_fd_sc_hd__nand3_1 _46777_ (.A(_17890_),
    .B(_17889_),
    .C(_17892_),
    .Y(_17893_));
 sky130_fd_sc_hd__and2_1 _46778_ (.A(_17891_),
    .B(_17893_),
    .X(_17894_));
 sky130_fd_sc_hd__clkbuf_1 _46779_ (.A(_17894_),
    .X(_00035_));
 sky130_fd_sc_hd__buf_1 _46780_ (.A(_23502_),
    .X(_17895_));
 sky130_fd_sc_hd__clkbuf_2 _46781_ (.A(_10339_),
    .X(_17896_));
 sky130_fd_sc_hd__clkbuf_2 _46782_ (.A(_17896_),
    .X(_17897_));
 sky130_fd_sc_hd__clkbuf_2 _46783_ (.A(_17897_),
    .X(_17898_));
 sky130_fd_sc_hd__and2b_1 _46784_ (.A_N(_17895_),
    .B(_17898_),
    .X(_17899_));
 sky130_fd_sc_hd__and2b_1 _46785_ (.A_N(_17898_),
    .B(_17895_),
    .X(_17900_));
 sky130_fd_sc_hd__nor2_2 _46786_ (.A(_15031_),
    .B(\delay_line[23][5] ),
    .Y(_17901_));
 sky130_fd_sc_hd__and2_1 _46787_ (.A(_15031_),
    .B(\delay_line[23][5] ),
    .X(_17902_));
 sky130_fd_sc_hd__clkbuf_4 _46788_ (.A(_17902_),
    .X(_17903_));
 sky130_fd_sc_hd__o22ai_2 _46789_ (.A1(_14965_),
    .A2(_15075_),
    .B1(_10394_),
    .B2(_14899_),
    .Y(_17904_));
 sky130_fd_sc_hd__buf_2 _46790_ (.A(_17904_),
    .X(_17905_));
 sky130_fd_sc_hd__clkbuf_2 _46791_ (.A(_17905_),
    .X(_17906_));
 sky130_fd_sc_hd__a21bo_1 _46792_ (.A1(_14779_),
    .A2(_14658_),
    .B1_N(_14669_),
    .X(_17907_));
 sky130_fd_sc_hd__a21o_1 _46793_ (.A1(_13416_),
    .A2(_14108_),
    .B1(_14207_),
    .X(_17908_));
 sky130_fd_sc_hd__nor2_2 _46794_ (.A(net414),
    .B(_11680_),
    .Y(_17909_));
 sky130_fd_sc_hd__inv_2 _46795_ (.A(net414),
    .Y(_17910_));
 sky130_fd_sc_hd__nor2_1 _46796_ (.A(net415),
    .B(_17910_),
    .Y(_17911_));
 sky130_fd_sc_hd__buf_1 _46797_ (.A(\delay_line[9][5] ),
    .X(_17912_));
 sky130_fd_sc_hd__clkbuf_2 _46798_ (.A(_17912_),
    .X(_17913_));
 sky130_fd_sc_hd__o21a_1 _46799_ (.A1(_17909_),
    .A2(_17911_),
    .B1(_17913_),
    .X(_17914_));
 sky130_fd_sc_hd__buf_2 _46800_ (.A(_17913_),
    .X(_17915_));
 sky130_fd_sc_hd__clkbuf_4 _46801_ (.A(_17915_),
    .X(_17916_));
 sky130_fd_sc_hd__nor3_1 _46802_ (.A(_17916_),
    .B(_17909_),
    .C(_17911_),
    .Y(_17917_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46803_ (.A(\delay_line[10][5] ),
    .X(_17918_));
 sky130_fd_sc_hd__buf_2 _46804_ (.A(_17918_),
    .X(_17919_));
 sky130_fd_sc_hd__and4_1 _46805_ (.A(_12174_),
    .B(_08470_),
    .C(_17919_),
    .D(_02414_),
    .X(_17920_));
 sky130_fd_sc_hd__clkbuf_4 _46806_ (.A(_17918_),
    .X(_17921_));
 sky130_fd_sc_hd__nor2_1 _46807_ (.A(_17921_),
    .B(_12163_),
    .Y(_17922_));
 sky130_fd_sc_hd__or3b_2 _46808_ (.A(_13031_),
    .B(_12152_),
    .C_N(_13042_),
    .X(_17923_));
 sky130_fd_sc_hd__or3_2 _46809_ (.A(_17920_),
    .B(_17922_),
    .C(_17923_),
    .X(_17924_));
 sky130_fd_sc_hd__buf_1 _46810_ (.A(_17920_),
    .X(_17925_));
 sky130_fd_sc_hd__o21ai_1 _46811_ (.A1(_17925_),
    .A2(_17922_),
    .B1(_17923_),
    .Y(_17926_));
 sky130_fd_sc_hd__a2bb2o_1 _46812_ (.A1_N(_17914_),
    .A2_N(net238),
    .B1(_17924_),
    .B2(_17926_),
    .X(_17927_));
 sky130_fd_sc_hd__or4bb_1 _46813_ (.A(_17914_),
    .B(net238),
    .C_N(_17924_),
    .D_N(_17926_),
    .X(_17928_));
 sky130_fd_sc_hd__clkbuf_2 _46814_ (.A(_17928_),
    .X(_17929_));
 sky130_fd_sc_hd__and3_1 _46815_ (.A(_13097_),
    .B(_17927_),
    .C(_17929_),
    .X(_17930_));
 sky130_fd_sc_hd__nand2_1 _46816_ (.A(_17927_),
    .B(_17928_),
    .Y(_17931_));
 sky130_fd_sc_hd__and3_1 _46817_ (.A(_17931_),
    .B(_13075_),
    .C(_13020_),
    .X(_17932_));
 sky130_fd_sc_hd__o21ai_1 _46818_ (.A1(_12339_),
    .A2(_12361_),
    .B1(_12416_),
    .Y(_17933_));
 sky130_fd_sc_hd__clkbuf_2 _46819_ (.A(\delay_line[4][2] ),
    .X(_17934_));
 sky130_fd_sc_hd__nor2_1 _46820_ (.A(\delay_line[4][0] ),
    .B(_17934_),
    .Y(_17935_));
 sky130_fd_sc_hd__and2_1 _46821_ (.A(\delay_line[4][0] ),
    .B(_17934_),
    .X(_17936_));
 sky130_fd_sc_hd__clkbuf_2 _46822_ (.A(\delay_line[11][3] ),
    .X(_17937_));
 sky130_fd_sc_hd__o21bai_1 _46823_ (.A1(_17935_),
    .A2(_17936_),
    .B1_N(_17937_),
    .Y(_17938_));
 sky130_fd_sc_hd__clkbuf_2 _46824_ (.A(_17938_),
    .X(_17939_));
 sky130_fd_sc_hd__inv_2 _46825_ (.A(\delay_line[4][2] ),
    .Y(_17940_));
 sky130_fd_sc_hd__clkbuf_2 _46826_ (.A(_17940_),
    .X(_17941_));
 sky130_fd_sc_hd__o21a_1 _46827_ (.A1(_07975_),
    .A2(_17934_),
    .B1(_17937_),
    .X(_17942_));
 sky130_fd_sc_hd__o21ai_1 _46828_ (.A1(_08140_),
    .A2(_17941_),
    .B1(_17942_),
    .Y(_17943_));
 sky130_fd_sc_hd__buf_1 _46829_ (.A(\delay_line[0][5] ),
    .X(_17944_));
 sky130_fd_sc_hd__a21o_1 _46830_ (.A1(_17939_),
    .A2(_17943_),
    .B1(_17944_),
    .X(_17945_));
 sky130_fd_sc_hd__clkbuf_2 _46831_ (.A(_17934_),
    .X(_17946_));
 sky130_fd_sc_hd__o21ai_2 _46832_ (.A1(_08052_),
    .A2(_17946_),
    .B1(_17937_),
    .Y(_17947_));
 sky130_fd_sc_hd__o211ai_2 _46833_ (.A1(_17936_),
    .A2(_17947_),
    .B1(_17944_),
    .C1(_17939_),
    .Y(_17948_));
 sky130_fd_sc_hd__and3_2 _46834_ (.A(_17933_),
    .B(_17945_),
    .C(_17948_),
    .X(_17949_));
 sky130_fd_sc_hd__clkbuf_2 _46835_ (.A(\delay_line[0][5] ),
    .X(_17950_));
 sky130_fd_sc_hd__a21oi_1 _46836_ (.A1(_17939_),
    .A2(_17943_),
    .B1(_17950_),
    .Y(_17951_));
 sky130_fd_sc_hd__o211a_1 _46837_ (.A1(_17936_),
    .A2(_17947_),
    .B1(\delay_line[0][5] ),
    .C1(_17939_),
    .X(_17952_));
 sky130_fd_sc_hd__o21a_1 _46838_ (.A1(_12339_),
    .A2(_12361_),
    .B1(_12416_),
    .X(_17953_));
 sky130_fd_sc_hd__o21ai_2 _46839_ (.A1(_17951_),
    .A2(_17952_),
    .B1(_17953_),
    .Y(_17954_));
 sky130_fd_sc_hd__buf_1 _46840_ (.A(_12383_),
    .X(_17955_));
 sky130_fd_sc_hd__clkbuf_2 _46841_ (.A(_17955_),
    .X(_17956_));
 sky130_fd_sc_hd__nand2_1 _46842_ (.A(_17954_),
    .B(_17956_),
    .Y(_17957_));
 sky130_fd_sc_hd__inv_2 _46843_ (.A(_12449_),
    .Y(_17958_));
 sky130_fd_sc_hd__a21oi_2 _46844_ (.A1(_08085_),
    .A2(_12559_),
    .B1(_17958_),
    .Y(_17959_));
 sky130_fd_sc_hd__nand3_1 _46845_ (.A(_17933_),
    .B(_17945_),
    .C(_17948_),
    .Y(_17960_));
 sky130_fd_sc_hd__a21o_1 _46846_ (.A1(_17954_),
    .A2(_17960_),
    .B1(_17955_),
    .X(_17961_));
 sky130_fd_sc_hd__o211a_2 _46847_ (.A1(_17949_),
    .A2(_17957_),
    .B1(_17959_),
    .C1(_17961_),
    .X(_17962_));
 sky130_fd_sc_hd__o21a_1 _46848_ (.A1(_12328_),
    .A2(_12394_),
    .B1(_08085_),
    .X(_17963_));
 sky130_fd_sc_hd__a21oi_1 _46849_ (.A1(_17954_),
    .A2(_17960_),
    .B1(_17956_),
    .Y(_17964_));
 sky130_fd_sc_hd__and3_1 _46850_ (.A(_17954_),
    .B(_17960_),
    .C(_17955_),
    .X(_17965_));
 sky130_fd_sc_hd__o22ai_4 _46851_ (.A1(_17958_),
    .A2(_17963_),
    .B1(_17964_),
    .B2(_17965_),
    .Y(_17966_));
 sky130_fd_sc_hd__xor2_2 _46852_ (.A(\delay_line[0][1] ),
    .B(net397),
    .X(_17967_));
 sky130_fd_sc_hd__and3_2 _46853_ (.A(_23161_),
    .B(_12207_),
    .C(_17967_),
    .X(_17968_));
 sky130_fd_sc_hd__a21oi_2 _46854_ (.A1(_23161_),
    .A2(_12207_),
    .B1(_17967_),
    .Y(_17969_));
 sky130_fd_sc_hd__nor2_1 _46855_ (.A(_17968_),
    .B(_17969_),
    .Y(_17970_));
 sky130_fd_sc_hd__nand2_1 _46856_ (.A(_17966_),
    .B(_17970_),
    .Y(_17971_));
 sky130_fd_sc_hd__o211ai_4 _46857_ (.A1(_17949_),
    .A2(_17957_),
    .B1(_17959_),
    .C1(_17961_),
    .Y(_17972_));
 sky130_fd_sc_hd__o2bb2ai_4 _46858_ (.A1_N(_17972_),
    .A2_N(_17966_),
    .B1(_17968_),
    .B2(_17969_),
    .Y(_17973_));
 sky130_fd_sc_hd__o221a_1 _46859_ (.A1(_12603_),
    .A2(_12724_),
    .B1(_17962_),
    .B2(_17971_),
    .C1(_17973_),
    .X(_17974_));
 sky130_fd_sc_hd__nand3_1 _46860_ (.A(_17972_),
    .B(_17966_),
    .C(_17970_),
    .Y(_17975_));
 sky130_fd_sc_hd__o31a_1 _46861_ (.A1(_12218_),
    .A2(_12229_),
    .A3(_12515_),
    .B1(_12636_),
    .X(_17976_));
 sky130_fd_sc_hd__a21boi_2 _46862_ (.A1(_17973_),
    .A2(_17975_),
    .B1_N(_17976_),
    .Y(_17977_));
 sky130_fd_sc_hd__clkbuf_2 _46863_ (.A(_08272_),
    .X(_17978_));
 sky130_fd_sc_hd__clkbuf_2 _46864_ (.A(_17978_),
    .X(_17979_));
 sky130_fd_sc_hd__o21ai_1 _46865_ (.A1(_17974_),
    .A2(_17977_),
    .B1(_17979_),
    .Y(_17980_));
 sky130_fd_sc_hd__inv_2 _46866_ (.A(_17978_),
    .Y(_17981_));
 sky130_fd_sc_hd__buf_2 _46867_ (.A(_17981_),
    .X(_17982_));
 sky130_fd_sc_hd__o221ai_4 _46868_ (.A1(_12603_),
    .A2(_12724_),
    .B1(_17962_),
    .B2(_17971_),
    .C1(_17973_),
    .Y(_17983_));
 sky130_fd_sc_hd__a21bo_1 _46869_ (.A1(_17973_),
    .A2(_17975_),
    .B1_N(_17976_),
    .X(_17984_));
 sky130_fd_sc_hd__nand3_1 _46870_ (.A(_17982_),
    .B(_17983_),
    .C(_17984_),
    .Y(_17985_));
 sky130_fd_sc_hd__o31a_1 _46871_ (.A1(_12691_),
    .A2(_12702_),
    .A3(_12724_),
    .B1(_12834_),
    .X(_17986_));
 sky130_fd_sc_hd__nand3_1 _46872_ (.A(_17980_),
    .B(_17985_),
    .C(_17986_),
    .Y(_17987_));
 sky130_fd_sc_hd__inv_2 _46873_ (.A(_12834_),
    .Y(_17988_));
 sky130_fd_sc_hd__nand3_1 _46874_ (.A(_17984_),
    .B(_17979_),
    .C(_17983_),
    .Y(_17989_));
 sky130_fd_sc_hd__o21ai_1 _46875_ (.A1(_17974_),
    .A2(_17977_),
    .B1(_17981_),
    .Y(_17990_));
 sky130_fd_sc_hd__o211ai_2 _46876_ (.A1(_12735_),
    .A2(_17988_),
    .B1(_17989_),
    .C1(_17990_),
    .Y(_17991_));
 sky130_fd_sc_hd__nand2_2 _46877_ (.A(_12130_),
    .B(net407),
    .Y(_17992_));
 sky130_fd_sc_hd__nor2_1 _46878_ (.A(\delay_line[12][4] ),
    .B(net406),
    .Y(_17993_));
 sky130_fd_sc_hd__nand2_1 _46879_ (.A(\delay_line[12][4] ),
    .B(net406),
    .Y(_17994_));
 sky130_fd_sc_hd__buf_2 _46880_ (.A(_17994_),
    .X(_17995_));
 sky130_fd_sc_hd__or2b_1 _46881_ (.A(_17993_),
    .B_N(_17995_),
    .X(_17996_));
 sky130_fd_sc_hd__nor2_2 _46882_ (.A(net406),
    .B(_17992_),
    .Y(_17997_));
 sky130_fd_sc_hd__a211oi_2 _46883_ (.A1(_17992_),
    .A2(_17996_),
    .B1(_17997_),
    .C1(_23260_),
    .Y(_17998_));
 sky130_fd_sc_hd__a21oi_2 _46884_ (.A1(_17992_),
    .A2(_17996_),
    .B1(_17997_),
    .Y(_17999_));
 sky130_fd_sc_hd__and2b_1 _46885_ (.A_N(_17999_),
    .B(_23260_),
    .X(_18000_));
 sky130_fd_sc_hd__o2bb2ai_2 _46886_ (.A1_N(_17987_),
    .A2_N(_17991_),
    .B1(_17998_),
    .B2(_18000_),
    .Y(_18001_));
 sky130_fd_sc_hd__o21a_2 _46887_ (.A1(_12867_),
    .A2(_12823_),
    .B1(_12888_),
    .X(_18002_));
 sky130_fd_sc_hd__and2_2 _46888_ (.A(_23227_),
    .B(_17999_),
    .X(_18003_));
 sky130_fd_sc_hd__nor2_2 _46889_ (.A(_23260_),
    .B(_17999_),
    .Y(_18004_));
 sky130_fd_sc_hd__clkbuf_2 _46890_ (.A(_17987_),
    .X(_18005_));
 sky130_fd_sc_hd__clkbuf_2 _46891_ (.A(_17991_),
    .X(_18006_));
 sky130_fd_sc_hd__o211ai_4 _46892_ (.A1(_18003_),
    .A2(_18004_),
    .B1(_18005_),
    .C1(_18006_),
    .Y(_18007_));
 sky130_fd_sc_hd__nand3_4 _46893_ (.A(_18001_),
    .B(_18002_),
    .C(_18007_),
    .Y(_18008_));
 sky130_fd_sc_hd__o21ai_2 _46894_ (.A1(_17930_),
    .A2(_17932_),
    .B1(_18008_),
    .Y(_18009_));
 sky130_fd_sc_hd__inv_2 _46895_ (.A(_18002_),
    .Y(_18010_));
 sky130_fd_sc_hd__o2bb2ai_2 _46896_ (.A1_N(_18005_),
    .A2_N(_18006_),
    .B1(_18003_),
    .B2(_18004_),
    .Y(_18011_));
 sky130_fd_sc_hd__o211ai_2 _46897_ (.A1(_17998_),
    .A2(_18000_),
    .B1(_18005_),
    .C1(_18006_),
    .Y(_18012_));
 sky130_fd_sc_hd__and3_2 _46898_ (.A(_18010_),
    .B(_18011_),
    .C(_18012_),
    .X(_18013_));
 sky130_fd_sc_hd__a32o_1 _46899_ (.A1(_12119_),
    .A2(_12856_),
    .A3(_12899_),
    .B1(_12954_),
    .B2(_13174_),
    .X(_18014_));
 sky130_fd_sc_hd__nand3_2 _46900_ (.A(_18010_),
    .B(_18011_),
    .C(_18012_),
    .Y(_18015_));
 sky130_fd_sc_hd__and4_1 _46901_ (.A(_17928_),
    .B(_13075_),
    .C(_13020_),
    .D(_17927_),
    .X(_18016_));
 sky130_fd_sc_hd__o41a_2 _46902_ (.A1(_12998_),
    .A2(_13009_),
    .A3(_13053_),
    .A4(_13064_),
    .B1(_17931_),
    .X(_18017_));
 sky130_fd_sc_hd__o2bb2ai_2 _46903_ (.A1_N(_18015_),
    .A2_N(_18008_),
    .B1(_18016_),
    .B2(_18017_),
    .Y(_18018_));
 sky130_fd_sc_hd__o211ai_4 _46904_ (.A1(_18009_),
    .A2(_18013_),
    .B1(_18014_),
    .C1(_18018_),
    .Y(_18019_));
 sky130_fd_sc_hd__o2bb2ai_1 _46905_ (.A1_N(_18015_),
    .A2_N(_18008_),
    .B1(_17930_),
    .B2(_17932_),
    .Y(_18020_));
 sky130_fd_sc_hd__a21oi_1 _46906_ (.A1(_13174_),
    .A2(_12954_),
    .B1(_13273_),
    .Y(_18021_));
 sky130_fd_sc_hd__o211ai_2 _46907_ (.A1(_18016_),
    .A2(_18017_),
    .B1(_18015_),
    .C1(_18008_),
    .Y(_18022_));
 sky130_fd_sc_hd__nand3_1 _46908_ (.A(_18020_),
    .B(_18021_),
    .C(_18022_),
    .Y(_18023_));
 sky130_fd_sc_hd__clkbuf_2 _46909_ (.A(_18023_),
    .X(_18024_));
 sky130_fd_sc_hd__clkbuf_2 _46910_ (.A(\delay_line[7][5] ),
    .X(_18025_));
 sky130_fd_sc_hd__clkbuf_4 _46911_ (.A(_18025_),
    .X(_18026_));
 sky130_fd_sc_hd__xnor2_2 _46912_ (.A(_18026_),
    .B(_11800_),
    .Y(_18027_));
 sky130_fd_sc_hd__o21a_1 _46913_ (.A1(_03172_),
    .A2(_08921_),
    .B1(\delay_line[8][1] ),
    .X(_18028_));
 sky130_fd_sc_hd__nor2_1 _46914_ (.A(\delay_line[8][3] ),
    .B(\delay_line[8][4] ),
    .Y(_18029_));
 sky130_fd_sc_hd__buf_1 _46915_ (.A(\delay_line[8][4] ),
    .X(_18030_));
 sky130_fd_sc_hd__nand2_1 _46916_ (.A(\delay_line[8][3] ),
    .B(_18030_),
    .Y(_18031_));
 sky130_fd_sc_hd__nand3b_1 _46917_ (.A_N(_18029_),
    .B(_18031_),
    .C(\delay_line[8][2] ),
    .Y(_18032_));
 sky130_fd_sc_hd__buf_1 _46918_ (.A(_18032_),
    .X(_18033_));
 sky130_fd_sc_hd__and2_1 _46919_ (.A(_08921_),
    .B(_18030_),
    .X(_18034_));
 sky130_fd_sc_hd__o21bai_1 _46920_ (.A1(_18029_),
    .A2(_18034_),
    .B1_N(_03172_),
    .Y(_18035_));
 sky130_fd_sc_hd__o211a_2 _46921_ (.A1(_11767_),
    .A2(_18028_),
    .B1(_18033_),
    .C1(_18035_),
    .X(_18036_));
 sky130_fd_sc_hd__a21o_1 _46922_ (.A1(_03205_),
    .A2(_08932_),
    .B1(_18028_),
    .X(_18037_));
 sky130_fd_sc_hd__a21o_1 _46923_ (.A1(_18033_),
    .A2(_18035_),
    .B1(_18037_),
    .X(_18038_));
 sky130_fd_sc_hd__buf_1 _46924_ (.A(\delay_line[8][5] ),
    .X(_18039_));
 sky130_fd_sc_hd__buf_2 _46925_ (.A(_18039_),
    .X(_18040_));
 sky130_fd_sc_hd__nand3b_1 _46926_ (.A_N(_18036_),
    .B(_18038_),
    .C(_18040_),
    .Y(_18041_));
 sky130_fd_sc_hd__buf_1 _46927_ (.A(_18041_),
    .X(_18042_));
 sky130_fd_sc_hd__a21oi_1 _46928_ (.A1(_18033_),
    .A2(_18035_),
    .B1(_18037_),
    .Y(_18043_));
 sky130_fd_sc_hd__buf_2 _46929_ (.A(_18040_),
    .X(_18044_));
 sky130_fd_sc_hd__o21bai_2 _46930_ (.A1(_18036_),
    .A2(_18043_),
    .B1_N(_18044_),
    .Y(_18045_));
 sky130_fd_sc_hd__and3_1 _46931_ (.A(_11855_),
    .B(_18042_),
    .C(_18045_),
    .X(_18046_));
 sky130_fd_sc_hd__a21oi_1 _46932_ (.A1(_18042_),
    .A2(_18045_),
    .B1(_11855_),
    .Y(_18047_));
 sky130_fd_sc_hd__nor2_1 _46933_ (.A(_18046_),
    .B(_18047_),
    .Y(_18048_));
 sky130_fd_sc_hd__xnor2_2 _46934_ (.A(_18027_),
    .B(_18048_),
    .Y(_18049_));
 sky130_fd_sc_hd__or2b_1 _46935_ (.A(_02876_),
    .B_N(_02854_),
    .X(_18050_));
 sky130_fd_sc_hd__and4_1 _46936_ (.A(_11691_),
    .B(_02876_),
    .C(_08668_),
    .D(_23084_),
    .X(_18051_));
 sky130_fd_sc_hd__buf_2 _46937_ (.A(_12987_),
    .X(_18052_));
 sky130_fd_sc_hd__clkbuf_2 _46938_ (.A(net422),
    .X(_18053_));
 sky130_fd_sc_hd__and2b_2 _46939_ (.A_N(\delay_line[9][2] ),
    .B(\delay_line[9][4] ),
    .X(_18054_));
 sky130_fd_sc_hd__or2b_1 _46940_ (.A(\delay_line[9][4] ),
    .B_N(\delay_line[9][2] ),
    .X(_18055_));
 sky130_fd_sc_hd__and2b_1 _46941_ (.A_N(_18054_),
    .B(_18055_),
    .X(_18056_));
 sky130_fd_sc_hd__o21a_1 _46942_ (.A1(_18053_),
    .A2(_08899_),
    .B1(_18056_),
    .X(_18057_));
 sky130_fd_sc_hd__buf_2 _46943_ (.A(_18056_),
    .X(_18058_));
 sky130_fd_sc_hd__nor3_1 _46944_ (.A(_18053_),
    .B(_08899_),
    .C(_18058_),
    .Y(_18059_));
 sky130_fd_sc_hd__a211oi_1 _46945_ (.A1(_25051_),
    .A2(_18052_),
    .B1(_18057_),
    .C1(_18059_),
    .Y(_18060_));
 sky130_fd_sc_hd__o211a_1 _46946_ (.A1(_18057_),
    .A2(_18059_),
    .B1(_25051_),
    .C1(_18052_),
    .X(_18061_));
 sky130_fd_sc_hd__nor2_1 _46947_ (.A(_18060_),
    .B(_18061_),
    .Y(_18062_));
 sky130_fd_sc_hd__a311o_1 _46948_ (.A1(_23117_),
    .A2(_11669_),
    .A3(_18050_),
    .B1(_18051_),
    .C1(_18062_),
    .X(_18063_));
 sky130_fd_sc_hd__a31o_1 _46949_ (.A1(_23106_),
    .A2(_11669_),
    .A3(_18050_),
    .B1(_18051_),
    .X(_18064_));
 sky130_fd_sc_hd__nand2_1 _46950_ (.A(_18062_),
    .B(_18064_),
    .Y(_18065_));
 sky130_fd_sc_hd__and2_1 _46951_ (.A(_18063_),
    .B(_18065_),
    .X(_18066_));
 sky130_fd_sc_hd__nand2_1 _46952_ (.A(_18049_),
    .B(_18066_),
    .Y(_18067_));
 sky130_fd_sc_hd__a31o_1 _46953_ (.A1(_13086_),
    .A2(_13097_),
    .A3(_13108_),
    .B1(_13152_),
    .X(_18068_));
 sky130_fd_sc_hd__o21a_1 _46954_ (.A1(_18049_),
    .A2(_18066_),
    .B1(_18068_),
    .X(_18069_));
 sky130_fd_sc_hd__or2_1 _46955_ (.A(_18049_),
    .B(_18066_),
    .X(_18070_));
 sky130_fd_sc_hd__a21oi_1 _46956_ (.A1(_18067_),
    .A2(_18070_),
    .B1(_18068_),
    .Y(_18071_));
 sky130_fd_sc_hd__a21o_1 _46957_ (.A1(_18067_),
    .A2(_18069_),
    .B1(_18071_),
    .X(_18072_));
 sky130_fd_sc_hd__xnor2_2 _46958_ (.A(_12064_),
    .B(_18072_),
    .Y(_18073_));
 sky130_fd_sc_hd__a21oi_1 _46959_ (.A1(_18019_),
    .A2(_18024_),
    .B1(_18073_),
    .Y(_18074_));
 sky130_fd_sc_hd__nand3_1 _46960_ (.A(_18019_),
    .B(_18024_),
    .C(_18073_),
    .Y(_18075_));
 sky130_fd_sc_hd__a21oi_1 _46961_ (.A1(_12108_),
    .A2(_13240_),
    .B1(_13306_),
    .Y(_18076_));
 sky130_fd_sc_hd__nand2_1 _46962_ (.A(_18075_),
    .B(_18076_),
    .Y(_18077_));
 sky130_fd_sc_hd__nor2_1 _46963_ (.A(_22963_),
    .B(_00062_),
    .Y(_18078_));
 sky130_fd_sc_hd__nor2_1 _46964_ (.A(_23018_),
    .B(_03447_),
    .Y(_18079_));
 sky130_fd_sc_hd__clkbuf_2 _46965_ (.A(net429),
    .X(_18080_));
 sky130_fd_sc_hd__or3b_2 _46966_ (.A(_18078_),
    .B(_18079_),
    .C_N(_18080_),
    .X(_18081_));
 sky130_fd_sc_hd__buf_2 _46967_ (.A(_18080_),
    .X(_18082_));
 sky130_fd_sc_hd__o21bai_1 _46968_ (.A1(_18078_),
    .A2(_18079_),
    .B1_N(_18082_),
    .Y(_18083_));
 sky130_fd_sc_hd__nand3b_1 _46969_ (.A_N(_11998_),
    .B(_18081_),
    .C(_18083_),
    .Y(_18084_));
 sky130_fd_sc_hd__a32o_1 _46970_ (.A1(_11899_),
    .A2(_11976_),
    .A3(_00095_),
    .B1(_18081_),
    .B2(_18083_),
    .X(_18085_));
 sky130_fd_sc_hd__nand2_1 _46971_ (.A(_18084_),
    .B(_18085_),
    .Y(_18086_));
 sky130_fd_sc_hd__xnor2_1 _46972_ (.A(_13482_),
    .B(_18086_),
    .Y(_18087_));
 sky130_fd_sc_hd__a21o_1 _46973_ (.A1(_11921_),
    .A2(_12031_),
    .B1(_18087_),
    .X(_18088_));
 sky130_fd_sc_hd__nand3_1 _46974_ (.A(_11921_),
    .B(_12031_),
    .C(_18087_),
    .Y(_18089_));
 sky130_fd_sc_hd__nand3b_1 _46975_ (.A_N(_13504_),
    .B(_18088_),
    .C(_18089_),
    .Y(_18090_));
 sky130_fd_sc_hd__a32o_1 _46976_ (.A1(_13471_),
    .A2(_13482_),
    .A3(_13493_),
    .B1(_18088_),
    .B2(_18089_),
    .X(_18091_));
 sky130_fd_sc_hd__nor2_1 _46977_ (.A(_24809_),
    .B(_03414_),
    .Y(_18092_));
 sky130_fd_sc_hd__o21a_1 _46978_ (.A1(_22908_),
    .A2(_18092_),
    .B1(_09228_),
    .X(_18093_));
 sky130_fd_sc_hd__buf_1 _46979_ (.A(\delay_line[6][3] ),
    .X(_18094_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46980_ (.A(_18094_),
    .X(_18095_));
 sky130_fd_sc_hd__inv_2 _46981_ (.A(\delay_line[6][0] ),
    .Y(_18096_));
 sky130_fd_sc_hd__o211a_1 _46982_ (.A1(_24809_),
    .A2(_03414_),
    .B1(_18095_),
    .C1(_18096_),
    .X(_18097_));
 sky130_fd_sc_hd__clkbuf_2 _46983_ (.A(_09481_),
    .X(_18098_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46984_ (.A(\delay_line[3][5] ),
    .X(_18099_));
 sky130_fd_sc_hd__nor2_1 _46985_ (.A(_18098_),
    .B(_18099_),
    .Y(_18100_));
 sky130_fd_sc_hd__clkbuf_2 _46986_ (.A(_09481_),
    .X(_18101_));
 sky130_fd_sc_hd__and2_1 _46987_ (.A(_18101_),
    .B(_18099_),
    .X(_18102_));
 sky130_fd_sc_hd__clkbuf_2 _46988_ (.A(_13559_),
    .X(_18103_));
 sky130_fd_sc_hd__buf_2 _46989_ (.A(\delay_line[5][5] ),
    .X(_18104_));
 sky130_fd_sc_hd__nor2_1 _46990_ (.A(_18103_),
    .B(_18104_),
    .Y(_18105_));
 sky130_fd_sc_hd__and2_1 _46991_ (.A(_13559_),
    .B(\delay_line[5][5] ),
    .X(_18106_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _46992_ (.A(_18106_),
    .X(_18107_));
 sky130_fd_sc_hd__o21a_1 _46993_ (.A1(_03535_),
    .A2(_18103_),
    .B1(_09481_),
    .X(_18108_));
 sky130_fd_sc_hd__o21ai_1 _46994_ (.A1(_18105_),
    .A2(_18107_),
    .B1(_18108_),
    .Y(_18109_));
 sky130_fd_sc_hd__or3_1 _46995_ (.A(_18105_),
    .B(_18106_),
    .C(_18108_),
    .X(_18110_));
 sky130_fd_sc_hd__o211a_1 _46996_ (.A1(_18100_),
    .A2(_18102_),
    .B1(_18109_),
    .C1(_18110_),
    .X(_18111_));
 sky130_fd_sc_hd__a211oi_1 _46997_ (.A1(_18109_),
    .A2(_18110_),
    .B1(_18100_),
    .C1(_18102_),
    .Y(_18112_));
 sky130_fd_sc_hd__nor4_1 _46998_ (.A(_18093_),
    .B(_18097_),
    .C(_18111_),
    .D(_18112_),
    .Y(_18113_));
 sky130_fd_sc_hd__o22a_1 _46999_ (.A1(_18093_),
    .A2(_18097_),
    .B1(_18111_),
    .B2(_18112_),
    .X(_18114_));
 sky130_fd_sc_hd__nor3_1 _47000_ (.A(_13735_),
    .B(net212),
    .C(_18114_),
    .Y(_18115_));
 sky130_fd_sc_hd__o32a_1 _47001_ (.A1(_13647_),
    .A2(_13702_),
    .A3(_13658_),
    .B1(_18114_),
    .B2(net212),
    .X(_18116_));
 sky130_fd_sc_hd__nor2_1 _47002_ (.A(_18115_),
    .B(_18116_),
    .Y(_18117_));
 sky130_fd_sc_hd__and3_1 _47003_ (.A(_03590_),
    .B(_03546_),
    .C(_13570_),
    .X(_18118_));
 sky130_fd_sc_hd__and2b_1 _47004_ (.A_N(net443),
    .B(net436),
    .X(_18119_));
 sky130_fd_sc_hd__nor2_1 _47005_ (.A(_03502_),
    .B(_13779_),
    .Y(_18120_));
 sky130_fd_sc_hd__nand2_1 _47006_ (.A(_13834_),
    .B(net443),
    .Y(_18121_));
 sky130_fd_sc_hd__nand3b_2 _47007_ (.A_N(_18119_),
    .B(_18120_),
    .C(_18121_),
    .Y(_18122_));
 sky130_fd_sc_hd__and2b_1 _47008_ (.A_N(net436),
    .B(\delay_line[2][5] ),
    .X(_18123_));
 sky130_fd_sc_hd__o22ai_2 _47009_ (.A1(_03502_),
    .A2(_13779_),
    .B1(_18123_),
    .B2(_18119_),
    .Y(_18124_));
 sky130_fd_sc_hd__nand4_1 _47010_ (.A(_18122_),
    .B(_18124_),
    .C(_03546_),
    .D(_13592_),
    .Y(_18125_));
 sky130_fd_sc_hd__a22o_1 _47011_ (.A1(_03535_),
    .A2(_13592_),
    .B1(_18122_),
    .B2(_18124_),
    .X(_18126_));
 sky130_fd_sc_hd__nand3b_1 _47012_ (.A_N(_13812_),
    .B(_18125_),
    .C(_18126_),
    .Y(_18127_));
 sky130_fd_sc_hd__a21bo_1 _47013_ (.A1(_18125_),
    .A2(_18126_),
    .B1_N(_13812_),
    .X(_18128_));
 sky130_fd_sc_hd__o211a_1 _47014_ (.A1(_13647_),
    .A2(_18118_),
    .B1(_18127_),
    .C1(_18128_),
    .X(_18129_));
 sky130_fd_sc_hd__a31o_1 _47015_ (.A1(_13581_),
    .A2(_13603_),
    .A3(_13636_),
    .B1(_18118_),
    .X(_18130_));
 sky130_fd_sc_hd__a21oi_1 _47016_ (.A1(_18127_),
    .A2(_18128_),
    .B1(_18130_),
    .Y(_18131_));
 sky130_fd_sc_hd__and2_1 _47017_ (.A(_13823_),
    .B(_13878_),
    .X(_18132_));
 sky130_fd_sc_hd__o21ai_1 _47018_ (.A1(_18129_),
    .A2(_18131_),
    .B1(_18132_),
    .Y(_18133_));
 sky130_fd_sc_hd__or3_1 _47019_ (.A(_18132_),
    .B(_18129_),
    .C(_18131_),
    .X(_18134_));
 sky130_fd_sc_hd__nand2_1 _47020_ (.A(_18133_),
    .B(_18134_),
    .Y(_18135_));
 sky130_fd_sc_hd__xnor2_2 _47021_ (.A(_18117_),
    .B(_18135_),
    .Y(_18136_));
 sky130_fd_sc_hd__a21o_1 _47022_ (.A1(_18090_),
    .A2(_18091_),
    .B1(_18136_),
    .X(_18137_));
 sky130_fd_sc_hd__nand3_1 _47023_ (.A(_18136_),
    .B(_18090_),
    .C(_18091_),
    .Y(_18138_));
 sky130_fd_sc_hd__o21bai_1 _47024_ (.A1(_09064_),
    .A2(_12075_),
    .B1_N(_12086_),
    .Y(_18139_));
 sky130_fd_sc_hd__a21oi_1 _47025_ (.A1(_18137_),
    .A2(_18138_),
    .B1(_18139_),
    .Y(_18140_));
 sky130_fd_sc_hd__nand3_1 _47026_ (.A(_18139_),
    .B(_18137_),
    .C(_18138_),
    .Y(_18141_));
 sky130_fd_sc_hd__and2b_1 _47027_ (.A_N(_18140_),
    .B(_18141_),
    .X(_18142_));
 sky130_fd_sc_hd__a31o_1 _47028_ (.A1(_09239_),
    .A2(_13515_),
    .A3(_13504_),
    .B1(_14031_),
    .X(_18143_));
 sky130_fd_sc_hd__inv_2 _47029_ (.A(_18143_),
    .Y(_18144_));
 sky130_fd_sc_hd__xnor2_2 _47030_ (.A(_18142_),
    .B(_18144_),
    .Y(_18145_));
 sky130_fd_sc_hd__o21a_1 _47031_ (.A1(_18074_),
    .A2(_18077_),
    .B1(_18145_),
    .X(_18146_));
 sky130_fd_sc_hd__nand2_1 _47032_ (.A(_18069_),
    .B(_18067_),
    .Y(_18147_));
 sky130_fd_sc_hd__nor2_1 _47033_ (.A(_12064_),
    .B(_18071_),
    .Y(_18148_));
 sky130_fd_sc_hd__and3_1 _47034_ (.A(_18068_),
    .B(_18067_),
    .C(_18070_),
    .X(_18149_));
 sky130_fd_sc_hd__o21a_1 _47035_ (.A1(_18149_),
    .A2(_18071_),
    .B1(_12064_),
    .X(_18150_));
 sky130_fd_sc_hd__a21oi_1 _47036_ (.A1(_18147_),
    .A2(_18148_),
    .B1(_18150_),
    .Y(_18151_));
 sky130_fd_sc_hd__nand2_1 _47037_ (.A(_18024_),
    .B(_18151_),
    .Y(_18152_));
 sky130_fd_sc_hd__o211a_2 _47038_ (.A1(_18009_),
    .A2(_18013_),
    .B1(_18014_),
    .C1(_18018_),
    .X(_18153_));
 sky130_fd_sc_hd__a21o_1 _47039_ (.A1(_12108_),
    .A2(_13240_),
    .B1(_13306_),
    .X(_18154_));
 sky130_fd_sc_hd__nor2_1 _47040_ (.A(_12064_),
    .B(_18072_),
    .Y(_18155_));
 sky130_fd_sc_hd__o2bb2ai_1 _47041_ (.A1_N(_18019_),
    .A2_N(_18023_),
    .B1(_18150_),
    .B2(_18155_),
    .Y(_18156_));
 sky130_fd_sc_hd__o211ai_2 _47042_ (.A1(_18152_),
    .A2(_18153_),
    .B1(_18154_),
    .C1(_18156_),
    .Y(_18157_));
 sky130_fd_sc_hd__nand2_1 _47043_ (.A(_18146_),
    .B(_18157_),
    .Y(_18158_));
 sky130_fd_sc_hd__a21o_1 _47044_ (.A1(_18019_),
    .A2(_18024_),
    .B1(_18073_),
    .X(_18159_));
 sky130_fd_sc_hd__nand3_1 _47045_ (.A(_18159_),
    .B(_18076_),
    .C(_18075_),
    .Y(_18160_));
 sky130_fd_sc_hd__a21o_1 _47046_ (.A1(_18157_),
    .A2(_18160_),
    .B1(_18145_),
    .X(_18161_));
 sky130_fd_sc_hd__nand3_4 _47047_ (.A(_17908_),
    .B(_18158_),
    .C(_18161_),
    .Y(_18162_));
 sky130_fd_sc_hd__clkbuf_2 _47048_ (.A(_18162_),
    .X(_18163_));
 sky130_fd_sc_hd__o211a_1 _47049_ (.A1(_18074_),
    .A2(_18077_),
    .B1(_18145_),
    .C1(_18157_),
    .X(_18164_));
 sky130_fd_sc_hd__a21oi_1 _47050_ (.A1(_18157_),
    .A2(_18160_),
    .B1(_18145_),
    .Y(_18165_));
 sky130_fd_sc_hd__o21bai_4 _47051_ (.A1(_18164_),
    .A2(_18165_),
    .B1_N(_17908_),
    .Y(_18166_));
 sky130_fd_sc_hd__clkbuf_2 _47052_ (.A(_18166_),
    .X(_18167_));
 sky130_fd_sc_hd__a32oi_2 _47053_ (.A1(_09514_),
    .A2(_13878_),
    .A3(_13867_),
    .B1(_13911_),
    .B2(_13932_),
    .Y(_18168_));
 sky130_fd_sc_hd__nor2_1 _47054_ (.A(net451),
    .B(\delay_line[1][5] ),
    .Y(_18169_));
 sky130_fd_sc_hd__nand2_2 _47055_ (.A(net451),
    .B(\delay_line[1][5] ),
    .Y(_18170_));
 sky130_fd_sc_hd__nand3b_2 _47056_ (.A_N(_18169_),
    .B(_18170_),
    .C(\delay_line[2][2] ),
    .Y(_18171_));
 sky130_fd_sc_hd__clkbuf_2 _47057_ (.A(_18169_),
    .X(_18172_));
 sky130_fd_sc_hd__and2_1 _47058_ (.A(net451),
    .B(\delay_line[1][5] ),
    .X(_18173_));
 sky130_fd_sc_hd__clkbuf_2 _47059_ (.A(_18173_),
    .X(_18174_));
 sky130_fd_sc_hd__o21ai_2 _47060_ (.A1(_18172_),
    .A2(_18174_),
    .B1(_03678_),
    .Y(_18175_));
 sky130_fd_sc_hd__o2111ai_2 _47061_ (.A1(_14328_),
    .A2(_14339_),
    .B1(_24930_),
    .C1(_18171_),
    .D1(_18175_),
    .Y(_18176_));
 sky130_fd_sc_hd__nor2_1 _47062_ (.A(_14328_),
    .B(_14339_),
    .Y(_18177_));
 sky130_fd_sc_hd__o2bb2ai_1 _47063_ (.A1_N(_18171_),
    .A2_N(_18175_),
    .B1(_14361_),
    .B2(_18177_),
    .Y(_18178_));
 sky130_fd_sc_hd__nand2_1 _47064_ (.A(_18176_),
    .B(_18178_),
    .Y(_18179_));
 sky130_fd_sc_hd__and2b_1 _47065_ (.A_N(\delay_line[1][1] ),
    .B(_09745_),
    .X(_18180_));
 sky130_fd_sc_hd__xnor2_1 _47066_ (.A(_14328_),
    .B(_18180_),
    .Y(_18181_));
 sky130_fd_sc_hd__nand2_1 _47067_ (.A(_18179_),
    .B(_18181_),
    .Y(_18182_));
 sky130_fd_sc_hd__nand3b_1 _47068_ (.A_N(_18181_),
    .B(_18176_),
    .C(_18178_),
    .Y(_18183_));
 sky130_fd_sc_hd__o21ai_1 _47069_ (.A1(_14405_),
    .A2(_14482_),
    .B1(_14449_),
    .Y(_18184_));
 sky130_fd_sc_hd__nand3_1 _47070_ (.A(_18182_),
    .B(_18183_),
    .C(_18184_),
    .Y(_18185_));
 sky130_fd_sc_hd__a21o_1 _47071_ (.A1(_18182_),
    .A2(_18183_),
    .B1(_18184_),
    .X(_18186_));
 sky130_fd_sc_hd__o2111ai_2 _47072_ (.A1(_03887_),
    .A2(_03909_),
    .B1(_14427_),
    .C1(_18185_),
    .D1(_18186_),
    .Y(_18187_));
 sky130_fd_sc_hd__nand2_1 _47073_ (.A(_18185_),
    .B(_18186_),
    .Y(_18188_));
 sky130_fd_sc_hd__o21ai_1 _47074_ (.A1(_03887_),
    .A2(_03909_),
    .B1(_14427_),
    .Y(_18189_));
 sky130_fd_sc_hd__nand2_1 _47075_ (.A(_18188_),
    .B(_18189_),
    .Y(_18190_));
 sky130_fd_sc_hd__nand3b_1 _47076_ (.A_N(_18168_),
    .B(_18187_),
    .C(_18190_),
    .Y(_18191_));
 sky130_fd_sc_hd__a21bo_1 _47077_ (.A1(_18187_),
    .A2(_18190_),
    .B1_N(_18168_),
    .X(_18192_));
 sky130_fd_sc_hd__a21o_1 _47078_ (.A1(_18191_),
    .A2(_18192_),
    .B1(_14537_),
    .X(_18193_));
 sky130_fd_sc_hd__nand3_1 _47079_ (.A(_18192_),
    .B(_14537_),
    .C(_18191_),
    .Y(_18194_));
 sky130_fd_sc_hd__a31o_1 _47080_ (.A1(_13965_),
    .A2(_13922_),
    .A3(_13943_),
    .B1(_13746_),
    .X(_18195_));
 sky130_fd_sc_hd__a21oi_1 _47081_ (.A1(_18193_),
    .A2(_18194_),
    .B1(_18195_),
    .Y(_18196_));
 sky130_fd_sc_hd__nand3_1 _47082_ (.A(_18195_),
    .B(_18193_),
    .C(_18194_),
    .Y(_18197_));
 sky130_fd_sc_hd__or2b_1 _47083_ (.A(_18196_),
    .B_N(_18197_),
    .X(_18198_));
 sky130_fd_sc_hd__o41a_2 _47084_ (.A1(_09393_),
    .A2(_09371_),
    .A3(_14537_),
    .A4(_14515_),
    .B1(_14581_),
    .X(_18199_));
 sky130_fd_sc_hd__o21bai_1 _47085_ (.A1(_14262_),
    .A2(_14592_),
    .B1_N(_09921_),
    .Y(_18200_));
 sky130_fd_sc_hd__a21boi_1 _47086_ (.A1(_14262_),
    .A2(_14592_),
    .B1_N(_18200_),
    .Y(_18201_));
 sky130_fd_sc_hd__a21boi_2 _47087_ (.A1(_18198_),
    .A2(_18199_),
    .B1_N(_18201_),
    .Y(_18202_));
 sky130_fd_sc_hd__xor2_1 _47088_ (.A(_18199_),
    .B(_18198_),
    .X(_18203_));
 sky130_fd_sc_hd__nor2_1 _47089_ (.A(_18201_),
    .B(_18203_),
    .Y(_18204_));
 sky130_fd_sc_hd__nand2_1 _47090_ (.A(_14075_),
    .B(_14053_),
    .Y(_18205_));
 sky130_fd_sc_hd__o211a_1 _47091_ (.A1(_18202_),
    .A2(_18204_),
    .B1(_14042_),
    .C1(_18205_),
    .X(_18206_));
 sky130_fd_sc_hd__a211oi_2 _47092_ (.A1(_14042_),
    .A2(_18205_),
    .B1(_18202_),
    .C1(_18204_),
    .Y(_18207_));
 sky130_fd_sc_hd__o22a_1 _47093_ (.A1(_09976_),
    .A2(_14603_),
    .B1(_18206_),
    .B2(_18207_),
    .X(_18208_));
 sky130_fd_sc_hd__nor4_1 _47094_ (.A(_09976_),
    .B(_18207_),
    .C(_14603_),
    .D(_18206_),
    .Y(_18209_));
 sky130_fd_sc_hd__nor2_2 _47095_ (.A(_18208_),
    .B(net98),
    .Y(_18210_));
 sky130_fd_sc_hd__a21oi_2 _47096_ (.A1(_18163_),
    .A2(_18167_),
    .B1(_18210_),
    .Y(_18211_));
 sky130_fd_sc_hd__nor2_1 _47097_ (.A(_14757_),
    .B(_14789_),
    .Y(_18212_));
 sky130_fd_sc_hd__a2111o_1 _47098_ (.A1(_03656_),
    .A2(_03755_),
    .B1(_09921_),
    .C1(_09932_),
    .D1(_14603_),
    .X(_18213_));
 sky130_fd_sc_hd__inv_2 _47099_ (.A(_18213_),
    .Y(_18214_));
 sky130_fd_sc_hd__o21a_1 _47100_ (.A1(_18206_),
    .A2(_18207_),
    .B1(_18214_),
    .X(_18215_));
 sky130_fd_sc_hd__clkbuf_2 _47101_ (.A(_18207_),
    .X(_18216_));
 sky130_fd_sc_hd__nor3_1 _47102_ (.A(_18214_),
    .B(_18206_),
    .C(_18216_),
    .Y(_18217_));
 sky130_fd_sc_hd__o211ai_2 _47103_ (.A1(_18215_),
    .A2(net94),
    .B1(_18162_),
    .C1(_18166_),
    .Y(_18218_));
 sky130_fd_sc_hd__o21ai_4 _47104_ (.A1(_14768_),
    .A2(_18212_),
    .B1(_18218_),
    .Y(_18219_));
 sky130_fd_sc_hd__o2bb2ai_1 _47105_ (.A1_N(_18162_),
    .A2_N(_18166_),
    .B1(_18215_),
    .B2(net94),
    .Y(_18220_));
 sky130_fd_sc_hd__a21oi_2 _47106_ (.A1(_14185_),
    .A2(_14691_),
    .B1(_14768_),
    .Y(_18221_));
 sky130_fd_sc_hd__o211ai_2 _47107_ (.A1(_18208_),
    .A2(net97),
    .B1(_18162_),
    .C1(_18167_),
    .Y(_18222_));
 sky130_fd_sc_hd__nand3_2 _47108_ (.A(_18220_),
    .B(_18221_),
    .C(_18222_),
    .Y(_18223_));
 sky130_fd_sc_hd__o21ai_2 _47109_ (.A1(_18211_),
    .A2(_18219_),
    .B1(_18223_),
    .Y(_18224_));
 sky130_fd_sc_hd__nand2_1 _47110_ (.A(_17907_),
    .B(_18224_),
    .Y(_18225_));
 sky130_fd_sc_hd__o2bb2a_2 _47111_ (.A1_N(_14844_),
    .A2_N(_14822_),
    .B1(_14735_),
    .B2(_14702_),
    .X(_18226_));
 sky130_fd_sc_hd__inv_2 _47112_ (.A(_17907_),
    .Y(_18227_));
 sky130_fd_sc_hd__o211ai_4 _47113_ (.A1(_18211_),
    .A2(_18219_),
    .B1(_18223_),
    .C1(_18227_),
    .Y(_18228_));
 sky130_fd_sc_hd__clkbuf_2 _47114_ (.A(_17907_),
    .X(_18229_));
 sky130_fd_sc_hd__clkbuf_2 _47115_ (.A(_18223_),
    .X(_18230_));
 sky130_fd_sc_hd__a31oi_4 _47116_ (.A1(_18163_),
    .A2(_18167_),
    .A3(_18210_),
    .B1(_18221_),
    .Y(_18231_));
 sky130_fd_sc_hd__a21o_1 _47117_ (.A1(_18163_),
    .A2(_18167_),
    .B1(_18210_),
    .X(_18232_));
 sky130_fd_sc_hd__nand2_2 _47118_ (.A(_18231_),
    .B(_18232_),
    .Y(_18233_));
 sky130_fd_sc_hd__a31oi_4 _47119_ (.A1(_18229_),
    .A2(_18230_),
    .A3(_18233_),
    .B1(_18226_),
    .Y(_18234_));
 sky130_fd_sc_hd__nand2_4 _47120_ (.A(_18224_),
    .B(_18227_),
    .Y(_18235_));
 sky130_fd_sc_hd__a32oi_4 _47121_ (.A1(_18225_),
    .A2(_18226_),
    .A3(_18228_),
    .B1(_18234_),
    .B2(_18235_),
    .Y(_18236_));
 sky130_fd_sc_hd__nand3_2 _47122_ (.A(_18225_),
    .B(_18226_),
    .C(_18228_),
    .Y(_18237_));
 sky130_fd_sc_hd__clkbuf_4 _47123_ (.A(_18237_),
    .X(_18238_));
 sky130_fd_sc_hd__nand2_2 _47124_ (.A(_17905_),
    .B(_18238_),
    .Y(_18239_));
 sky130_fd_sc_hd__o221ai_4 _47125_ (.A1(_17901_),
    .A2(_17903_),
    .B1(_17906_),
    .B2(_18236_),
    .C1(_18239_),
    .Y(_18240_));
 sky130_fd_sc_hd__o211ai_2 _47126_ (.A1(_18211_),
    .A2(_18219_),
    .B1(_18230_),
    .C1(_18229_),
    .Y(_18241_));
 sky130_fd_sc_hd__nand3b_4 _47127_ (.A_N(_18226_),
    .B(_18235_),
    .C(_18241_),
    .Y(_18242_));
 sky130_fd_sc_hd__a21oi_2 _47128_ (.A1(_18238_),
    .A2(_18242_),
    .B1(_17906_),
    .Y(_18243_));
 sky130_fd_sc_hd__and2_1 _47129_ (.A(_17905_),
    .B(_18238_),
    .X(_18244_));
 sky130_fd_sc_hd__nor2_1 _47130_ (.A(_17901_),
    .B(_17903_),
    .Y(_18245_));
 sky130_fd_sc_hd__o21ai_2 _47131_ (.A1(_18243_),
    .A2(_18244_),
    .B1(_18245_),
    .Y(_18246_));
 sky130_fd_sc_hd__a2bb2oi_4 _47132_ (.A1_N(_17800_),
    .A2_N(_17804_),
    .B1(_18240_),
    .B2(_18246_),
    .Y(_18247_));
 sky130_fd_sc_hd__o221a_2 _47133_ (.A1(_15031_),
    .A2(_17896_),
    .B1(_10405_),
    .B2(_14899_),
    .C1(_14987_),
    .X(_18248_));
 sky130_fd_sc_hd__a21o_1 _47134_ (.A1(_18238_),
    .A2(_18242_),
    .B1(_17906_),
    .X(_18249_));
 sky130_fd_sc_hd__or2_2 _47135_ (.A(_17901_),
    .B(_17902_),
    .X(_18250_));
 sky130_fd_sc_hd__a21oi_4 _47136_ (.A1(_18249_),
    .A2(_18239_),
    .B1(_18250_),
    .Y(_18251_));
 sky130_fd_sc_hd__a21oi_1 _47137_ (.A1(_17783_),
    .A2(_17799_),
    .B1(_17804_),
    .Y(_18252_));
 sky130_fd_sc_hd__nand2_2 _47138_ (.A(_18240_),
    .B(_18252_),
    .Y(_18253_));
 sky130_fd_sc_hd__o22ai_4 _47139_ (.A1(_15020_),
    .A2(_18248_),
    .B1(_18251_),
    .B2(_18253_),
    .Y(_18254_));
 sky130_fd_sc_hd__o21ai_2 _47140_ (.A1(_18243_),
    .A2(_18244_),
    .B1(_18250_),
    .Y(_18255_));
 sky130_fd_sc_hd__o211ai_2 _47141_ (.A1(_17906_),
    .A2(_18236_),
    .B1(_18239_),
    .C1(_18245_),
    .Y(_18256_));
 sky130_fd_sc_hd__o211ai_4 _47142_ (.A1(_17800_),
    .A2(_17804_),
    .B1(_18255_),
    .C1(_18256_),
    .Y(_18257_));
 sky130_fd_sc_hd__nand3_2 _47143_ (.A(_18246_),
    .B(_18252_),
    .C(_18240_),
    .Y(_18258_));
 sky130_fd_sc_hd__buf_2 _47144_ (.A(_15031_),
    .X(_18259_));
 sky130_fd_sc_hd__a21o_1 _47145_ (.A1(_18259_),
    .A2(_17896_),
    .B1(_18248_),
    .X(_18260_));
 sky130_fd_sc_hd__a21o_1 _47146_ (.A1(_18257_),
    .A2(_18258_),
    .B1(_18260_),
    .X(_18261_));
 sky130_fd_sc_hd__o221ai_4 _47147_ (.A1(_17767_),
    .A2(_17807_),
    .B1(_18247_),
    .B2(_18254_),
    .C1(_18261_),
    .Y(_18262_));
 sky130_fd_sc_hd__a21oi_4 _47148_ (.A1(_18257_),
    .A2(_18258_),
    .B1(_18260_),
    .Y(_18263_));
 sky130_fd_sc_hd__o221a_1 _47149_ (.A1(_15020_),
    .A2(_18248_),
    .B1(_18251_),
    .B2(_18253_),
    .C1(_18257_),
    .X(_18264_));
 sky130_fd_sc_hd__a31o_1 _47150_ (.A1(_17488_),
    .A2(_17758_),
    .A3(_17765_),
    .B1(_17807_),
    .X(_18265_));
 sky130_fd_sc_hd__o21bai_4 _47151_ (.A1(_18263_),
    .A2(_18264_),
    .B1_N(_18265_),
    .Y(_18266_));
 sky130_fd_sc_hd__a21o_2 _47152_ (.A1(_15207_),
    .A2(_15174_),
    .B1(_15119_),
    .X(_18267_));
 sky130_fd_sc_hd__a21oi_4 _47153_ (.A1(_18262_),
    .A2(_18266_),
    .B1(_18267_),
    .Y(_18268_));
 sky130_fd_sc_hd__o221ai_4 _47154_ (.A1(_15020_),
    .A2(_18248_),
    .B1(_18251_),
    .B2(_18253_),
    .C1(_18257_),
    .Y(_18269_));
 sky130_fd_sc_hd__a21oi_4 _47155_ (.A1(_18261_),
    .A2(_18269_),
    .B1(_18265_),
    .Y(_18270_));
 sky130_fd_sc_hd__o22ai_4 _47156_ (.A1(_17767_),
    .A2(_17807_),
    .B1(_18247_),
    .B2(_18254_),
    .Y(_18271_));
 sky130_fd_sc_hd__o21ai_4 _47157_ (.A1(_18263_),
    .A2(_18271_),
    .B1(_18267_),
    .Y(_18272_));
 sky130_fd_sc_hd__o2bb2ai_4 _47158_ (.A1_N(_15328_),
    .A2_N(_15339_),
    .B1(_18270_),
    .B2(_18272_),
    .Y(_18273_));
 sky130_fd_sc_hd__inv_2 _47159_ (.A(_15229_),
    .Y(_18274_));
 sky130_fd_sc_hd__nor2_2 _47160_ (.A(_18263_),
    .B(_18271_),
    .Y(_18275_));
 sky130_fd_sc_hd__o22ai_2 _47161_ (.A1(_15119_),
    .A2(_18274_),
    .B1(_18275_),
    .B2(_18270_),
    .Y(_18276_));
 sky130_fd_sc_hd__a21oi_2 _47162_ (.A1(_15284_),
    .A2(_15317_),
    .B1(_15273_),
    .Y(_18277_));
 sky130_fd_sc_hd__o2111ai_4 _47163_ (.A1(_18271_),
    .A2(_18263_),
    .B1(_15229_),
    .C1(_15196_),
    .D1(_18266_),
    .Y(_18278_));
 sky130_fd_sc_hd__nand3_4 _47164_ (.A(_18276_),
    .B(_18277_),
    .C(_18278_),
    .Y(_18279_));
 sky130_fd_sc_hd__o21ai_1 _47165_ (.A1(_18268_),
    .A2(_18273_),
    .B1(_18279_),
    .Y(_18280_));
 sky130_fd_sc_hd__o21ai_1 _47166_ (.A1(_17899_),
    .A2(_17900_),
    .B1(_18280_),
    .Y(_18281_));
 sky130_fd_sc_hd__a21o_1 _47167_ (.A1(_17477_),
    .A2(_17862_),
    .B1(_17864_),
    .X(_18282_));
 sky130_fd_sc_hd__inv_2 _47168_ (.A(_18282_),
    .Y(_18283_));
 sky130_fd_sc_hd__nor2_1 _47169_ (.A(_17899_),
    .B(_17900_),
    .Y(_18284_));
 sky130_fd_sc_hd__o211ai_1 _47170_ (.A1(_18268_),
    .A2(_18273_),
    .B1(_18279_),
    .C1(_18284_),
    .Y(_18285_));
 sky130_fd_sc_hd__nand3_2 _47171_ (.A(_18281_),
    .B(_18283_),
    .C(_18285_),
    .Y(_18286_));
 sky130_fd_sc_hd__o22ai_1 _47172_ (.A1(_17899_),
    .A2(_17900_),
    .B1(_18268_),
    .B2(_18273_),
    .Y(_18287_));
 sky130_fd_sc_hd__and3_2 _47173_ (.A(_18276_),
    .B(_18277_),
    .C(_18278_),
    .X(_18288_));
 sky130_fd_sc_hd__nand2_1 _47174_ (.A(_18284_),
    .B(_18280_),
    .Y(_18289_));
 sky130_fd_sc_hd__o211ai_2 _47175_ (.A1(_18287_),
    .A2(_18288_),
    .B1(_18282_),
    .C1(_18289_),
    .Y(_18290_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47176_ (.A(_18290_),
    .X(_18291_));
 sky130_fd_sc_hd__a21oi_2 _47177_ (.A1(_15394_),
    .A2(_15416_),
    .B1(_15361_),
    .Y(_18292_));
 sky130_fd_sc_hd__a21oi_1 _47178_ (.A1(_18286_),
    .A2(_18291_),
    .B1(_18292_),
    .Y(_18293_));
 sky130_fd_sc_hd__o211a_1 _47179_ (.A1(_18273_),
    .A2(_18268_),
    .B1(_18284_),
    .C1(_18279_),
    .X(_18294_));
 sky130_fd_sc_hd__and3_1 _47180_ (.A(_15284_),
    .B(_15317_),
    .C(_15328_),
    .X(_18295_));
 sky130_fd_sc_hd__o21bai_2 _47181_ (.A1(_18275_),
    .A2(_18270_),
    .B1_N(_18267_),
    .Y(_18296_));
 sky130_fd_sc_hd__o221ai_4 _47182_ (.A1(_18270_),
    .A2(_18272_),
    .B1(_15273_),
    .B2(_18295_),
    .C1(_18296_),
    .Y(_18297_));
 sky130_fd_sc_hd__a21oi_1 _47183_ (.A1(_18279_),
    .A2(_18297_),
    .B1(_18284_),
    .Y(_18298_));
 sky130_fd_sc_hd__o311a_1 _47184_ (.A1(_18282_),
    .A2(_18294_),
    .A3(_18298_),
    .B1(_18290_),
    .C1(_18292_),
    .X(_18299_));
 sky130_fd_sc_hd__a22o_1 _47185_ (.A1(_17379_),
    .A2(_17401_),
    .B1(_17434_),
    .B2(_16316_),
    .X(_18300_));
 sky130_fd_sc_hd__inv_2 _47186_ (.A(_16996_),
    .Y(_18301_));
 sky130_fd_sc_hd__nand4_1 _47187_ (.A(_17117_),
    .B(_17128_),
    .C(_17281_),
    .D(_17292_),
    .Y(_18302_));
 sky130_fd_sc_hd__nor2_1 _47188_ (.A(_16481_),
    .B(net173),
    .Y(_18303_));
 sky130_fd_sc_hd__inv_2 _47189_ (.A(net346),
    .Y(_18304_));
 sky130_fd_sc_hd__clkbuf_2 _47190_ (.A(_18304_),
    .X(_18305_));
 sky130_fd_sc_hd__inv_2 _47191_ (.A(_01435_),
    .Y(_18306_));
 sky130_fd_sc_hd__nand2_1 _47192_ (.A(_18305_),
    .B(_18306_),
    .Y(_18307_));
 sky130_fd_sc_hd__nand2_2 _47193_ (.A(net346),
    .B(_01446_),
    .Y(_18308_));
 sky130_fd_sc_hd__buf_1 _47194_ (.A(net343),
    .X(_18309_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47195_ (.A(_18309_),
    .X(_18310_));
 sky130_fd_sc_hd__a21o_1 _47196_ (.A1(_18307_),
    .A2(_18308_),
    .B1(_18310_),
    .X(_18311_));
 sky130_fd_sc_hd__nand3_1 _47197_ (.A(_18307_),
    .B(_18308_),
    .C(_18310_),
    .Y(_18312_));
 sky130_fd_sc_hd__clkbuf_2 _47198_ (.A(_18312_),
    .X(_18313_));
 sky130_fd_sc_hd__nand4_2 _47199_ (.A(_18311_),
    .B(_17029_),
    .C(_23687_),
    .D(_18313_),
    .Y(_18314_));
 sky130_fd_sc_hd__a22o_1 _47200_ (.A1(_23698_),
    .A2(_17040_),
    .B1(_18313_),
    .B2(_18311_),
    .X(_18315_));
 sky130_fd_sc_hd__clkbuf_2 _47201_ (.A(\delay_line[22][4] ),
    .X(_18316_));
 sky130_fd_sc_hd__buf_1 _47202_ (.A(_18316_),
    .X(_18317_));
 sky130_fd_sc_hd__buf_2 _47203_ (.A(_18317_),
    .X(_18318_));
 sky130_fd_sc_hd__xor2_1 _47204_ (.A(_23676_),
    .B(_18318_),
    .X(_18319_));
 sky130_fd_sc_hd__a21oi_1 _47205_ (.A1(_18314_),
    .A2(_18315_),
    .B1(_18319_),
    .Y(_18320_));
 sky130_fd_sc_hd__and3_1 _47206_ (.A(_18315_),
    .B(_18319_),
    .C(_18314_),
    .X(_18321_));
 sky130_fd_sc_hd__clkbuf_2 _47207_ (.A(_17215_),
    .X(_18322_));
 sky130_fd_sc_hd__clkbuf_2 _47208_ (.A(\delay_line[25][5] ),
    .X(_18323_));
 sky130_fd_sc_hd__buf_1 _47209_ (.A(_18323_),
    .X(_18324_));
 sky130_fd_sc_hd__nor2_1 _47210_ (.A(_06766_),
    .B(_18324_),
    .Y(_18325_));
 sky130_fd_sc_hd__and2_1 _47211_ (.A(\delay_line[25][3] ),
    .B(\delay_line[25][5] ),
    .X(_18326_));
 sky130_fd_sc_hd__or4bb_4 _47212_ (.A(_18325_),
    .B(_18326_),
    .C_N(_17139_),
    .D_N(_17248_),
    .X(_18327_));
 sky130_fd_sc_hd__a2bb2o_1 _47213_ (.A1_N(_18325_),
    .A2_N(_18326_),
    .B1(_01490_),
    .B2(_17248_),
    .X(_18328_));
 sky130_fd_sc_hd__a21o_1 _47214_ (.A1(_18327_),
    .A2(_18328_),
    .B1(_22358_),
    .X(_18329_));
 sky130_fd_sc_hd__nand3_1 _47215_ (.A(_18327_),
    .B(_18328_),
    .C(_22358_),
    .Y(_18330_));
 sky130_fd_sc_hd__clkbuf_2 _47216_ (.A(_18330_),
    .X(_18331_));
 sky130_fd_sc_hd__nand4_1 _47217_ (.A(_17270_),
    .B(_18329_),
    .C(_17193_),
    .D(_18331_),
    .Y(_18332_));
 sky130_fd_sc_hd__buf_1 _47218_ (.A(_18332_),
    .X(_18333_));
 sky130_fd_sc_hd__a32o_1 _47219_ (.A1(_23742_),
    .A2(_17270_),
    .A3(_06799_),
    .B1(_18329_),
    .B2(_18331_),
    .X(_18334_));
 sky130_fd_sc_hd__a2bb2o_1 _47220_ (.A1_N(_06854_),
    .A2_N(_18322_),
    .B1(_18333_),
    .B2(_18334_),
    .X(_18335_));
 sky130_fd_sc_hd__or4bb_2 _47221_ (.A(_18322_),
    .B(_06854_),
    .C_N(_18334_),
    .D_N(_18333_),
    .X(_18336_));
 sky130_fd_sc_hd__and4bb_1 _47222_ (.A_N(_18320_),
    .B_N(_18321_),
    .C(_18335_),
    .D(_18336_),
    .X(_18337_));
 sky130_fd_sc_hd__a2bb2oi_1 _47223_ (.A1_N(_18320_),
    .A2_N(_18321_),
    .B1(_18335_),
    .B2(_18336_),
    .Y(_18338_));
 sky130_fd_sc_hd__nor2_1 _47224_ (.A(_18337_),
    .B(_18338_),
    .Y(_18339_));
 sky130_fd_sc_hd__xor2_1 _47225_ (.A(_18303_),
    .B(_18339_),
    .X(_18340_));
 sky130_fd_sc_hd__a21oi_2 _47226_ (.A1(_17128_),
    .A2(_18302_),
    .B1(_18340_),
    .Y(_18341_));
 sky130_fd_sc_hd__o311a_1 _47227_ (.A1(_17106_),
    .A2(_17051_),
    .A3(_17062_),
    .B1(_18302_),
    .C1(_18340_),
    .X(_18342_));
 sky130_fd_sc_hd__nor2_2 _47228_ (.A(_18341_),
    .B(_18342_),
    .Y(_18343_));
 sky130_fd_sc_hd__inv_2 _47229_ (.A(_16941_),
    .Y(_18344_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47230_ (.A(\delay_line[21][3] ),
    .X(_18345_));
 sky130_fd_sc_hd__and2b_1 _47231_ (.A_N(net361),
    .B(_18345_),
    .X(_18346_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47232_ (.A(net360),
    .X(_18347_));
 sky130_fd_sc_hd__clkbuf_2 _47233_ (.A(_18347_),
    .X(_18348_));
 sky130_fd_sc_hd__buf_1 _47234_ (.A(_18348_),
    .X(_18349_));
 sky130_fd_sc_hd__clkbuf_2 _47235_ (.A(_18349_),
    .X(_18350_));
 sky130_fd_sc_hd__clkbuf_2 _47236_ (.A(_18350_),
    .X(_18351_));
 sky130_fd_sc_hd__clkbuf_2 _47237_ (.A(_16503_),
    .X(_18352_));
 sky130_fd_sc_hd__buf_1 _47238_ (.A(_18352_),
    .X(_18353_));
 sky130_fd_sc_hd__and3b_1 _47239_ (.A_N(_18353_),
    .B(_07580_),
    .C(_07294_),
    .X(_18354_));
 sky130_fd_sc_hd__nand2_1 _47240_ (.A(_18351_),
    .B(_18354_),
    .Y(_18355_));
 sky130_fd_sc_hd__or2b_1 _47241_ (.A(_18345_),
    .B_N(_18347_),
    .X(_18356_));
 sky130_fd_sc_hd__or2b_1 _47242_ (.A(net360),
    .B_N(_18345_),
    .X(_18357_));
 sky130_fd_sc_hd__nand2_1 _47243_ (.A(_18356_),
    .B(_18357_),
    .Y(_18358_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47244_ (.A(_18358_),
    .X(_18359_));
 sky130_fd_sc_hd__nand2_1 _47245_ (.A(_18353_),
    .B(_07580_),
    .Y(_18360_));
 sky130_fd_sc_hd__clkbuf_2 _47246_ (.A(_18353_),
    .X(_18361_));
 sky130_fd_sc_hd__o2111a_1 _47247_ (.A1(_16492_),
    .A2(_18361_),
    .B1(_07602_),
    .C1(_18356_),
    .D1(_18357_),
    .X(_18362_));
 sky130_fd_sc_hd__a21o_1 _47248_ (.A1(_18359_),
    .A2(_18360_),
    .B1(_18362_),
    .X(_18363_));
 sky130_fd_sc_hd__a32o_1 _47249_ (.A1(_24017_),
    .A2(_16492_),
    .A3(_18346_),
    .B1(_18355_),
    .B2(_18363_),
    .X(_18364_));
 sky130_fd_sc_hd__or4b_1 _47250_ (.A(_07591_),
    .B(_18350_),
    .C(_07349_),
    .D_N(_18353_),
    .X(_18365_));
 sky130_fd_sc_hd__buf_1 _47251_ (.A(_18365_),
    .X(_18366_));
 sky130_fd_sc_hd__clkbuf_2 _47252_ (.A(\delay_line[19][3] ),
    .X(_18367_));
 sky130_fd_sc_hd__buf_2 _47253_ (.A(_18367_),
    .X(_18368_));
 sky130_fd_sc_hd__and3b_1 _47254_ (.A_N(_18368_),
    .B(_07459_),
    .C(_07415_),
    .X(_18369_));
 sky130_fd_sc_hd__inv_2 _47255_ (.A(net371),
    .Y(_18370_));
 sky130_fd_sc_hd__nand2_1 _47256_ (.A(_18370_),
    .B(_16382_),
    .Y(_18371_));
 sky130_fd_sc_hd__or2b_1 _47257_ (.A(_16382_),
    .B_N(net371),
    .X(_18372_));
 sky130_fd_sc_hd__nand2_1 _47258_ (.A(_18371_),
    .B(_18372_),
    .Y(_18373_));
 sky130_fd_sc_hd__clkbuf_2 _47259_ (.A(\delay_line[19][4] ),
    .X(_18374_));
 sky130_fd_sc_hd__buf_1 _47260_ (.A(_18374_),
    .X(_18375_));
 sky130_fd_sc_hd__buf_1 _47261_ (.A(_18375_),
    .X(_18376_));
 sky130_fd_sc_hd__and2_1 _47262_ (.A(_18367_),
    .B(_07382_),
    .X(_18377_));
 sky130_fd_sc_hd__mux2_1 _47263_ (.A0(_18373_),
    .A1(_18376_),
    .S(_18377_),
    .X(_18378_));
 sky130_fd_sc_hd__o2111a_2 _47264_ (.A1(_18369_),
    .A2(_18378_),
    .B1(_23896_),
    .C1(_07426_),
    .D1(_16404_),
    .X(_18379_));
 sky130_fd_sc_hd__buf_1 _47265_ (.A(_18368_),
    .X(_18380_));
 sky130_fd_sc_hd__and4b_1 _47266_ (.A_N(_18380_),
    .B(_07459_),
    .C(_18376_),
    .D(_07415_),
    .X(_18381_));
 sky130_fd_sc_hd__o21ba_1 _47267_ (.A1(_18369_),
    .A2(_18378_),
    .B1_N(_18381_),
    .X(_18382_));
 sky130_fd_sc_hd__a31oi_4 _47268_ (.A1(_23907_),
    .A2(_07426_),
    .A3(_16404_),
    .B1(_18382_),
    .Y(_18383_));
 sky130_fd_sc_hd__buf_1 _47269_ (.A(\delay_line[18][4] ),
    .X(_18384_));
 sky130_fd_sc_hd__buf_2 _47270_ (.A(_18384_),
    .X(_18385_));
 sky130_fd_sc_hd__nor2_1 _47271_ (.A(_23863_),
    .B(_18385_),
    .Y(_18386_));
 sky130_fd_sc_hd__inv_2 _47272_ (.A(\delay_line[18][4] ),
    .Y(_18387_));
 sky130_fd_sc_hd__clkbuf_2 _47273_ (.A(_18387_),
    .X(_18388_));
 sky130_fd_sc_hd__clkbuf_2 _47274_ (.A(_18388_),
    .X(_18389_));
 sky130_fd_sc_hd__nor2_1 _47275_ (.A(_23951_),
    .B(_18389_),
    .Y(_18390_));
 sky130_fd_sc_hd__o22ai_4 _47276_ (.A1(_18379_),
    .A2(_18383_),
    .B1(_18386_),
    .B2(_18390_),
    .Y(_18391_));
 sky130_fd_sc_hd__or4_1 _47277_ (.A(_18379_),
    .B(_18383_),
    .C(_18386_),
    .D(_18390_),
    .X(_18392_));
 sky130_fd_sc_hd__nand2_1 _47278_ (.A(_18391_),
    .B(_18392_),
    .Y(_18393_));
 sky130_fd_sc_hd__a21bo_2 _47279_ (.A1(_18364_),
    .A2(_18366_),
    .B1_N(_18392_),
    .X(_18394_));
 sky130_fd_sc_hd__inv_2 _47280_ (.A(_18394_),
    .Y(_18395_));
 sky130_fd_sc_hd__a32o_1 _47281_ (.A1(_18364_),
    .A2(_18366_),
    .A3(_18393_),
    .B1(_18395_),
    .B2(_18391_),
    .X(_18396_));
 sky130_fd_sc_hd__or2_1 _47282_ (.A(\delay_line[16][0] ),
    .B(_01864_),
    .X(_18397_));
 sky130_fd_sc_hd__nand2_1 _47283_ (.A(_24127_),
    .B(_01875_),
    .Y(_18398_));
 sky130_fd_sc_hd__buf_1 _47284_ (.A(\delay_line[16][4] ),
    .X(_18399_));
 sky130_fd_sc_hd__clkbuf_2 _47285_ (.A(_18399_),
    .X(_18400_));
 sky130_fd_sc_hd__nand3_2 _47286_ (.A(_18397_),
    .B(_18398_),
    .C(_18400_),
    .Y(_18401_));
 sky130_fd_sc_hd__a21o_1 _47287_ (.A1(_18397_),
    .A2(_18398_),
    .B1(_18400_),
    .X(_18402_));
 sky130_fd_sc_hd__a22o_1 _47288_ (.A1(_24138_),
    .A2(_16612_),
    .B1(_18401_),
    .B2(_18402_),
    .X(_18403_));
 sky130_fd_sc_hd__nand4_4 _47289_ (.A(_18402_),
    .B(_16612_),
    .C(_24127_),
    .D(_18401_),
    .Y(_18404_));
 sky130_fd_sc_hd__buf_1 _47290_ (.A(\delay_line[14][4] ),
    .X(_18405_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47291_ (.A(_18405_),
    .X(_18406_));
 sky130_fd_sc_hd__clkbuf_2 _47292_ (.A(_18406_),
    .X(_18407_));
 sky130_fd_sc_hd__clkbuf_2 _47293_ (.A(_18407_),
    .X(_18408_));
 sky130_fd_sc_hd__and2_1 _47294_ (.A(_24072_),
    .B(_18408_),
    .X(_18409_));
 sky130_fd_sc_hd__nor2_1 _47295_ (.A(_24072_),
    .B(_18408_),
    .Y(_18410_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47296_ (.A(_16733_),
    .X(_18411_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47297_ (.A(_18411_),
    .X(_18412_));
 sky130_fd_sc_hd__clkbuf_2 _47298_ (.A(_18412_),
    .X(_18413_));
 sky130_fd_sc_hd__buf_1 _47299_ (.A(\delay_line[15][5] ),
    .X(_18414_));
 sky130_fd_sc_hd__and2_1 _47300_ (.A(\delay_line[15][3] ),
    .B(_18414_),
    .X(_18415_));
 sky130_fd_sc_hd__buf_2 _47301_ (.A(_18414_),
    .X(_18416_));
 sky130_fd_sc_hd__o211ai_2 _47302_ (.A1(\delay_line[15][3] ),
    .A2(_18416_),
    .B1(_01787_),
    .C1(_16733_),
    .Y(_18417_));
 sky130_fd_sc_hd__nor2_1 _47303_ (.A(\delay_line[15][3] ),
    .B(_18414_),
    .Y(_18418_));
 sky130_fd_sc_hd__a2bb2o_1 _47304_ (.A1_N(_18415_),
    .A2_N(_18418_),
    .B1(_01787_),
    .B2(_16733_),
    .X(_18419_));
 sky130_fd_sc_hd__o211a_1 _47305_ (.A1(_18415_),
    .A2(_18417_),
    .B1(_22391_),
    .C1(_18419_),
    .X(_18420_));
 sky130_fd_sc_hd__clkbuf_2 _47306_ (.A(_18420_),
    .X(_18421_));
 sky130_fd_sc_hd__buf_1 _47307_ (.A(_18416_),
    .X(_18422_));
 sky130_fd_sc_hd__buf_1 _47308_ (.A(_18422_),
    .X(_18423_));
 sky130_fd_sc_hd__a21o_1 _47309_ (.A1(_07096_),
    .A2(_18423_),
    .B1(_18417_),
    .X(_18424_));
 sky130_fd_sc_hd__a21oi_1 _47310_ (.A1(_18424_),
    .A2(_18419_),
    .B1(_22402_),
    .Y(_18425_));
 sky130_fd_sc_hd__o2bb2a_1 _47311_ (.A1_N(_16766_),
    .A2_N(_16799_),
    .B1(_18421_),
    .B2(_18425_),
    .X(_18426_));
 sky130_fd_sc_hd__a2111oi_1 _47312_ (.A1(_16711_),
    .A2(_16755_),
    .B1(_16854_),
    .C1(_18421_),
    .D1(_18425_),
    .Y(_18427_));
 sky130_fd_sc_hd__o22ai_1 _47313_ (.A1(_07151_),
    .A2(_18413_),
    .B1(_18426_),
    .B2(net182),
    .Y(_18428_));
 sky130_fd_sc_hd__clkbuf_2 _47314_ (.A(_16689_),
    .X(_18429_));
 sky130_fd_sc_hd__o211a_1 _47315_ (.A1(_07085_),
    .A2(_07129_),
    .B1(_18429_),
    .C1(_01809_),
    .X(_18430_));
 sky130_fd_sc_hd__a2111o_2 _47316_ (.A1(_16711_),
    .A2(_16755_),
    .B1(_16854_),
    .C1(_18421_),
    .D1(_18425_),
    .X(_18431_));
 sky130_fd_sc_hd__nand3b_2 _47317_ (.A_N(_18426_),
    .B(_18430_),
    .C(_18431_),
    .Y(_18432_));
 sky130_fd_sc_hd__or4bb_4 _47318_ (.A(_18409_),
    .B(_18410_),
    .C_N(_18428_),
    .D_N(_18432_),
    .X(_18433_));
 sky130_fd_sc_hd__a2bb2o_2 _47319_ (.A1_N(_18409_),
    .A2_N(_18410_),
    .B1(_18428_),
    .B2(_18432_),
    .X(_18434_));
 sky130_fd_sc_hd__and4_1 _47320_ (.A(_18403_),
    .B(_18404_),
    .C(_18433_),
    .D(_18434_),
    .X(_18435_));
 sky130_fd_sc_hd__a22oi_4 _47321_ (.A1(_18403_),
    .A2(_18404_),
    .B1(_18433_),
    .B2(_18434_),
    .Y(_18436_));
 sky130_fd_sc_hd__nand3_2 _47322_ (.A(_16810_),
    .B(_16843_),
    .C(_16865_),
    .Y(_18437_));
 sky130_fd_sc_hd__o211ai_4 _47323_ (.A1(_18435_),
    .A2(_18436_),
    .B1(_18437_),
    .C1(_16898_),
    .Y(_18438_));
 sky130_fd_sc_hd__a211o_2 _47324_ (.A1(_18437_),
    .A2(_16898_),
    .B1(_18435_),
    .C1(_18436_),
    .X(_18439_));
 sky130_fd_sc_hd__and3b_1 _47325_ (.A_N(_18396_),
    .B(_18438_),
    .C(_18439_),
    .X(_18440_));
 sky130_fd_sc_hd__a21boi_1 _47326_ (.A1(_18438_),
    .A2(_18439_),
    .B1_N(_18396_),
    .Y(_18441_));
 sky130_fd_sc_hd__nor2_1 _47327_ (.A(_18440_),
    .B(_18441_),
    .Y(_18442_));
 sky130_fd_sc_hd__o311a_1 _47328_ (.A1(_16568_),
    .A2(_16579_),
    .A3(_16930_),
    .B1(_18344_),
    .C1(_18442_),
    .X(_18443_));
 sky130_fd_sc_hd__a21oi_2 _47329_ (.A1(_18344_),
    .A2(_16952_),
    .B1(_18442_),
    .Y(_18444_));
 sky130_fd_sc_hd__nor2_1 _47330_ (.A(_18443_),
    .B(_18444_),
    .Y(_18445_));
 sky130_fd_sc_hd__and2_1 _47331_ (.A(_18343_),
    .B(_18445_),
    .X(_18446_));
 sky130_fd_sc_hd__nor2_1 _47332_ (.A(_18343_),
    .B(_18445_),
    .Y(_18447_));
 sky130_fd_sc_hd__or2_1 _47333_ (.A(_18446_),
    .B(_18447_),
    .X(_18448_));
 sky130_fd_sc_hd__a21oi_1 _47334_ (.A1(_18301_),
    .A2(_17412_),
    .B1(_18448_),
    .Y(_18449_));
 sky130_fd_sc_hd__inv_2 _47335_ (.A(\delay_line[29][3] ),
    .Y(_18450_));
 sky130_fd_sc_hd__clkbuf_2 _47336_ (.A(_18450_),
    .X(_18451_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47337_ (.A(\delay_line[30][5] ),
    .X(_18452_));
 sky130_fd_sc_hd__clkbuf_2 _47338_ (.A(_18452_),
    .X(_18453_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47339_ (.A(\delay_line[30][2] ),
    .X(_18454_));
 sky130_fd_sc_hd__and2b_1 _47340_ (.A_N(_18454_),
    .B(\delay_line[30][0] ),
    .X(_18455_));
 sky130_fd_sc_hd__and2b_1 _47341_ (.A_N(_22281_),
    .B(_18454_),
    .X(_18456_));
 sky130_fd_sc_hd__nor3_2 _47342_ (.A(_18453_),
    .B(_18455_),
    .C(_18456_),
    .Y(_18457_));
 sky130_fd_sc_hd__o21a_1 _47343_ (.A1(_18455_),
    .A2(_18456_),
    .B1(_18452_),
    .X(_18458_));
 sky130_fd_sc_hd__or4_2 _47344_ (.A(_15602_),
    .B(_15624_),
    .C(_18457_),
    .D(_18458_),
    .X(_18459_));
 sky130_fd_sc_hd__o22ai_4 _47345_ (.A1(_15602_),
    .A2(_15624_),
    .B1(_18457_),
    .B2(_18458_),
    .Y(_18460_));
 sky130_fd_sc_hd__and3_1 _47346_ (.A(_18451_),
    .B(_18459_),
    .C(_18460_),
    .X(_18461_));
 sky130_fd_sc_hd__a21oi_4 _47347_ (.A1(_18459_),
    .A2(_18460_),
    .B1(_18451_),
    .Y(_18462_));
 sky130_fd_sc_hd__nor2_2 _47348_ (.A(_18461_),
    .B(_18462_),
    .Y(_18463_));
 sky130_fd_sc_hd__or3b_1 _47349_ (.A(_15844_),
    .B(_15866_),
    .C_N(_15767_),
    .X(_18464_));
 sky130_fd_sc_hd__buf_1 _47350_ (.A(\delay_line[31][5] ),
    .X(_18465_));
 sky130_fd_sc_hd__nor2_1 _47351_ (.A(net318),
    .B(_18465_),
    .Y(_18466_));
 sky130_fd_sc_hd__nand2_1 _47352_ (.A(_15789_),
    .B(_18465_),
    .Y(_18467_));
 sky130_fd_sc_hd__nand3b_1 _47353_ (.A_N(_18466_),
    .B(_18467_),
    .C(_06205_),
    .Y(_18468_));
 sky130_fd_sc_hd__and2_1 _47354_ (.A(net318),
    .B(_18465_),
    .X(_18469_));
 sky130_fd_sc_hd__o21ai_1 _47355_ (.A1(_18466_),
    .A2(_18469_),
    .B1(_06249_),
    .Y(_18470_));
 sky130_fd_sc_hd__o21ai_1 _47356_ (.A1(_15701_),
    .A2(_15778_),
    .B1(_15800_),
    .Y(_18471_));
 sky130_fd_sc_hd__and3_1 _47357_ (.A(_18468_),
    .B(_18470_),
    .C(_18471_),
    .X(_18472_));
 sky130_fd_sc_hd__nand2_1 _47358_ (.A(_18468_),
    .B(_18470_),
    .Y(_18473_));
 sky130_fd_sc_hd__and3_1 _47359_ (.A(_15800_),
    .B(_15811_),
    .C(_18473_),
    .X(_18474_));
 sky130_fd_sc_hd__nor2_1 _47360_ (.A(_18472_),
    .B(_18474_),
    .Y(_18475_));
 sky130_fd_sc_hd__nor2_1 _47361_ (.A(_15844_),
    .B(_15855_),
    .Y(_18476_));
 sky130_fd_sc_hd__a21oi_1 _47362_ (.A1(_15756_),
    .A2(_18476_),
    .B1(_15866_),
    .Y(_18477_));
 sky130_fd_sc_hd__nand2_1 _47363_ (.A(_18475_),
    .B(_18477_),
    .Y(_18478_));
 sky130_fd_sc_hd__o21bai_1 _47364_ (.A1(_18472_),
    .A2(_18474_),
    .B1_N(_18477_),
    .Y(_18479_));
 sky130_fd_sc_hd__and3_1 _47365_ (.A(_18464_),
    .B(_18478_),
    .C(_18479_),
    .X(_18480_));
 sky130_fd_sc_hd__a21oi_2 _47366_ (.A1(_18478_),
    .A2(_18479_),
    .B1(_18464_),
    .Y(_18481_));
 sky130_fd_sc_hd__nor2_2 _47367_ (.A(_18480_),
    .B(_18481_),
    .Y(_18482_));
 sky130_fd_sc_hd__and2_2 _47368_ (.A(_18463_),
    .B(_18482_),
    .X(_18483_));
 sky130_fd_sc_hd__nor2_1 _47369_ (.A(_18463_),
    .B(_18482_),
    .Y(_18484_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47370_ (.A(\delay_line[26][0] ),
    .X(_18485_));
 sky130_fd_sc_hd__clkbuf_2 _47371_ (.A(\delay_line[26][4] ),
    .X(_18486_));
 sky130_fd_sc_hd__nor2_2 _47372_ (.A(_18485_),
    .B(_18486_),
    .Y(_18487_));
 sky130_fd_sc_hd__buf_1 _47373_ (.A(\delay_line[26][4] ),
    .X(_18488_));
 sky130_fd_sc_hd__and2_1 _47374_ (.A(_18485_),
    .B(_18488_),
    .X(_18489_));
 sky130_fd_sc_hd__buf_1 _47375_ (.A(_18489_),
    .X(_18490_));
 sky130_fd_sc_hd__clkbuf_2 _47376_ (.A(net333),
    .X(_18491_));
 sky130_fd_sc_hd__nor2_1 _47377_ (.A(\delay_line[27][3] ),
    .B(_18491_),
    .Y(_18492_));
 sky130_fd_sc_hd__nand2_1 _47378_ (.A(\delay_line[27][3] ),
    .B(net333),
    .Y(_18493_));
 sky130_fd_sc_hd__nand3b_2 _47379_ (.A_N(_18492_),
    .B(_18493_),
    .C(_16075_),
    .Y(_18494_));
 sky130_fd_sc_hd__and2_1 _47380_ (.A(\delay_line[27][3] ),
    .B(net333),
    .X(_18495_));
 sky130_fd_sc_hd__nand2_1 _47381_ (.A(\delay_line[27][2] ),
    .B(_16042_),
    .Y(_18496_));
 sky130_fd_sc_hd__o21ai_1 _47382_ (.A1(_18492_),
    .A2(_18495_),
    .B1(_18496_),
    .Y(_18497_));
 sky130_fd_sc_hd__nand2_1 _47383_ (.A(_18494_),
    .B(_18497_),
    .Y(_18498_));
 sky130_fd_sc_hd__clkbuf_2 _47384_ (.A(_18498_),
    .X(_18499_));
 sky130_fd_sc_hd__nor2_1 _47385_ (.A(_18491_),
    .B(_16086_),
    .Y(_18500_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47386_ (.A(_18500_),
    .X(_18501_));
 sky130_fd_sc_hd__a21o_1 _47387_ (.A1(_16108_),
    .A2(_18499_),
    .B1(_18501_),
    .X(_18502_));
 sky130_fd_sc_hd__o21ai_1 _47388_ (.A1(_16053_),
    .A2(_06579_),
    .B1(_18502_),
    .Y(_18503_));
 sky130_fd_sc_hd__a2111o_1 _47389_ (.A1(_16108_),
    .A2(_18499_),
    .B1(_18501_),
    .C1(_16053_),
    .D1(_06579_),
    .X(_18504_));
 sky130_fd_sc_hd__a2bb2oi_1 _47390_ (.A1_N(_18487_),
    .A2_N(_18490_),
    .B1(_18503_),
    .B2(_18504_),
    .Y(_18505_));
 sky130_fd_sc_hd__inv_2 _47391_ (.A(_18505_),
    .Y(_18506_));
 sky130_fd_sc_hd__or4bb_4 _47392_ (.A(_18487_),
    .B(_18490_),
    .C_N(_18503_),
    .D_N(_18504_),
    .X(_18507_));
 sky130_fd_sc_hd__inv_2 _47393_ (.A(net327),
    .Y(_18508_));
 sky130_fd_sc_hd__and3_1 _47394_ (.A(_18508_),
    .B(net328),
    .C(\delay_line[28][2] ),
    .X(_18509_));
 sky130_fd_sc_hd__buf_1 _47395_ (.A(\delay_line[28][5] ),
    .X(_18510_));
 sky130_fd_sc_hd__nand3b_1 _47396_ (.A_N(_18510_),
    .B(net328),
    .C(_15965_),
    .Y(_18511_));
 sky130_fd_sc_hd__nor2_1 _47397_ (.A(net327),
    .B(_18510_),
    .Y(_18512_));
 sky130_fd_sc_hd__and2_1 _47398_ (.A(net327),
    .B(\delay_line[28][5] ),
    .X(_18513_));
 sky130_fd_sc_hd__o2bb2ai_1 _47399_ (.A1_N(_15965_),
    .A2_N(net328),
    .B1(_18512_),
    .B2(_18513_),
    .Y(_18514_));
 sky130_fd_sc_hd__and3b_1 _47400_ (.A_N(\delay_line[28][0] ),
    .B(_18511_),
    .C(_18514_),
    .X(_18515_));
 sky130_fd_sc_hd__a21boi_1 _47401_ (.A1(_18511_),
    .A2(_18514_),
    .B1_N(_22248_),
    .Y(_18516_));
 sky130_fd_sc_hd__nor3_1 _47402_ (.A(_18509_),
    .B(_18515_),
    .C(_18516_),
    .Y(_18517_));
 sky130_fd_sc_hd__o21ai_1 _47403_ (.A1(_18515_),
    .A2(_18516_),
    .B1(_18509_),
    .Y(_18518_));
 sky130_fd_sc_hd__buf_1 _47404_ (.A(_18518_),
    .X(_18519_));
 sky130_fd_sc_hd__or4b_4 _47405_ (.A(_15976_),
    .B(_15954_),
    .C(_18517_),
    .D_N(_18519_),
    .X(_18520_));
 sky130_fd_sc_hd__inv_2 _47406_ (.A(_18517_),
    .Y(_18521_));
 sky130_fd_sc_hd__nand3_1 _47407_ (.A(_18521_),
    .B(_15932_),
    .C(_15965_),
    .Y(_18522_));
 sky130_fd_sc_hd__a22o_1 _47408_ (.A1(_15976_),
    .A2(_15932_),
    .B1(_18521_),
    .B2(_18519_),
    .X(_18523_));
 sky130_fd_sc_hd__a2bb2o_2 _47409_ (.A1_N(_15976_),
    .A2_N(_15954_),
    .B1(_18522_),
    .B2(_18523_),
    .X(_18524_));
 sky130_fd_sc_hd__a22o_2 _47410_ (.A1(_18506_),
    .A2(_18507_),
    .B1(_18520_),
    .B2(_18524_),
    .X(_18525_));
 sky130_fd_sc_hd__nand4_4 _47411_ (.A(_18506_),
    .B(_18507_),
    .C(_18520_),
    .D(_18524_),
    .Y(_18526_));
 sky130_fd_sc_hd__a21o_2 _47412_ (.A1(_16031_),
    .A2(_16141_),
    .B1(_16184_),
    .X(_18527_));
 sky130_fd_sc_hd__a21oi_1 _47413_ (.A1(_18525_),
    .A2(_18526_),
    .B1(_18527_),
    .Y(_18528_));
 sky130_fd_sc_hd__and3_1 _47414_ (.A(_18527_),
    .B(_18525_),
    .C(_18526_),
    .X(_18529_));
 sky130_fd_sc_hd__nor4_1 _47415_ (.A(_18483_),
    .B(_18484_),
    .C(_18528_),
    .D(_18529_),
    .Y(_18530_));
 sky130_fd_sc_hd__o22a_1 _47416_ (.A1(_18483_),
    .A2(_18484_),
    .B1(_18528_),
    .B2(_18529_),
    .X(_18531_));
 sky130_fd_sc_hd__nor2_1 _47417_ (.A(_18530_),
    .B(_18531_),
    .Y(_18532_));
 sky130_fd_sc_hd__or3_1 _47418_ (.A(_17336_),
    .B(_17346_),
    .C(_18532_),
    .X(_18533_));
 sky130_fd_sc_hd__o21ai_1 _47419_ (.A1(_17336_),
    .A2(_17346_),
    .B1(_18532_),
    .Y(_18534_));
 sky130_fd_sc_hd__and2_1 _47420_ (.A(_18533_),
    .B(_18534_),
    .X(_18535_));
 sky130_fd_sc_hd__o31ai_2 _47421_ (.A1(_15899_),
    .A2(_15910_),
    .A3(_16228_),
    .B1(_16195_),
    .Y(_18536_));
 sky130_fd_sc_hd__xnor2_2 _47422_ (.A(_18535_),
    .B(net119),
    .Y(_18537_));
 sky130_fd_sc_hd__and3_1 _47423_ (.A(_18301_),
    .B(_17412_),
    .C(_18448_),
    .X(_18538_));
 sky130_fd_sc_hd__nor3_1 _47424_ (.A(_18449_),
    .B(_18537_),
    .C(_18538_),
    .Y(_18539_));
 sky130_fd_sc_hd__o21ai_1 _47425_ (.A1(_18538_),
    .A2(_18449_),
    .B1(_18537_),
    .Y(_18540_));
 sky130_fd_sc_hd__or2b_1 _47426_ (.A(_18539_),
    .B_N(_18540_),
    .X(_18541_));
 sky130_fd_sc_hd__and2b_1 _47427_ (.A_N(_18300_),
    .B(_18541_),
    .X(_18542_));
 sky130_fd_sc_hd__and2b_1 _47428_ (.A_N(_18541_),
    .B(_18300_),
    .X(_18543_));
 sky130_fd_sc_hd__nor2_1 _47429_ (.A(_18542_),
    .B(_18543_),
    .Y(_18544_));
 sky130_fd_sc_hd__buf_1 _47430_ (.A(\delay_line[36][2] ),
    .X(_18545_));
 sky130_fd_sc_hd__buf_1 _47431_ (.A(_18545_),
    .X(_18546_));
 sky130_fd_sc_hd__and2b_1 _47432_ (.A_N(_18546_),
    .B(\delay_line[36][0] ),
    .X(_18547_));
 sky130_fd_sc_hd__and2b_1 _47433_ (.A_N(_05931_),
    .B(_18546_),
    .X(_18548_));
 sky130_fd_sc_hd__inv_2 _47434_ (.A(_17597_),
    .Y(_18549_));
 sky130_fd_sc_hd__buf_1 _47435_ (.A(\delay_line[35][5] ),
    .X(_18550_));
 sky130_fd_sc_hd__a21oi_1 _47436_ (.A1(_18549_),
    .A2(_18550_),
    .B1(_05909_),
    .Y(_18551_));
 sky130_fd_sc_hd__buf_1 _47437_ (.A(\delay_line[35][4] ),
    .X(_18552_));
 sky130_fd_sc_hd__or2b_1 _47438_ (.A(_18550_),
    .B_N(_18552_),
    .X(_18553_));
 sky130_fd_sc_hd__buf_1 _47439_ (.A(\delay_line[35][5] ),
    .X(_18554_));
 sky130_fd_sc_hd__o21ai_2 _47440_ (.A1(_17597_),
    .A2(_18554_),
    .B1(_05799_),
    .Y(_18555_));
 sky130_fd_sc_hd__a21oi_1 _47441_ (.A1(_18552_),
    .A2(_18550_),
    .B1(_18555_),
    .Y(_18556_));
 sky130_fd_sc_hd__a21oi_2 _47442_ (.A1(_18551_),
    .A2(_18553_),
    .B1(_18556_),
    .Y(_18557_));
 sky130_fd_sc_hd__nand2_1 _47443_ (.A(_17619_),
    .B(_17630_),
    .Y(_18558_));
 sky130_fd_sc_hd__xnor2_1 _47444_ (.A(_18557_),
    .B(_18558_),
    .Y(_18559_));
 sky130_fd_sc_hd__nand2_1 _47445_ (.A(_05887_),
    .B(_17695_),
    .Y(_18560_));
 sky130_fd_sc_hd__and3b_1 _47446_ (.A_N(_18559_),
    .B(_18560_),
    .C(_17673_),
    .X(_18561_));
 sky130_fd_sc_hd__buf_1 _47447_ (.A(_18559_),
    .X(_18562_));
 sky130_fd_sc_hd__a21boi_2 _47448_ (.A1(_17673_),
    .A2(_18560_),
    .B1_N(_18562_),
    .Y(_18563_));
 sky130_fd_sc_hd__a211o_1 _47449_ (.A1(_17716_),
    .A2(_17695_),
    .B1(_18561_),
    .C1(_18563_),
    .X(_18564_));
 sky130_fd_sc_hd__o211ai_4 _47450_ (.A1(_18561_),
    .A2(_18563_),
    .B1(_17716_),
    .C1(_17695_),
    .Y(_18565_));
 sky130_fd_sc_hd__o211a_1 _47451_ (.A1(_18547_),
    .A2(_18548_),
    .B1(_18564_),
    .C1(_18565_),
    .X(_18566_));
 sky130_fd_sc_hd__a211oi_1 _47452_ (.A1(_18564_),
    .A2(_18565_),
    .B1(_18547_),
    .C1(_18548_),
    .Y(_18567_));
 sky130_fd_sc_hd__nor2_1 _47453_ (.A(_18566_),
    .B(_18567_),
    .Y(_18568_));
 sky130_fd_sc_hd__and2b_1 _47454_ (.A_N(_05986_),
    .B(\delay_line[37][5] ),
    .X(_18569_));
 sky130_fd_sc_hd__buf_1 _47455_ (.A(\delay_line[37][5] ),
    .X(_18570_));
 sky130_fd_sc_hd__and2b_1 _47456_ (.A_N(_18570_),
    .B(_05986_),
    .X(_18571_));
 sky130_fd_sc_hd__nor2_1 _47457_ (.A(_18569_),
    .B(_18571_),
    .Y(_18572_));
 sky130_fd_sc_hd__and2b_1 _47458_ (.A_N(\delay_line[37][1] ),
    .B(_05986_),
    .X(_18573_));
 sky130_fd_sc_hd__a21oi_1 _47459_ (.A1(_18573_),
    .A2(_17543_),
    .B1(_17521_),
    .Y(_18574_));
 sky130_fd_sc_hd__xnor2_1 _47460_ (.A(_18572_),
    .B(_18574_),
    .Y(_18575_));
 sky130_fd_sc_hd__buf_1 _47461_ (.A(\delay_line[37][4] ),
    .X(_18576_));
 sky130_fd_sc_hd__a41oi_1 _47462_ (.A1(_04294_),
    .A2(_18576_),
    .A3(_05975_),
    .A4(_06008_),
    .B1(_17586_),
    .Y(_18577_));
 sky130_fd_sc_hd__or2b_1 _47463_ (.A(_18575_),
    .B_N(_18577_),
    .X(_18578_));
 sky130_fd_sc_hd__or2b_1 _47464_ (.A(_18577_),
    .B_N(_18575_),
    .X(_18579_));
 sky130_fd_sc_hd__and3_1 _47465_ (.A(_18568_),
    .B(_18578_),
    .C(_18579_),
    .X(_18580_));
 sky130_fd_sc_hd__o2bb2a_1 _47466_ (.A1_N(_18579_),
    .A2_N(_18578_),
    .B1(_18566_),
    .B2(_18567_),
    .X(_18581_));
 sky130_fd_sc_hd__o211a_1 _47467_ (.A1(_18580_),
    .A2(_18581_),
    .B1(_17748_),
    .C1(_17765_),
    .X(_18582_));
 sky130_fd_sc_hd__a211oi_2 _47468_ (.A1(_17748_),
    .A2(_17765_),
    .B1(_18580_),
    .C1(_18581_),
    .Y(_18583_));
 sky130_fd_sc_hd__nor2_1 _47469_ (.A(_18582_),
    .B(_18583_),
    .Y(_18584_));
 sky130_fd_sc_hd__inv_2 _47470_ (.A(\delay_line[40][5] ),
    .Y(_18585_));
 sky130_fd_sc_hd__or3b_1 _47471_ (.A(\delay_line[40][3] ),
    .B(_18585_),
    .C_N(_17769_),
    .X(_18586_));
 sky130_fd_sc_hd__or2_1 _47472_ (.A(\delay_line[40][5] ),
    .B(_17772_),
    .X(_18587_));
 sky130_fd_sc_hd__nand3_1 _47473_ (.A(_18586_),
    .B(_24776_),
    .C(_18587_),
    .Y(_18588_));
 sky130_fd_sc_hd__a21o_1 _47474_ (.A1(_18587_),
    .A2(_18586_),
    .B1(\delay_line[40][1] ),
    .X(_18589_));
 sky130_fd_sc_hd__and2b_1 _47475_ (.A_N(_17773_),
    .B(_22776_),
    .X(_18590_));
 sky130_fd_sc_hd__a211o_1 _47476_ (.A1(_18588_),
    .A2(_18589_),
    .B1(_17770_),
    .C1(_18590_),
    .X(_18591_));
 sky130_fd_sc_hd__o211ai_2 _47477_ (.A1(_17770_),
    .A2(_18590_),
    .B1(_18588_),
    .C1(_18589_),
    .Y(_18592_));
 sky130_fd_sc_hd__o2111a_1 _47478_ (.A1(_17774_),
    .A2(_17775_),
    .B1(_05722_),
    .C1(_05700_),
    .D1(_05711_),
    .X(_18593_));
 sky130_fd_sc_hd__and3_1 _47479_ (.A(_18591_),
    .B(_18592_),
    .C(_18593_),
    .X(_18594_));
 sky130_fd_sc_hd__a21oi_1 _47480_ (.A1(_18591_),
    .A2(_18592_),
    .B1(_18593_),
    .Y(_18595_));
 sky130_fd_sc_hd__and2_1 _47481_ (.A(net290),
    .B(\delay_line[38][5] ),
    .X(_18596_));
 sky130_fd_sc_hd__nor2_1 _47482_ (.A(net290),
    .B(\delay_line[38][5] ),
    .Y(_18597_));
 sky130_fd_sc_hd__nor2_1 _47483_ (.A(_18596_),
    .B(_18597_),
    .Y(_18598_));
 sky130_fd_sc_hd__buf_1 _47484_ (.A(_18598_),
    .X(_18599_));
 sky130_fd_sc_hd__o21ai_1 _47485_ (.A1(_17780_),
    .A2(_17781_),
    .B1(_18599_),
    .Y(_18600_));
 sky130_fd_sc_hd__or3_1 _47486_ (.A(_17780_),
    .B(_17781_),
    .C(_18599_),
    .X(_18601_));
 sky130_fd_sc_hd__nand2_1 _47487_ (.A(_17784_),
    .B(_17798_),
    .Y(_18602_));
 sky130_fd_sc_hd__clkbuf_2 _47488_ (.A(\delay_line[39][4] ),
    .X(_18603_));
 sky130_fd_sc_hd__o21a_1 _47489_ (.A1(_18603_),
    .A2(_05601_),
    .B1(_04118_),
    .X(_18604_));
 sky130_fd_sc_hd__nor2_1 _47490_ (.A(_17788_),
    .B(\delay_line[39][5] ),
    .Y(_18605_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47491_ (.A(\delay_line[39][5] ),
    .X(_18606_));
 sky130_fd_sc_hd__nand2_1 _47492_ (.A(_17788_),
    .B(_18606_),
    .Y(_18607_));
 sky130_fd_sc_hd__nand3b_1 _47493_ (.A_N(_18605_),
    .B(_18607_),
    .C(_05612_),
    .Y(_18608_));
 sky130_fd_sc_hd__and2_1 _47494_ (.A(_17788_),
    .B(\delay_line[39][5] ),
    .X(_18609_));
 sky130_fd_sc_hd__o21bai_1 _47495_ (.A1(_18605_),
    .A2(_18609_),
    .B1_N(_05612_),
    .Y(_18610_));
 sky130_fd_sc_hd__o211a_1 _47496_ (.A1(_17787_),
    .A2(_18604_),
    .B1(_18608_),
    .C1(_18610_),
    .X(_18611_));
 sky130_fd_sc_hd__a221oi_2 _47497_ (.A1(_18603_),
    .A2(_05612_),
    .B1(_18608_),
    .B2(_18610_),
    .C1(_18604_),
    .Y(_18612_));
 sky130_fd_sc_hd__or3b_2 _47498_ (.A(_18611_),
    .B(_18612_),
    .C_N(_04118_),
    .X(_18613_));
 sky130_fd_sc_hd__o21bai_2 _47499_ (.A1(_18611_),
    .A2(_18612_),
    .B1_N(_04129_),
    .Y(_18614_));
 sky130_fd_sc_hd__o31a_1 _47500_ (.A1(_04118_),
    .A2(_18603_),
    .A3(_05623_),
    .B1(_00392_),
    .X(_18615_));
 sky130_fd_sc_hd__a211o_1 _47501_ (.A1(_18613_),
    .A2(_18614_),
    .B1(_17795_),
    .C1(_18615_),
    .X(_18616_));
 sky130_fd_sc_hd__o211ai_4 _47502_ (.A1(_17795_),
    .A2(_18615_),
    .B1(_18613_),
    .C1(_18614_),
    .Y(_18617_));
 sky130_fd_sc_hd__o31a_1 _47503_ (.A1(_00403_),
    .A2(_04129_),
    .A3(_05634_),
    .B1(_17785_),
    .X(_18618_));
 sky130_fd_sc_hd__nand4_4 _47504_ (.A(_18602_),
    .B(_18616_),
    .C(_18617_),
    .D(_18618_),
    .Y(_18619_));
 sky130_fd_sc_hd__a22o_1 _47505_ (.A1(_18616_),
    .A2(_18617_),
    .B1(_18602_),
    .B2(_18618_),
    .X(_18620_));
 sky130_fd_sc_hd__and4_2 _47506_ (.A(_18600_),
    .B(_18601_),
    .C(_18619_),
    .D(_18620_),
    .X(_18621_));
 sky130_fd_sc_hd__a22oi_1 _47507_ (.A1(_18600_),
    .A2(_18601_),
    .B1(_18619_),
    .B2(_18620_),
    .Y(_18622_));
 sky130_fd_sc_hd__o22ai_1 _47508_ (.A1(_18594_),
    .A2(_18595_),
    .B1(_18621_),
    .B2(_18622_),
    .Y(_18623_));
 sky130_fd_sc_hd__or4_1 _47509_ (.A(_18594_),
    .B(_18595_),
    .C(_18621_),
    .D(_18622_),
    .X(_18624_));
 sky130_fd_sc_hd__and3_1 _47510_ (.A(_18584_),
    .B(_18623_),
    .C(_18624_),
    .X(_18625_));
 sky130_fd_sc_hd__a21oi_1 _47511_ (.A1(_18624_),
    .A2(_18623_),
    .B1(_18584_),
    .Y(_18626_));
 sky130_fd_sc_hd__nor2_4 _47512_ (.A(_18625_),
    .B(_18626_),
    .Y(_18627_));
 sky130_fd_sc_hd__o21bai_1 _47513_ (.A1(_17855_),
    .A2(_17852_),
    .B1_N(_17853_),
    .Y(_18628_));
 sky130_fd_sc_hd__or2_4 _47514_ (.A(_15657_),
    .B(_15910_),
    .X(_18629_));
 sky130_fd_sc_hd__buf_1 _47515_ (.A(\delay_line[34][3] ),
    .X(_18630_));
 sky130_fd_sc_hd__buf_1 _47516_ (.A(\delay_line[34][5] ),
    .X(_18631_));
 sky130_fd_sc_hd__and2_1 _47517_ (.A(_18630_),
    .B(_18631_),
    .X(_18632_));
 sky130_fd_sc_hd__clkbuf_2 _47518_ (.A(\delay_line[34][5] ),
    .X(_18633_));
 sky130_fd_sc_hd__nor2_1 _47519_ (.A(_18630_),
    .B(_18633_),
    .Y(_18634_));
 sky130_fd_sc_hd__o21ai_1 _47520_ (.A1(_18632_),
    .A2(_18634_),
    .B1(_17811_),
    .Y(_18635_));
 sky130_fd_sc_hd__nor2_1 _47521_ (.A(net308),
    .B(_02238_),
    .Y(_18636_));
 sky130_fd_sc_hd__and2_1 _47522_ (.A(net308),
    .B(\delay_line[34][2] ),
    .X(_18637_));
 sky130_fd_sc_hd__nor2_1 _47523_ (.A(_18636_),
    .B(_18637_),
    .Y(_18638_));
 sky130_fd_sc_hd__nand2_1 _47524_ (.A(_05392_),
    .B(_18633_),
    .Y(_18639_));
 sky130_fd_sc_hd__nand3b_2 _47525_ (.A_N(_18634_),
    .B(_17814_),
    .C(_18639_),
    .Y(_18640_));
 sky130_fd_sc_hd__nand3_2 _47526_ (.A(_18635_),
    .B(_18638_),
    .C(_18640_),
    .Y(_18641_));
 sky130_fd_sc_hd__a2bb2o_1 _47527_ (.A1_N(_18636_),
    .A2_N(_18637_),
    .B1(_18640_),
    .B2(_18635_),
    .X(_18642_));
 sky130_fd_sc_hd__a22o_1 _47528_ (.A1(_17811_),
    .A2(_17813_),
    .B1(_17816_),
    .B2(_17809_),
    .X(_18643_));
 sky130_fd_sc_hd__a21o_1 _47529_ (.A1(_18641_),
    .A2(_18642_),
    .B1(_18643_),
    .X(_18644_));
 sky130_fd_sc_hd__nand3_2 _47530_ (.A(_18643_),
    .B(_18641_),
    .C(_18642_),
    .Y(_18645_));
 sky130_fd_sc_hd__a22o_1 _47531_ (.A1(_22611_),
    .A2(_00612_),
    .B1(_18644_),
    .B2(_18645_),
    .X(_18646_));
 sky130_fd_sc_hd__nand4_2 _47532_ (.A(_18644_),
    .B(_18645_),
    .C(_22611_),
    .D(_00612_),
    .Y(_18647_));
 sky130_fd_sc_hd__and3_1 _47533_ (.A(_17819_),
    .B(_18646_),
    .C(_18647_),
    .X(_18648_));
 sky130_fd_sc_hd__a21oi_1 _47534_ (.A1(_18646_),
    .A2(_18647_),
    .B1(_17819_),
    .Y(_18649_));
 sky130_fd_sc_hd__inv_2 _47535_ (.A(net312),
    .Y(_18650_));
 sky130_fd_sc_hd__clkbuf_2 _47536_ (.A(_18650_),
    .X(_18651_));
 sky130_fd_sc_hd__buf_1 _47537_ (.A(\delay_line[33][1] ),
    .X(_18652_));
 sky130_fd_sc_hd__nand2b_1 _47538_ (.A_N(_18652_),
    .B(net315),
    .Y(_18653_));
 sky130_fd_sc_hd__or2b_1 _47539_ (.A(net315),
    .B_N(_18652_),
    .X(_18654_));
 sky130_fd_sc_hd__and3_1 _47540_ (.A(_18651_),
    .B(_18653_),
    .C(_18654_),
    .X(_18655_));
 sky130_fd_sc_hd__a21oi_1 _47541_ (.A1(_18653_),
    .A2(_18654_),
    .B1(_18650_),
    .Y(_18656_));
 sky130_fd_sc_hd__and4bb_1 _47542_ (.A_N(_18655_),
    .B_N(_18656_),
    .C(net315),
    .D(_17824_),
    .X(_18657_));
 sky130_fd_sc_hd__o2bb2a_1 _47543_ (.A1_N(_22534_),
    .A2_N(_17825_),
    .B1(_18655_),
    .B2(_18656_),
    .X(_18658_));
 sky130_fd_sc_hd__clkbuf_2 _47544_ (.A(_17831_),
    .X(_18659_));
 sky130_fd_sc_hd__clkbuf_2 _47545_ (.A(_18659_),
    .X(_18660_));
 sky130_fd_sc_hd__or4_1 _47546_ (.A(_24501_),
    .B(_24545_),
    .C(_05227_),
    .D(_05271_),
    .X(_18661_));
 sky130_fd_sc_hd__a21oi_1 _47547_ (.A1(_17831_),
    .A2(_05304_),
    .B1(_17833_),
    .Y(_18662_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47548_ (.A(\delay_line[32][5] ),
    .X(_18663_));
 sky130_fd_sc_hd__nor2_1 _47549_ (.A(_17832_),
    .B(_18663_),
    .Y(_18664_));
 sky130_fd_sc_hd__nand2_1 _47550_ (.A(_17832_),
    .B(_18663_),
    .Y(_18665_));
 sky130_fd_sc_hd__nand3b_2 _47551_ (.A_N(_18664_),
    .B(_18665_),
    .C(_05304_),
    .Y(_18666_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47552_ (.A(_18663_),
    .X(_18667_));
 sky130_fd_sc_hd__and2_1 _47553_ (.A(_17832_),
    .B(_18667_),
    .X(_18668_));
 sky130_fd_sc_hd__o21ai_2 _47554_ (.A1(_18664_),
    .A2(_18668_),
    .B1(_05249_),
    .Y(_18669_));
 sky130_fd_sc_hd__o211a_1 _47555_ (.A1(_17835_),
    .A2(_18662_),
    .B1(_18666_),
    .C1(_18669_),
    .X(_18670_));
 sky130_fd_sc_hd__inv_2 _47556_ (.A(\delay_line[32][4] ),
    .Y(_18671_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47557_ (.A(_18671_),
    .X(_18672_));
 sky130_fd_sc_hd__o21a_1 _47558_ (.A1(_18672_),
    .A2(_05238_),
    .B1(_17833_),
    .X(_18673_));
 sky130_fd_sc_hd__a21boi_2 _47559_ (.A1(_18666_),
    .A2(_18669_),
    .B1_N(_18673_),
    .Y(_18674_));
 sky130_fd_sc_hd__o21ai_1 _47560_ (.A1(_18670_),
    .A2(_18674_),
    .B1(_05227_),
    .Y(_18675_));
 sky130_fd_sc_hd__o211ai_2 _47561_ (.A1(_17835_),
    .A2(_18662_),
    .B1(_18666_),
    .C1(_18669_),
    .Y(_18676_));
 sky130_fd_sc_hd__nand3b_1 _47562_ (.A_N(_18674_),
    .B(_02106_),
    .C(_18676_),
    .Y(_18677_));
 sky130_fd_sc_hd__nand2_1 _47563_ (.A(_18675_),
    .B(_18677_),
    .Y(_18678_));
 sky130_fd_sc_hd__o21ba_1 _47564_ (.A1(_24534_),
    .A2(_17840_),
    .B1_N(_17841_),
    .X(_18679_));
 sky130_fd_sc_hd__nand2_1 _47565_ (.A(_18678_),
    .B(_18679_),
    .Y(_18680_));
 sky130_fd_sc_hd__nand3b_2 _47566_ (.A_N(_18679_),
    .B(_18675_),
    .C(_18677_),
    .Y(_18681_));
 sky130_fd_sc_hd__nand2_1 _47567_ (.A(_18680_),
    .B(_18681_),
    .Y(_18682_));
 sky130_fd_sc_hd__buf_1 _47568_ (.A(_18682_),
    .X(_18683_));
 sky130_fd_sc_hd__o221a_1 _47569_ (.A1(_18660_),
    .A2(_18661_),
    .B1(_17829_),
    .B2(_17844_),
    .C1(_18683_),
    .X(_18684_));
 sky130_fd_sc_hd__nand3b_1 _47570_ (.A_N(_17829_),
    .B(_17842_),
    .C(_17843_),
    .Y(_18685_));
 sky130_fd_sc_hd__or4b_1 _47571_ (.A(_05227_),
    .B(_18660_),
    .C(_05271_),
    .D_N(_24556_),
    .X(_18686_));
 sky130_fd_sc_hd__a21oi_1 _47572_ (.A1(_18685_),
    .A2(_18686_),
    .B1(_18683_),
    .Y(_18687_));
 sky130_fd_sc_hd__nor4_1 _47573_ (.A(_18657_),
    .B(_18658_),
    .C(_18684_),
    .D(_18687_),
    .Y(_18688_));
 sky130_fd_sc_hd__o22a_1 _47574_ (.A1(_18657_),
    .A2(_18658_),
    .B1(_18684_),
    .B2(_18687_),
    .X(_18689_));
 sky130_fd_sc_hd__o22a_1 _47575_ (.A1(_18648_),
    .A2(_18649_),
    .B1(_18688_),
    .B2(_18689_),
    .X(_18690_));
 sky130_fd_sc_hd__nor4_1 _47576_ (.A(_18648_),
    .B(_18649_),
    .C(net138),
    .D(_18689_),
    .Y(_18691_));
 sky130_fd_sc_hd__nor2_1 _47577_ (.A(_18690_),
    .B(_18691_),
    .Y(_18692_));
 sky130_fd_sc_hd__xnor2_1 _47578_ (.A(_18629_),
    .B(_18692_),
    .Y(_18693_));
 sky130_fd_sc_hd__and3_1 _47579_ (.A(_17847_),
    .B(_17850_),
    .C(_18693_),
    .X(_18694_));
 sky130_fd_sc_hd__a21oi_1 _47580_ (.A1(_17847_),
    .A2(_17850_),
    .B1(_18693_),
    .Y(_18695_));
 sky130_fd_sc_hd__nor2_1 _47581_ (.A(_18694_),
    .B(_18695_),
    .Y(_18696_));
 sky130_fd_sc_hd__or2_1 _47582_ (.A(_18628_),
    .B(_18696_),
    .X(_18697_));
 sky130_fd_sc_hd__nand2_1 _47583_ (.A(_18696_),
    .B(_18628_),
    .Y(_18698_));
 sky130_fd_sc_hd__and2_1 _47584_ (.A(_18697_),
    .B(_18698_),
    .X(_18699_));
 sky130_fd_sc_hd__xnor2_1 _47585_ (.A(_18627_),
    .B(_18699_),
    .Y(_18700_));
 sky130_fd_sc_hd__nand3_1 _47586_ (.A(_16261_),
    .B(_16305_),
    .C(_18700_),
    .Y(_18701_));
 sky130_fd_sc_hd__a21o_1 _47587_ (.A1(_16261_),
    .A2(_16305_),
    .B1(_18700_),
    .X(_18702_));
 sky130_fd_sc_hd__or2_1 _47588_ (.A(_17859_),
    .B(_17860_),
    .X(_18703_));
 sky130_fd_sc_hd__a21oi_1 _47589_ (.A1(_18701_),
    .A2(_18702_),
    .B1(_18703_),
    .Y(_18704_));
 sky130_fd_sc_hd__and3_1 _47590_ (.A(_18703_),
    .B(_18701_),
    .C(_18702_),
    .X(_18705_));
 sky130_fd_sc_hd__nor2_1 _47591_ (.A(_18704_),
    .B(_18705_),
    .Y(_18706_));
 sky130_fd_sc_hd__xnor2_1 _47592_ (.A(_18544_),
    .B(_18706_),
    .Y(_18707_));
 sky130_fd_sc_hd__or2b_1 _47593_ (.A(_17445_),
    .B_N(_17456_),
    .X(_18708_));
 sky130_fd_sc_hd__a21bo_1 _47594_ (.A1(_17467_),
    .A2(_17866_),
    .B1_N(_18708_),
    .X(_18709_));
 sky130_fd_sc_hd__and2b_1 _47595_ (.A_N(_18707_),
    .B(_18709_),
    .X(_18710_));
 sky130_fd_sc_hd__and2b_1 _47596_ (.A_N(_18709_),
    .B(_18707_),
    .X(_18711_));
 sky130_fd_sc_hd__or2_1 _47597_ (.A(_18710_),
    .B(_18711_),
    .X(_18712_));
 sky130_fd_sc_hd__o21ai_4 _47598_ (.A1(_18293_),
    .A2(_18299_),
    .B1(_18712_),
    .Y(_18713_));
 sky130_fd_sc_hd__a31oi_2 _47599_ (.A1(_18286_),
    .A2(_18291_),
    .A3(_18292_),
    .B1(_18712_),
    .Y(_18714_));
 sky130_fd_sc_hd__a21o_1 _47600_ (.A1(_18286_),
    .A2(_18291_),
    .B1(_18292_),
    .X(_18715_));
 sky130_fd_sc_hd__nand2_2 _47601_ (.A(_18714_),
    .B(_18715_),
    .Y(_18716_));
 sky130_fd_sc_hd__a31o_1 _47602_ (.A1(_17872_),
    .A2(_17874_),
    .A3(_17875_),
    .B1(_17868_),
    .X(_18717_));
 sky130_fd_sc_hd__a21oi_2 _47603_ (.A1(_18713_),
    .A2(_18716_),
    .B1(_18717_),
    .Y(_18718_));
 sky130_fd_sc_hd__a21oi_2 _47604_ (.A1(_15482_),
    .A2(_15537_),
    .B1(_17870_),
    .Y(_18719_));
 sky130_fd_sc_hd__o211a_1 _47605_ (.A1(_17868_),
    .A2(_18719_),
    .B1(_18713_),
    .C1(_18716_),
    .X(_18720_));
 sky130_fd_sc_hd__o21ai_1 _47606_ (.A1(_15526_),
    .A2(_15460_),
    .B1(_17873_),
    .Y(_18721_));
 sky130_fd_sc_hd__inv_2 _47607_ (.A(_11295_),
    .Y(_18722_));
 sky130_fd_sc_hd__o21ai_1 _47608_ (.A1(_10778_),
    .A2(_18722_),
    .B1(_11361_),
    .Y(_18723_));
 sky130_fd_sc_hd__and3_1 _47609_ (.A(_18722_),
    .B(_10811_),
    .C(_10778_),
    .X(_18724_));
 sky130_fd_sc_hd__nor2_1 _47610_ (.A(_11295_),
    .B(\delay_line[17][5] ),
    .Y(_18725_));
 sky130_fd_sc_hd__nand2_1 _47611_ (.A(\delay_line[17][4] ),
    .B(\delay_line[17][5] ),
    .Y(_18726_));
 sky130_fd_sc_hd__nor2b_2 _47612_ (.A(_18725_),
    .B_N(_18726_),
    .Y(_18727_));
 sky130_fd_sc_hd__and4_1 _47613_ (.A(_11328_),
    .B(_18727_),
    .C(_22183_),
    .D(_23622_),
    .X(_18728_));
 sky130_fd_sc_hd__buf_2 _47614_ (.A(_10932_),
    .X(_18729_));
 sky130_fd_sc_hd__o21ai_1 _47615_ (.A1(_23611_),
    .A2(_18729_),
    .B1(_22161_),
    .Y(_18730_));
 sky130_fd_sc_hd__a21o_1 _47616_ (.A1(_23611_),
    .A2(_18729_),
    .B1(_22172_),
    .X(_18731_));
 sky130_fd_sc_hd__a21oi_1 _47617_ (.A1(_18730_),
    .A2(_18731_),
    .B1(_18727_),
    .Y(_18732_));
 sky130_fd_sc_hd__and3_1 _47618_ (.A(_18727_),
    .B(_18730_),
    .C(_18731_),
    .X(_18733_));
 sky130_fd_sc_hd__o21a_1 _47619_ (.A1(_18732_),
    .A2(_18733_),
    .B1(_11317_),
    .X(_18734_));
 sky130_fd_sc_hd__nor4_1 _47620_ (.A(_18723_),
    .B(_18724_),
    .C(_18728_),
    .D(_18734_),
    .Y(_18735_));
 sky130_fd_sc_hd__o22a_1 _47621_ (.A1(_18723_),
    .A2(_18724_),
    .B1(_18728_),
    .B2(_18734_),
    .X(_18736_));
 sky130_fd_sc_hd__and2_1 _47622_ (.A(_11416_),
    .B(net366),
    .X(_18737_));
 sky130_fd_sc_hd__nor2_1 _47623_ (.A(_11416_),
    .B(net366),
    .Y(_18738_));
 sky130_fd_sc_hd__o2bb2a_1 _47624_ (.A1_N(_11042_),
    .A2_N(_11449_),
    .B1(_18737_),
    .B2(_18738_),
    .X(_18739_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47625_ (.A(net366),
    .X(_18740_));
 sky130_fd_sc_hd__and3b_1 _47626_ (.A_N(_18740_),
    .B(_11449_),
    .C(_11042_),
    .X(_18741_));
 sky130_fd_sc_hd__nor2_1 _47627_ (.A(_10899_),
    .B(_10921_),
    .Y(_18742_));
 sky130_fd_sc_hd__xnor2_1 _47628_ (.A(_23600_),
    .B(_18742_),
    .Y(_18743_));
 sky130_fd_sc_hd__clkbuf_2 _47629_ (.A(_18743_),
    .X(_18744_));
 sky130_fd_sc_hd__nor3_2 _47630_ (.A(_18739_),
    .B(_18741_),
    .C(_18744_),
    .Y(_18745_));
 sky130_fd_sc_hd__o21a_1 _47631_ (.A1(_18739_),
    .A2(_18741_),
    .B1(_18744_),
    .X(_18746_));
 sky130_fd_sc_hd__o2111ai_4 _47632_ (.A1(_10910_),
    .A2(_11438_),
    .B1(_11460_),
    .C1(_04865_),
    .D1(_04832_),
    .Y(_18747_));
 sky130_fd_sc_hd__o211ai_2 _47633_ (.A1(_18745_),
    .A2(_18746_),
    .B1(_11460_),
    .C1(_18747_),
    .Y(_18748_));
 sky130_fd_sc_hd__a211o_1 _47634_ (.A1(_11460_),
    .A2(_18747_),
    .B1(_18745_),
    .C1(_18746_),
    .X(_18749_));
 sky130_fd_sc_hd__nand2_2 _47635_ (.A(_18748_),
    .B(_18749_),
    .Y(_18750_));
 sky130_fd_sc_hd__xnor2_1 _47636_ (.A(_11504_),
    .B(_18750_),
    .Y(_18751_));
 sky130_fd_sc_hd__nor3b_2 _47637_ (.A(net210),
    .B(_18736_),
    .C_N(_18751_),
    .Y(_18752_));
 sky130_fd_sc_hd__o21ba_1 _47638_ (.A1(net210),
    .A2(_18736_),
    .B1_N(_18751_),
    .X(_18753_));
 sky130_fd_sc_hd__or2_2 _47639_ (.A(_18752_),
    .B(_18753_),
    .X(_18754_));
 sky130_fd_sc_hd__inv_2 _47640_ (.A(_18754_),
    .Y(_18755_));
 sky130_fd_sc_hd__nand2_1 _47641_ (.A(_18721_),
    .B(_18755_),
    .Y(_18756_));
 sky130_fd_sc_hd__o211ai_2 _47642_ (.A1(_15526_),
    .A2(_15460_),
    .B1(_17873_),
    .C1(_18754_),
    .Y(_18757_));
 sky130_fd_sc_hd__nand2_1 _47643_ (.A(_18756_),
    .B(_18757_),
    .Y(_18758_));
 sky130_fd_sc_hd__a2bb2o_1 _47644_ (.A1_N(_11625_),
    .A2_N(_11647_),
    .B1(_15449_),
    .B2(_15493_),
    .X(_18759_));
 sky130_fd_sc_hd__a21oi_1 _47645_ (.A1(_17873_),
    .A2(_18759_),
    .B1(_18754_),
    .Y(_18760_));
 sky130_fd_sc_hd__a31o_1 _47646_ (.A1(_17873_),
    .A2(_18759_),
    .A3(_18754_),
    .B1(_11537_),
    .X(_18761_));
 sky130_fd_sc_hd__o2bb2ai_2 _47647_ (.A1_N(_11537_),
    .A2_N(_18758_),
    .B1(_18760_),
    .B2(_18761_),
    .Y(_18762_));
 sky130_fd_sc_hd__o21bai_1 _47648_ (.A1(_18718_),
    .A2(_18720_),
    .B1_N(_18762_),
    .Y(_18763_));
 sky130_fd_sc_hd__o31a_1 _47649_ (.A1(_11592_),
    .A2(_11614_),
    .A3(_17879_),
    .B1(_17883_),
    .X(_18764_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47650_ (.A(_11394_),
    .X(_18765_));
 sky130_fd_sc_hd__o41a_1 _47651_ (.A1(_11383_),
    .A2(_18765_),
    .A3(_11504_),
    .A4(_11526_),
    .B1(_18758_),
    .X(_18766_));
 sky130_fd_sc_hd__inv_2 _47652_ (.A(_11537_),
    .Y(_18767_));
 sky130_fd_sc_hd__and3_1 _47653_ (.A(_18756_),
    .B(_18757_),
    .C(_18767_),
    .X(_18768_));
 sky130_fd_sc_hd__a21o_1 _47654_ (.A1(_18713_),
    .A2(_18716_),
    .B1(_18717_),
    .X(_18769_));
 sky130_fd_sc_hd__o211ai_4 _47655_ (.A1(_17868_),
    .A2(_18719_),
    .B1(_18713_),
    .C1(_18716_),
    .Y(_18770_));
 sky130_fd_sc_hd__o211ai_1 _47656_ (.A1(_18766_),
    .A2(_18768_),
    .B1(_18769_),
    .C1(_18770_),
    .Y(_18771_));
 sky130_fd_sc_hd__nand3_2 _47657_ (.A(_18763_),
    .B(_18764_),
    .C(_18771_),
    .Y(_18772_));
 sky130_fd_sc_hd__a21o_1 _47658_ (.A1(_17881_),
    .A2(_17882_),
    .B1(_17877_),
    .X(_18773_));
 sky130_fd_sc_hd__o21ai_2 _47659_ (.A1(_18718_),
    .A2(_18720_),
    .B1(_18762_),
    .Y(_18774_));
 sky130_fd_sc_hd__nand3b_2 _47660_ (.A_N(_18762_),
    .B(_18769_),
    .C(_18770_),
    .Y(_18775_));
 sky130_fd_sc_hd__nand3_1 _47661_ (.A(_18773_),
    .B(_18774_),
    .C(_18775_),
    .Y(_18776_));
 sky130_fd_sc_hd__or3b_1 _47662_ (.A(_10679_),
    .B(_18767_),
    .C_N(_11559_),
    .X(_18777_));
 sky130_fd_sc_hd__inv_2 _47663_ (.A(_18777_),
    .Y(_18778_));
 sky130_fd_sc_hd__clkbuf_2 _47664_ (.A(_11361_),
    .X(_18779_));
 sky130_fd_sc_hd__clkbuf_2 _47665_ (.A(_18779_),
    .X(_18780_));
 sky130_fd_sc_hd__o21ai_1 _47666_ (.A1(_18780_),
    .A2(_10866_),
    .B1(_22150_),
    .Y(_18781_));
 sky130_fd_sc_hd__or3_2 _47667_ (.A(_18779_),
    .B(_10866_),
    .C(_22150_),
    .X(_18782_));
 sky130_fd_sc_hd__a21oi_1 _47668_ (.A1(_18781_),
    .A2(_18782_),
    .B1(_18765_),
    .Y(_18783_));
 sky130_fd_sc_hd__a21oi_2 _47669_ (.A1(_05161_),
    .A2(_18765_),
    .B1(_18783_),
    .Y(_18784_));
 sky130_fd_sc_hd__o21a_1 _47670_ (.A1(_18778_),
    .A2(_11614_),
    .B1(_18784_),
    .X(_18785_));
 sky130_fd_sc_hd__a311oi_2 _47671_ (.A1(_10690_),
    .A2(_11537_),
    .A3(_11559_),
    .B1(_11614_),
    .C1(_18784_),
    .Y(_18786_));
 sky130_fd_sc_hd__o2bb2ai_1 _47672_ (.A1_N(_18772_),
    .A2_N(_18776_),
    .B1(_18785_),
    .B2(_18786_),
    .Y(_18787_));
 sky130_fd_sc_hd__nor2_1 _47673_ (.A(_18785_),
    .B(_18786_),
    .Y(_18788_));
 sky130_fd_sc_hd__nand3_1 _47674_ (.A(_18772_),
    .B(_18776_),
    .C(_18788_),
    .Y(_18789_));
 sky130_fd_sc_hd__o21a_1 _47675_ (.A1(_11273_),
    .A2(_17885_),
    .B1(_17886_),
    .X(_18790_));
 sky130_fd_sc_hd__a21boi_1 _47676_ (.A1(_18787_),
    .A2(_18789_),
    .B1_N(_18790_),
    .Y(_18791_));
 sky130_fd_sc_hd__nand3b_1 _47677_ (.A_N(_18790_),
    .B(_18787_),
    .C(_18789_),
    .Y(_18792_));
 sky130_fd_sc_hd__and2b_1 _47678_ (.A_N(_18791_),
    .B(_18792_),
    .X(_18793_));
 sky130_fd_sc_hd__xor2_1 _47679_ (.A(_11251_),
    .B(_18793_),
    .X(_18794_));
 sky130_fd_sc_hd__a21oi_2 _47680_ (.A1(_17890_),
    .A2(_17893_),
    .B1(_18794_),
    .Y(_18795_));
 sky130_fd_sc_hd__and3_1 _47681_ (.A(_18794_),
    .B(_17893_),
    .C(_17890_),
    .X(_18796_));
 sky130_fd_sc_hd__nor2_1 _47682_ (.A(_18795_),
    .B(_18796_),
    .Y(_00036_));
 sky130_fd_sc_hd__nand2_1 _47683_ (.A(_18286_),
    .B(_18292_),
    .Y(_18797_));
 sky130_fd_sc_hd__xnor2_1 _47684_ (.A(_10932_),
    .B(_11438_),
    .Y(_18798_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47685_ (.A(_18798_),
    .X(_18799_));
 sky130_fd_sc_hd__xor2_2 _47686_ (.A(net366),
    .B(net365),
    .X(_18800_));
 sky130_fd_sc_hd__nand2_1 _47687_ (.A(_18737_),
    .B(_18800_),
    .Y(_18801_));
 sky130_fd_sc_hd__a21o_1 _47688_ (.A1(_11449_),
    .A2(_18740_),
    .B1(_18800_),
    .X(_18802_));
 sky130_fd_sc_hd__nand3b_1 _47689_ (.A_N(_18799_),
    .B(_18801_),
    .C(_18802_),
    .Y(_18803_));
 sky130_fd_sc_hd__a21bo_1 _47690_ (.A1(_18802_),
    .A2(_18801_),
    .B1_N(_18799_),
    .X(_18804_));
 sky130_fd_sc_hd__and2_1 _47691_ (.A(_18803_),
    .B(_18804_),
    .X(_18805_));
 sky130_fd_sc_hd__or3_1 _47692_ (.A(_18741_),
    .B(_18745_),
    .C(_18805_),
    .X(_18806_));
 sky130_fd_sc_hd__o21ai_2 _47693_ (.A1(_18741_),
    .A2(_18745_),
    .B1(_18805_),
    .Y(_18807_));
 sky130_fd_sc_hd__nand2_2 _47694_ (.A(_18806_),
    .B(_18807_),
    .Y(_18808_));
 sky130_fd_sc_hd__o21ai_1 _47695_ (.A1(_11548_),
    .A2(_18750_),
    .B1(_18749_),
    .Y(_18809_));
 sky130_fd_sc_hd__xor2_1 _47696_ (.A(_18808_),
    .B(_18809_),
    .X(_18810_));
 sky130_fd_sc_hd__clkbuf_2 _47697_ (.A(\delay_line[17][5] ),
    .X(_18811_));
 sky130_fd_sc_hd__nor2_1 _47698_ (.A(_18811_),
    .B(\delay_line[17][6] ),
    .Y(_18812_));
 sky130_fd_sc_hd__and2_2 _47699_ (.A(\delay_line[17][5] ),
    .B(\delay_line[17][6] ),
    .X(_18813_));
 sky130_fd_sc_hd__a21oi_2 _47700_ (.A1(_23600_),
    .A2(_18742_),
    .B1(_10899_),
    .Y(_18814_));
 sky130_fd_sc_hd__or2b_1 _47701_ (.A(_18814_),
    .B_N(_11020_),
    .X(_18815_));
 sky130_fd_sc_hd__a211o_1 _47702_ (.A1(_23600_),
    .A2(_18742_),
    .B1(_10910_),
    .C1(_11009_),
    .X(_18816_));
 sky130_fd_sc_hd__a21bo_1 _47703_ (.A1(_18815_),
    .A2(_18816_),
    .B1_N(_18730_),
    .X(_18817_));
 sky130_fd_sc_hd__o2111ai_4 _47704_ (.A1(_23611_),
    .A2(_18729_),
    .B1(_18816_),
    .C1(_22172_),
    .D1(_18815_),
    .Y(_18818_));
 sky130_fd_sc_hd__or4bb_4 _47705_ (.A(_18812_),
    .B(_18813_),
    .C_N(_18817_),
    .D_N(_18818_),
    .X(_18819_));
 sky130_fd_sc_hd__a2bb2o_1 _47706_ (.A1_N(_18812_),
    .A2_N(_18813_),
    .B1(_18817_),
    .B2(_18818_),
    .X(_18820_));
 sky130_fd_sc_hd__and3_1 _47707_ (.A(_18819_),
    .B(_18820_),
    .C(_18733_),
    .X(_18821_));
 sky130_fd_sc_hd__a21oi_1 _47708_ (.A1(_18819_),
    .A2(_18820_),
    .B1(_18733_),
    .Y(_18822_));
 sky130_fd_sc_hd__nor2_2 _47709_ (.A(_18811_),
    .B(_18722_),
    .Y(_18823_));
 sky130_fd_sc_hd__nand2_2 _47710_ (.A(_11295_),
    .B(_10811_),
    .Y(_18824_));
 sky130_fd_sc_hd__mux2_1 _47711_ (.A0(_18811_),
    .A1(_18823_),
    .S(_18824_),
    .X(_18825_));
 sky130_fd_sc_hd__nor3b_1 _47712_ (.A(_18821_),
    .B(_18822_),
    .C_N(_18825_),
    .Y(_18826_));
 sky130_fd_sc_hd__o21ba_1 _47713_ (.A1(_18821_),
    .A2(_18822_),
    .B1_N(_18825_),
    .X(_18827_));
 sky130_fd_sc_hd__or2_1 _47714_ (.A(_18826_),
    .B(_18827_),
    .X(_18828_));
 sky130_fd_sc_hd__xnor2_1 _47715_ (.A(_18810_),
    .B(_18828_),
    .Y(_18829_));
 sky130_fd_sc_hd__a21oi_1 _47716_ (.A1(_18291_),
    .A2(_18797_),
    .B1(_18829_),
    .Y(_18830_));
 sky130_fd_sc_hd__nand3_1 _47717_ (.A(_18291_),
    .B(_18797_),
    .C(_18829_),
    .Y(_18831_));
 sky130_fd_sc_hd__nand2b_1 _47718_ (.A_N(_18830_),
    .B(_18831_),
    .Y(_18832_));
 sky130_fd_sc_hd__xor2_1 _47719_ (.A(_18752_),
    .B(_18832_),
    .X(_18833_));
 sky130_fd_sc_hd__inv_2 _47720_ (.A(_18833_),
    .Y(_18834_));
 sky130_fd_sc_hd__a21o_1 _47721_ (.A1(_18714_),
    .A2(_18715_),
    .B1(_18710_),
    .X(_18835_));
 sky130_fd_sc_hd__buf_2 _47722_ (.A(\delay_line[23][5] ),
    .X(_18836_));
 sky130_fd_sc_hd__o221a_1 _47723_ (.A1(_18259_),
    .A2(_18836_),
    .B1(_17906_),
    .B2(_18236_),
    .C1(_18239_),
    .X(_18837_));
 sky130_fd_sc_hd__inv_2 _47724_ (.A(_18624_),
    .Y(_18838_));
 sky130_fd_sc_hd__a22o_1 _47725_ (.A1(_18232_),
    .A2(_18231_),
    .B1(_18230_),
    .B2(_18229_),
    .X(_18839_));
 sky130_fd_sc_hd__nor2_2 _47726_ (.A(_18213_),
    .B(_18206_),
    .Y(_18840_));
 sky130_fd_sc_hd__o211a_1 _47727_ (.A1(_18152_),
    .A2(_18153_),
    .B1(_18154_),
    .C1(_18156_),
    .X(_18841_));
 sky130_fd_sc_hd__a2bb2o_1 _47728_ (.A1_N(_02865_),
    .A2_N(_18065_),
    .B1(_18066_),
    .B2(_18049_),
    .X(_18842_));
 sky130_fd_sc_hd__xor2_1 _47729_ (.A(_22996_),
    .B(_18036_),
    .X(_18843_));
 sky130_fd_sc_hd__buf_2 _47730_ (.A(_08976_),
    .X(_18844_));
 sky130_fd_sc_hd__buf_1 _47731_ (.A(\delay_line[8][6] ),
    .X(_18845_));
 sky130_fd_sc_hd__o21a_1 _47732_ (.A1(_18039_),
    .A2(_18845_),
    .B1(_18030_),
    .X(_18846_));
 sky130_fd_sc_hd__nand2_1 _47733_ (.A(_18039_),
    .B(_18845_),
    .Y(_18847_));
 sky130_fd_sc_hd__nand2_1 _47734_ (.A(_18846_),
    .B(_18847_),
    .Y(_18848_));
 sky130_fd_sc_hd__and2_1 _47735_ (.A(\delay_line[8][5] ),
    .B(\delay_line[8][6] ),
    .X(_18849_));
 sky130_fd_sc_hd__nor2_1 _47736_ (.A(_18039_),
    .B(_18845_),
    .Y(_18850_));
 sky130_fd_sc_hd__o21ai_2 _47737_ (.A1(_18849_),
    .A2(_18850_),
    .B1(_11811_),
    .Y(_18851_));
 sky130_fd_sc_hd__a22o_1 _47738_ (.A1(_18031_),
    .A2(_18033_),
    .B1(_18848_),
    .B2(_18851_),
    .X(_18852_));
 sky130_fd_sc_hd__o2111ai_1 _47739_ (.A1(_08976_),
    .A2(_11822_),
    .B1(_18033_),
    .C1(_18848_),
    .D1(_18851_),
    .Y(_18853_));
 sky130_fd_sc_hd__nand3_2 _47740_ (.A(_18844_),
    .B(_18852_),
    .C(_18853_),
    .Y(_18854_));
 sky130_fd_sc_hd__o21ai_1 _47741_ (.A1(_08976_),
    .A2(_11811_),
    .B1(_18032_),
    .Y(_18855_));
 sky130_fd_sc_hd__a21o_1 _47742_ (.A1(_18848_),
    .A2(_18851_),
    .B1(_18855_),
    .X(_18856_));
 sky130_fd_sc_hd__nand3_1 _47743_ (.A(_18855_),
    .B(_18848_),
    .C(_18851_),
    .Y(_18857_));
 sky130_fd_sc_hd__nand3_2 _47744_ (.A(_18856_),
    .B(_09020_),
    .C(_18857_),
    .Y(_18858_));
 sky130_fd_sc_hd__nand3_2 _47745_ (.A(_18854_),
    .B(_23084_),
    .C(_18858_),
    .Y(_18859_));
 sky130_fd_sc_hd__a21o_1 _47746_ (.A1(_18858_),
    .A2(_18854_),
    .B1(_23073_),
    .X(_18860_));
 sky130_fd_sc_hd__nand3b_2 _47747_ (.A_N(_18041_),
    .B(_18859_),
    .C(_18860_),
    .Y(_18861_));
 sky130_fd_sc_hd__nand2_1 _47748_ (.A(_18859_),
    .B(_18860_),
    .Y(_18862_));
 sky130_fd_sc_hd__nand2_1 _47749_ (.A(_18042_),
    .B(_18862_),
    .Y(_18863_));
 sky130_fd_sc_hd__nand3b_2 _47750_ (.A_N(_18843_),
    .B(_18861_),
    .C(_18863_),
    .Y(_18864_));
 sky130_fd_sc_hd__a21bo_1 _47751_ (.A1(_18861_),
    .A2(_18863_),
    .B1_N(_18843_),
    .X(_18865_));
 sky130_fd_sc_hd__o311a_1 _47752_ (.A1(_13009_),
    .A2(_18057_),
    .A3(_18059_),
    .B1(_02865_),
    .C1(_08668_),
    .X(_18866_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47753_ (.A(net421),
    .X(_18867_));
 sky130_fd_sc_hd__nor2_1 _47754_ (.A(_17912_),
    .B(_18867_),
    .Y(_18868_));
 sky130_fd_sc_hd__buf_1 _47755_ (.A(_18868_),
    .X(_18869_));
 sky130_fd_sc_hd__and2_1 _47756_ (.A(_17912_),
    .B(_18867_),
    .X(_18870_));
 sky130_fd_sc_hd__nand3b_1 _47757_ (.A_N(\delay_line[9][4] ),
    .B(net422),
    .C(_02843_),
    .Y(_18871_));
 sky130_fd_sc_hd__or2b_1 _47758_ (.A(net422),
    .B_N(_12976_),
    .X(_18872_));
 sky130_fd_sc_hd__o211ai_1 _47759_ (.A1(_18869_),
    .A2(_18870_),
    .B1(_18871_),
    .C1(_18872_),
    .Y(_18873_));
 sky130_fd_sc_hd__a211o_1 _47760_ (.A1(_18872_),
    .A2(_18871_),
    .B1(_18870_),
    .C1(_18868_),
    .X(_18874_));
 sky130_fd_sc_hd__a21oi_1 _47761_ (.A1(_18873_),
    .A2(_18874_),
    .B1(_17914_),
    .Y(_18875_));
 sky130_fd_sc_hd__nand4b_1 _47762_ (.A_N(_18053_),
    .B(_12987_),
    .C(_02854_),
    .D(_25073_),
    .Y(_18876_));
 sky130_fd_sc_hd__and3_1 _47763_ (.A(_18874_),
    .B(_17914_),
    .C(_18873_),
    .X(_18877_));
 sky130_fd_sc_hd__nor3_1 _47764_ (.A(_18875_),
    .B(_18876_),
    .C(_18877_),
    .Y(_18878_));
 sky130_fd_sc_hd__o21ai_1 _47765_ (.A1(_18877_),
    .A2(_18875_),
    .B1(_18876_),
    .Y(_18879_));
 sky130_fd_sc_hd__and2b_1 _47766_ (.A_N(_18878_),
    .B(_18879_),
    .X(_18880_));
 sky130_fd_sc_hd__nor3_1 _47767_ (.A(_18061_),
    .B(_18866_),
    .C(_18880_),
    .Y(_18881_));
 sky130_fd_sc_hd__o21a_1 _47768_ (.A1(_18061_),
    .A2(_18866_),
    .B1(_18880_),
    .X(_18882_));
 sky130_fd_sc_hd__nor2_1 _47769_ (.A(_18881_),
    .B(_18882_),
    .Y(_18883_));
 sky130_fd_sc_hd__a21oi_1 _47770_ (.A1(_18864_),
    .A2(_18865_),
    .B1(_18883_),
    .Y(_18884_));
 sky130_fd_sc_hd__or4b_1 _47771_ (.A(_13053_),
    .B(_13064_),
    .C(_17931_),
    .D_N(_13020_),
    .X(_18885_));
 sky130_fd_sc_hd__nand3_1 _47772_ (.A(_18883_),
    .B(_18864_),
    .C(_18865_),
    .Y(_18886_));
 sky130_fd_sc_hd__inv_2 _47773_ (.A(_18886_),
    .Y(_18887_));
 sky130_fd_sc_hd__or3_1 _47774_ (.A(_18884_),
    .B(_18885_),
    .C(_18887_),
    .X(_18888_));
 sky130_fd_sc_hd__o21ai_1 _47775_ (.A1(_18887_),
    .A2(_18884_),
    .B1(_18885_),
    .Y(_18889_));
 sky130_fd_sc_hd__and3_1 _47776_ (.A(_18842_),
    .B(_18888_),
    .C(_18889_),
    .X(_18890_));
 sky130_fd_sc_hd__a21oi_1 _47777_ (.A1(_18888_),
    .A2(_18889_),
    .B1(_18842_),
    .Y(_18891_));
 sky130_fd_sc_hd__nor2_1 _47778_ (.A(_18890_),
    .B(_18891_),
    .Y(_18892_));
 sky130_fd_sc_hd__nor2_1 _47779_ (.A(_17930_),
    .B(_17932_),
    .Y(_18893_));
 sky130_fd_sc_hd__a31oi_2 _47780_ (.A1(_18001_),
    .A2(_18002_),
    .A3(_18007_),
    .B1(_18893_),
    .Y(_18894_));
 sky130_fd_sc_hd__or3_1 _47781_ (.A(_25303_),
    .B(_17997_),
    .C(_18003_),
    .X(_18895_));
 sky130_fd_sc_hd__o21ai_2 _47782_ (.A1(_17997_),
    .A2(_18003_),
    .B1(_25303_),
    .Y(_18896_));
 sky130_fd_sc_hd__and3_1 _47783_ (.A(_18895_),
    .B(_18896_),
    .C(_17925_),
    .X(_18897_));
 sky130_fd_sc_hd__a21oi_1 _47784_ (.A1(_18895_),
    .A2(_18896_),
    .B1(_17925_),
    .Y(_18898_));
 sky130_fd_sc_hd__nor2_1 _47785_ (.A(_18897_),
    .B(_18898_),
    .Y(_18899_));
 sky130_fd_sc_hd__and2b_1 _47786_ (.A_N(\delay_line[10][3] ),
    .B(\delay_line[10][1] ),
    .X(_18900_));
 sky130_fd_sc_hd__clkbuf_2 _47787_ (.A(_18900_),
    .X(_18901_));
 sky130_fd_sc_hd__and2b_1 _47788_ (.A_N(\delay_line[10][1] ),
    .B(\delay_line[10][3] ),
    .X(_18902_));
 sky130_fd_sc_hd__nor3_1 _47789_ (.A(\delay_line[10][6] ),
    .B(_18901_),
    .C(_18902_),
    .Y(_18903_));
 sky130_fd_sc_hd__o21a_1 _47790_ (.A1(_18900_),
    .A2(_18902_),
    .B1(\delay_line[10][6] ),
    .X(_18904_));
 sky130_fd_sc_hd__nor2_2 _47791_ (.A(_18903_),
    .B(_18904_),
    .Y(_18905_));
 sky130_fd_sc_hd__xnor2_4 _47792_ (.A(_17909_),
    .B(_18905_),
    .Y(_18906_));
 sky130_fd_sc_hd__xnor2_2 _47793_ (.A(_18899_),
    .B(_18906_),
    .Y(_18907_));
 sky130_fd_sc_hd__o311a_1 _47794_ (.A1(_17923_),
    .A2(_17925_),
    .A3(_17922_),
    .B1(_17929_),
    .C1(_18907_),
    .X(_18908_));
 sky130_fd_sc_hd__a21oi_2 _47795_ (.A1(_17924_),
    .A2(_17929_),
    .B1(_18907_),
    .Y(_18909_));
 sky130_fd_sc_hd__nor2_1 _47796_ (.A(_18003_),
    .B(_18004_),
    .Y(_18910_));
 sky130_fd_sc_hd__a21boi_1 _47797_ (.A1(_18005_),
    .A2(_18910_),
    .B1_N(_18006_),
    .Y(_18911_));
 sky130_fd_sc_hd__o21ai_1 _47798_ (.A1(_17982_),
    .A2(_17977_),
    .B1(_17983_),
    .Y(_18912_));
 sky130_fd_sc_hd__buf_1 _47799_ (.A(\delay_line[13][6] ),
    .X(_18913_));
 sky130_fd_sc_hd__nand2_1 _47800_ (.A(\delay_line[13][4] ),
    .B(_18913_),
    .Y(_18914_));
 sky130_fd_sc_hd__clkbuf_2 _47801_ (.A(_12207_),
    .X(_18915_));
 sky130_fd_sc_hd__or2_1 _47802_ (.A(_18915_),
    .B(_18913_),
    .X(_18916_));
 sky130_fd_sc_hd__a21oi_2 _47803_ (.A1(_18914_),
    .A2(_18916_),
    .B1(_17968_),
    .Y(_18917_));
 sky130_fd_sc_hd__buf_2 _47804_ (.A(_18913_),
    .X(_18918_));
 sky130_fd_sc_hd__and4b_1 _47805_ (.A_N(_18918_),
    .B(_17967_),
    .C(_23172_),
    .D(_18915_),
    .X(_18919_));
 sky130_fd_sc_hd__buf_2 _47806_ (.A(_18919_),
    .X(_18920_));
 sky130_fd_sc_hd__a21oi_2 _47807_ (.A1(_08052_),
    .A2(_17946_),
    .B1(_17947_),
    .Y(_18921_));
 sky130_fd_sc_hd__and2_1 _47808_ (.A(_17938_),
    .B(_17944_),
    .X(_18922_));
 sky130_fd_sc_hd__clkbuf_2 _47809_ (.A(\delay_line[4][3] ),
    .X(_18923_));
 sky130_fd_sc_hd__nor2b_1 _47810_ (.A(_12240_),
    .B_N(_18923_),
    .Y(_18924_));
 sky130_fd_sc_hd__clkbuf_2 _47811_ (.A(_18924_),
    .X(_18925_));
 sky130_fd_sc_hd__and2b_1 _47812_ (.A_N(_18923_),
    .B(_12251_),
    .X(_18926_));
 sky130_fd_sc_hd__o22ai_2 _47813_ (.A1(_08129_),
    .A2(_17946_),
    .B1(_18925_),
    .B2(_18926_),
    .Y(_18927_));
 sky130_fd_sc_hd__buf_6 _47814_ (.A(\delay_line[4][3] ),
    .X(_18928_));
 sky130_fd_sc_hd__nand2b_2 _47815_ (.A_N(\delay_line[4][1] ),
    .B(_18928_),
    .Y(_18929_));
 sky130_fd_sc_hd__clkbuf_2 _47816_ (.A(_18929_),
    .X(_18930_));
 sky130_fd_sc_hd__nand2b_1 _47817_ (.A_N(_18923_),
    .B(\delay_line[4][1] ),
    .Y(_18931_));
 sky130_fd_sc_hd__nand4_2 _47818_ (.A(_17941_),
    .B(_18930_),
    .C(_18931_),
    .D(_08052_),
    .Y(_18932_));
 sky130_fd_sc_hd__clkbuf_2 _47819_ (.A(\delay_line[11][4] ),
    .X(_18933_));
 sky130_fd_sc_hd__clkbuf_2 _47820_ (.A(_18933_),
    .X(_18934_));
 sky130_fd_sc_hd__nor2_1 _47821_ (.A(\delay_line[11][0] ),
    .B(_18934_),
    .Y(_18935_));
 sky130_fd_sc_hd__clkbuf_2 _47822_ (.A(_18935_),
    .X(_18936_));
 sky130_fd_sc_hd__nand2_1 _47823_ (.A(_02502_),
    .B(_18934_),
    .Y(_18937_));
 sky130_fd_sc_hd__nand2b_1 _47824_ (.A_N(_18936_),
    .B(_18937_),
    .Y(_18938_));
 sky130_fd_sc_hd__a21oi_1 _47825_ (.A1(_18927_),
    .A2(_18932_),
    .B1(_18938_),
    .Y(_18939_));
 sky130_fd_sc_hd__and2_1 _47826_ (.A(_02502_),
    .B(_18934_),
    .X(_18940_));
 sky130_fd_sc_hd__o211a_2 _47827_ (.A1(_18936_),
    .A2(_18940_),
    .B1(_18927_),
    .C1(_18932_),
    .X(_18941_));
 sky130_fd_sc_hd__o22ai_4 _47828_ (.A1(_18921_),
    .A2(_18922_),
    .B1(_18939_),
    .B2(_18941_),
    .Y(_18942_));
 sky130_fd_sc_hd__a21o_1 _47829_ (.A1(_18927_),
    .A2(_18932_),
    .B1(_18938_),
    .X(_18943_));
 sky130_fd_sc_hd__o211ai_1 _47830_ (.A1(_18936_),
    .A2(_18940_),
    .B1(_18927_),
    .C1(_18932_),
    .Y(_18944_));
 sky130_fd_sc_hd__a21oi_1 _47831_ (.A1(_17939_),
    .A2(_17950_),
    .B1(_18921_),
    .Y(_18945_));
 sky130_fd_sc_hd__nand3_2 _47832_ (.A(_18943_),
    .B(_18944_),
    .C(_18945_),
    .Y(_18946_));
 sky130_fd_sc_hd__and2_1 _47833_ (.A(_17944_),
    .B(\delay_line[0][6] ),
    .X(_18947_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47834_ (.A(\delay_line[0][6] ),
    .X(_18948_));
 sky130_fd_sc_hd__nor2_1 _47835_ (.A(_17944_),
    .B(_18948_),
    .Y(_18949_));
 sky130_fd_sc_hd__nor2_1 _47836_ (.A(_18947_),
    .B(_18949_),
    .Y(_18950_));
 sky130_fd_sc_hd__a21oi_2 _47837_ (.A1(_18942_),
    .A2(_18946_),
    .B1(_18950_),
    .Y(_18951_));
 sky130_fd_sc_hd__nand2_1 _47838_ (.A(_17945_),
    .B(_17948_),
    .Y(_18952_));
 sky130_fd_sc_hd__a21boi_1 _47839_ (.A1(_18952_),
    .A2(_17953_),
    .B1_N(_17955_),
    .Y(_18953_));
 sky130_fd_sc_hd__nand3_1 _47840_ (.A(_18942_),
    .B(_18946_),
    .C(_18950_),
    .Y(_18954_));
 sky130_fd_sc_hd__o21ai_2 _47841_ (.A1(_17949_),
    .A2(_18953_),
    .B1(_18954_),
    .Y(_18955_));
 sky130_fd_sc_hd__or2_1 _47842_ (.A(_18947_),
    .B(_18949_),
    .X(_18956_));
 sky130_fd_sc_hd__a21o_1 _47843_ (.A1(_18942_),
    .A2(_18946_),
    .B1(_18956_),
    .X(_18957_));
 sky130_fd_sc_hd__o211ai_1 _47844_ (.A1(_18947_),
    .A2(_18949_),
    .B1(_18942_),
    .C1(_18946_),
    .Y(_18958_));
 sky130_fd_sc_hd__a21boi_1 _47845_ (.A1(_17954_),
    .A2(_17955_),
    .B1_N(_17960_),
    .Y(_18959_));
 sky130_fd_sc_hd__nand3_2 _47846_ (.A(_18957_),
    .B(_18958_),
    .C(_18959_),
    .Y(_18960_));
 sky130_fd_sc_hd__o21ai_1 _47847_ (.A1(_18951_),
    .A2(_18955_),
    .B1(_18960_),
    .Y(_18961_));
 sky130_fd_sc_hd__clkbuf_2 _47848_ (.A(net397),
    .X(_18962_));
 sky130_fd_sc_hd__a21oi_1 _47849_ (.A1(_25161_),
    .A2(_18962_),
    .B1(_08118_),
    .Y(_18963_));
 sky130_fd_sc_hd__and3_1 _47850_ (.A(_25161_),
    .B(_08118_),
    .C(_18962_),
    .X(_18964_));
 sky130_fd_sc_hd__nor2_1 _47851_ (.A(_18963_),
    .B(_18964_),
    .Y(_18965_));
 sky130_fd_sc_hd__nand2_1 _47852_ (.A(_18961_),
    .B(_18965_),
    .Y(_18966_));
 sky130_fd_sc_hd__buf_1 _47853_ (.A(_18964_),
    .X(_18967_));
 sky130_fd_sc_hd__o221ai_2 _47854_ (.A1(_18963_),
    .A2(_18967_),
    .B1(_18951_),
    .B2(_18955_),
    .C1(_18960_),
    .Y(_18968_));
 sky130_fd_sc_hd__a21oi_1 _47855_ (.A1(_17966_),
    .A2(_17970_),
    .B1(_17962_),
    .Y(_18969_));
 sky130_fd_sc_hd__nand3_2 _47856_ (.A(_18966_),
    .B(_18968_),
    .C(_18969_),
    .Y(_18970_));
 sky130_fd_sc_hd__a21o_1 _47857_ (.A1(_17966_),
    .A2(_17970_),
    .B1(_17962_),
    .X(_18971_));
 sky130_fd_sc_hd__o211ai_1 _47858_ (.A1(_18951_),
    .A2(_18955_),
    .B1(_18960_),
    .C1(_18965_),
    .Y(_18972_));
 sky130_fd_sc_hd__o21ai_1 _47859_ (.A1(_18963_),
    .A2(_18967_),
    .B1(_18961_),
    .Y(_18973_));
 sky130_fd_sc_hd__nand3_1 _47860_ (.A(_18971_),
    .B(_18972_),
    .C(_18973_),
    .Y(_18974_));
 sky130_fd_sc_hd__nand2_1 _47861_ (.A(_18970_),
    .B(_18974_),
    .Y(_18975_));
 sky130_fd_sc_hd__o21ai_1 _47862_ (.A1(_18917_),
    .A2(_18920_),
    .B1(_18975_),
    .Y(_18976_));
 sky130_fd_sc_hd__nor2_1 _47863_ (.A(_18917_),
    .B(_18920_),
    .Y(_18977_));
 sky130_fd_sc_hd__nand3_1 _47864_ (.A(_18974_),
    .B(_18977_),
    .C(_18970_),
    .Y(_18978_));
 sky130_fd_sc_hd__nand3_1 _47865_ (.A(_18912_),
    .B(_18976_),
    .C(_18978_),
    .Y(_18979_));
 sky130_fd_sc_hd__o21a_1 _47866_ (.A1(_17982_),
    .A2(_17977_),
    .B1(_17983_),
    .X(_18980_));
 sky130_fd_sc_hd__o211ai_2 _47867_ (.A1(_18917_),
    .A2(_18920_),
    .B1(_18970_),
    .C1(_18974_),
    .Y(_18981_));
 sky130_fd_sc_hd__nand2_1 _47868_ (.A(_18975_),
    .B(_18977_),
    .Y(_18982_));
 sky130_fd_sc_hd__nand3_1 _47869_ (.A(_18980_),
    .B(_18981_),
    .C(_18982_),
    .Y(_18983_));
 sky130_fd_sc_hd__clkbuf_2 _47870_ (.A(\delay_line[12][6] ),
    .X(_18984_));
 sky130_fd_sc_hd__clkbuf_2 _47871_ (.A(_18984_),
    .X(_18985_));
 sky130_fd_sc_hd__buf_2 _47872_ (.A(_18985_),
    .X(_18986_));
 sky130_fd_sc_hd__buf_2 _47873_ (.A(net406),
    .X(_18987_));
 sky130_fd_sc_hd__buf_2 _47874_ (.A(_18987_),
    .X(_18988_));
 sky130_fd_sc_hd__and2_1 _47875_ (.A(_12174_),
    .B(_18988_),
    .X(_18989_));
 sky130_fd_sc_hd__xnor2_1 _47876_ (.A(_18986_),
    .B(_18989_),
    .Y(_18990_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47877_ (.A(_18990_),
    .X(_18991_));
 sky130_fd_sc_hd__nor2_1 _47878_ (.A(_08525_),
    .B(_18991_),
    .Y(_18992_));
 sky130_fd_sc_hd__and2_1 _47879_ (.A(_08525_),
    .B(_18990_),
    .X(_18993_));
 sky130_fd_sc_hd__o2bb2ai_1 _47880_ (.A1_N(_18979_),
    .A2_N(_18983_),
    .B1(_18992_),
    .B2(_18993_),
    .Y(_18994_));
 sky130_fd_sc_hd__nor2_1 _47881_ (.A(_18992_),
    .B(_18993_),
    .Y(_18995_));
 sky130_fd_sc_hd__nand3_1 _47882_ (.A(_18979_),
    .B(_18983_),
    .C(_18995_),
    .Y(_18996_));
 sky130_fd_sc_hd__nand3_2 _47883_ (.A(_18911_),
    .B(_18994_),
    .C(_18996_),
    .Y(_18997_));
 sky130_fd_sc_hd__o21ai_1 _47884_ (.A1(_17998_),
    .A2(_18000_),
    .B1(_18005_),
    .Y(_18998_));
 sky130_fd_sc_hd__nand2_1 _47885_ (.A(_18006_),
    .B(_18998_),
    .Y(_18999_));
 sky130_fd_sc_hd__or2_1 _47886_ (.A(_18992_),
    .B(_18993_),
    .X(_19000_));
 sky130_fd_sc_hd__a21o_1 _47887_ (.A1(_18979_),
    .A2(_18983_),
    .B1(_19000_),
    .X(_19001_));
 sky130_fd_sc_hd__a31oi_2 _47888_ (.A1(_18980_),
    .A2(_18981_),
    .A3(_18982_),
    .B1(_18995_),
    .Y(_19002_));
 sky130_fd_sc_hd__nand2_1 _47889_ (.A(_19002_),
    .B(_18979_),
    .Y(_19003_));
 sky130_fd_sc_hd__nand3_2 _47890_ (.A(_18999_),
    .B(_19001_),
    .C(_19003_),
    .Y(_19004_));
 sky130_fd_sc_hd__o211ai_2 _47891_ (.A1(_18908_),
    .A2(_18909_),
    .B1(_18997_),
    .C1(_19004_),
    .Y(_19005_));
 sky130_fd_sc_hd__a21boi_2 _47892_ (.A1(_17924_),
    .A2(_17929_),
    .B1_N(_18907_),
    .Y(_19006_));
 sky130_fd_sc_hd__inv_2 _47893_ (.A(_18907_),
    .Y(_19007_));
 sky130_fd_sc_hd__o311a_1 _47894_ (.A1(_17923_),
    .A2(_17925_),
    .A3(_17922_),
    .B1(_17929_),
    .C1(_19007_),
    .X(_19008_));
 sky130_fd_sc_hd__o2bb2ai_1 _47895_ (.A1_N(_18997_),
    .A2_N(_19004_),
    .B1(_19006_),
    .B2(_19008_),
    .Y(_19009_));
 sky130_fd_sc_hd__o211ai_4 _47896_ (.A1(_18013_),
    .A2(_18894_),
    .B1(_19005_),
    .C1(_19009_),
    .Y(_19010_));
 sky130_fd_sc_hd__o2bb2ai_1 _47897_ (.A1_N(_18997_),
    .A2_N(_19004_),
    .B1(_18908_),
    .B2(_18909_),
    .Y(_19011_));
 sky130_fd_sc_hd__nor2_1 _47898_ (.A(_18016_),
    .B(_18017_),
    .Y(_19012_));
 sky130_fd_sc_hd__a32oi_2 _47899_ (.A1(_18010_),
    .A2(_18011_),
    .A3(_18012_),
    .B1(_18008_),
    .B2(_19012_),
    .Y(_19013_));
 sky130_fd_sc_hd__o211ai_1 _47900_ (.A1(_19006_),
    .A2(_19008_),
    .B1(_18997_),
    .C1(_19004_),
    .Y(_19014_));
 sky130_fd_sc_hd__nand3_2 _47901_ (.A(_19011_),
    .B(_19013_),
    .C(_19014_),
    .Y(_19015_));
 sky130_fd_sc_hd__nand2_1 _47902_ (.A(_19010_),
    .B(_19015_),
    .Y(_19016_));
 sky130_fd_sc_hd__nand2_1 _47903_ (.A(_18892_),
    .B(_19016_),
    .Y(_19017_));
 sky130_fd_sc_hd__o211ai_1 _47904_ (.A1(_18890_),
    .A2(_18891_),
    .B1(_19015_),
    .C1(_19010_),
    .Y(_19018_));
 sky130_fd_sc_hd__a21oi_1 _47905_ (.A1(_18024_),
    .A2(_18151_),
    .B1(_18153_),
    .Y(_19019_));
 sky130_fd_sc_hd__and3_2 _47906_ (.A(_19017_),
    .B(_19018_),
    .C(_19019_),
    .X(_19020_));
 sky130_fd_sc_hd__nand2_1 _47907_ (.A(_03128_),
    .B(\delay_line[7][1] ),
    .Y(_19021_));
 sky130_fd_sc_hd__nand2b_1 _47908_ (.A_N(\delay_line[7][1] ),
    .B(\delay_line[7][2] ),
    .Y(_19022_));
 sky130_fd_sc_hd__a21boi_1 _47909_ (.A1(_19021_),
    .A2(_19022_),
    .B1_N(\delay_line[7][6] ),
    .Y(_19023_));
 sky130_fd_sc_hd__buf_1 _47910_ (.A(_19023_),
    .X(_19024_));
 sky130_fd_sc_hd__and3b_1 _47911_ (.A_N(\delay_line[7][6] ),
    .B(_19021_),
    .C(_19022_),
    .X(_19025_));
 sky130_fd_sc_hd__or4_2 _47912_ (.A(_22963_),
    .B(_03447_),
    .C(_19024_),
    .D(_19025_),
    .X(_19026_));
 sky130_fd_sc_hd__a2bb2o_1 _47913_ (.A1_N(_19024_),
    .A2_N(_19025_),
    .B1(_23018_),
    .B2(_00062_),
    .X(_19027_));
 sky130_fd_sc_hd__nand4_4 _47914_ (.A(_19026_),
    .B(_19027_),
    .C(_18026_),
    .D(_11800_),
    .Y(_19028_));
 sky130_fd_sc_hd__a22o_1 _47915_ (.A1(_18026_),
    .A2(_11800_),
    .B1(_19026_),
    .B2(_19027_),
    .X(_19029_));
 sky130_fd_sc_hd__nand3b_2 _47916_ (.A_N(_18081_),
    .B(_19028_),
    .C(_19029_),
    .Y(_19030_));
 sky130_fd_sc_hd__a21bo_1 _47917_ (.A1(_19028_),
    .A2(_19029_),
    .B1_N(_18081_),
    .X(_19031_));
 sky130_fd_sc_hd__nand3_1 _47918_ (.A(_11855_),
    .B(_18042_),
    .C(_18045_),
    .Y(_19032_));
 sky130_fd_sc_hd__o21ai_1 _47919_ (.A1(_18027_),
    .A2(_18047_),
    .B1(_19032_),
    .Y(_19033_));
 sky130_fd_sc_hd__a21o_1 _47920_ (.A1(_19030_),
    .A2(_19031_),
    .B1(_19033_),
    .X(_19034_));
 sky130_fd_sc_hd__nand3_2 _47921_ (.A(_19033_),
    .B(_19030_),
    .C(_19031_),
    .Y(_19035_));
 sky130_fd_sc_hd__o21ai_1 _47922_ (.A1(_13482_),
    .A2(_18086_),
    .B1(_18084_),
    .Y(_19036_));
 sky130_fd_sc_hd__a21o_1 _47923_ (.A1(_19034_),
    .A2(_19035_),
    .B1(_19036_),
    .X(_19037_));
 sky130_fd_sc_hd__nand3_2 _47924_ (.A(_19036_),
    .B(_19034_),
    .C(_19035_),
    .Y(_19038_));
 sky130_fd_sc_hd__a21bo_1 _47925_ (.A1(_19037_),
    .A2(_19038_),
    .B1_N(_18088_),
    .X(_19039_));
 sky130_fd_sc_hd__nand3b_1 _47926_ (.A_N(_18088_),
    .B(_19037_),
    .C(_19038_),
    .Y(_19040_));
 sky130_fd_sc_hd__and2_1 _47927_ (.A(_18125_),
    .B(_18127_),
    .X(_19041_));
 sky130_fd_sc_hd__a211o_1 _47928_ (.A1(_18109_),
    .A2(_18110_),
    .B1(_18100_),
    .C1(_18102_),
    .X(_19042_));
 sky130_fd_sc_hd__inv_2 _47929_ (.A(\delay_line[5][5] ),
    .Y(_19043_));
 sky130_fd_sc_hd__buf_2 _47930_ (.A(_19043_),
    .X(_19044_));
 sky130_fd_sc_hd__clkbuf_2 _47931_ (.A(_18103_),
    .X(_19045_));
 sky130_fd_sc_hd__or4b_2 _47932_ (.A(_03568_),
    .B(_19044_),
    .C(_19045_),
    .D_N(_18098_),
    .X(_19046_));
 sky130_fd_sc_hd__buf_1 _47933_ (.A(\delay_line[3][6] ),
    .X(_19047_));
 sky130_fd_sc_hd__or2b_1 _47934_ (.A(\delay_line[3][4] ),
    .B_N(_19047_),
    .X(_19048_));
 sky130_fd_sc_hd__or2b_1 _47935_ (.A(\delay_line[3][6] ),
    .B_N(_13592_),
    .X(_19049_));
 sky130_fd_sc_hd__a22o_1 _47936_ (.A1(_13834_),
    .A2(net443),
    .B1(_19048_),
    .B2(_19049_),
    .X(_19050_));
 sky130_fd_sc_hd__clkbuf_2 _47937_ (.A(net443),
    .X(_19051_));
 sky130_fd_sc_hd__nand4_1 _47938_ (.A(_13834_),
    .B(_19048_),
    .C(_19049_),
    .D(_19051_),
    .Y(_19052_));
 sky130_fd_sc_hd__nand4_1 _47939_ (.A(_19050_),
    .B(_18101_),
    .C(_19052_),
    .D(_18099_),
    .Y(_19053_));
 sky130_fd_sc_hd__a22o_1 _47940_ (.A1(_18101_),
    .A2(_18099_),
    .B1(_19052_),
    .B2(_19050_),
    .X(_19054_));
 sky130_fd_sc_hd__nand3b_1 _47941_ (.A_N(_18122_),
    .B(_19053_),
    .C(_19054_),
    .Y(_19055_));
 sky130_fd_sc_hd__a21bo_1 _47942_ (.A1(_19053_),
    .A2(_19054_),
    .B1_N(_18122_),
    .X(_19056_));
 sky130_fd_sc_hd__nand2_1 _47943_ (.A(_19055_),
    .B(_19056_),
    .Y(_19057_));
 sky130_fd_sc_hd__a21o_1 _47944_ (.A1(_19042_),
    .A2(_19046_),
    .B1(_19057_),
    .X(_19058_));
 sky130_fd_sc_hd__nand3_1 _47945_ (.A(_19042_),
    .B(_19057_),
    .C(_19046_),
    .Y(_19059_));
 sky130_fd_sc_hd__and3b_1 _47946_ (.A_N(_19041_),
    .B(_19058_),
    .C(_19059_),
    .X(_19060_));
 sky130_fd_sc_hd__a21boi_1 _47947_ (.A1(_19058_),
    .A2(_19059_),
    .B1_N(_19041_),
    .Y(_19061_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _47948_ (.A(\delay_line[6][2] ),
    .X(_19062_));
 sky130_fd_sc_hd__nor2_1 _47949_ (.A(_19062_),
    .B(_18094_),
    .Y(_19063_));
 sky130_fd_sc_hd__nor2_1 _47950_ (.A(_13449_),
    .B(net428),
    .Y(_19064_));
 sky130_fd_sc_hd__and2_1 _47951_ (.A(\delay_line[6][4] ),
    .B(net428),
    .X(_19065_));
 sky130_fd_sc_hd__clkbuf_2 _47952_ (.A(_19065_),
    .X(_19066_));
 sky130_fd_sc_hd__o22a_1 _47953_ (.A1(_13680_),
    .A2(_19063_),
    .B1(_19064_),
    .B2(_19066_),
    .X(_19067_));
 sky130_fd_sc_hd__nor4_1 _47954_ (.A(_09437_),
    .B(_19063_),
    .C(_19064_),
    .D(_19066_),
    .Y(_19068_));
 sky130_fd_sc_hd__o32a_1 _47955_ (.A1(_18096_),
    .A2(_18095_),
    .A3(_18092_),
    .B1(_19067_),
    .B2(_19068_),
    .X(_19069_));
 sky130_fd_sc_hd__buf_1 _47956_ (.A(\delay_line[5][6] ),
    .X(_19070_));
 sky130_fd_sc_hd__a211oi_1 _47957_ (.A1(_19045_),
    .A2(_18101_),
    .B1(_19070_),
    .C1(_18107_),
    .Y(_19071_));
 sky130_fd_sc_hd__o211a_1 _47958_ (.A1(_09481_),
    .A2(_18104_),
    .B1(_19070_),
    .C1(_18103_),
    .X(_19072_));
 sky130_fd_sc_hd__nor3_2 _47959_ (.A(\delay_line[5][0] ),
    .B(_18105_),
    .C(_18106_),
    .Y(_19073_));
 sky130_fd_sc_hd__o21a_1 _47960_ (.A1(_18105_),
    .A2(_18106_),
    .B1(_22831_),
    .X(_19074_));
 sky130_fd_sc_hd__nor4_1 _47961_ (.A(_19071_),
    .B(_19072_),
    .C(_19073_),
    .D(_19074_),
    .Y(_19075_));
 sky130_fd_sc_hd__o22a_1 _47962_ (.A1(_19071_),
    .A2(_19072_),
    .B1(_19073_),
    .B2(_19074_),
    .X(_19076_));
 sky130_fd_sc_hd__nor2_1 _47963_ (.A(_19075_),
    .B(_19076_),
    .Y(_19077_));
 sky130_fd_sc_hd__o21ai_1 _47964_ (.A1(_09437_),
    .A2(_03403_),
    .B1(_22908_),
    .Y(_19078_));
 sky130_fd_sc_hd__or4_2 _47965_ (.A(_18095_),
    .B(_19078_),
    .C(_19067_),
    .D(net275),
    .X(_19079_));
 sky130_fd_sc_hd__nand3b_2 _47966_ (.A_N(_19069_),
    .B(_19077_),
    .C(_19079_),
    .Y(_19080_));
 sky130_fd_sc_hd__clkbuf_2 _47967_ (.A(_18095_),
    .X(_19081_));
 sky130_fd_sc_hd__nor4_1 _47968_ (.A(_19081_),
    .B(_19078_),
    .C(_19067_),
    .D(net275),
    .Y(_19082_));
 sky130_fd_sc_hd__o22ai_2 _47969_ (.A1(_19075_),
    .A2(_19076_),
    .B1(net261),
    .B2(_19069_),
    .Y(_19083_));
 sky130_fd_sc_hd__nand2_1 _47970_ (.A(_19080_),
    .B(_19083_),
    .Y(_19084_));
 sky130_fd_sc_hd__xor2_1 _47971_ (.A(net211),
    .B(_19084_),
    .X(_19085_));
 sky130_fd_sc_hd__o21a_1 _47972_ (.A1(_19060_),
    .A2(_19061_),
    .B1(_19085_),
    .X(_19086_));
 sky130_fd_sc_hd__nor3_1 _47973_ (.A(_19060_),
    .B(_19061_),
    .C(_19085_),
    .Y(_19087_));
 sky130_fd_sc_hd__nor2_1 _47974_ (.A(_19086_),
    .B(_19087_),
    .Y(_19088_));
 sky130_fd_sc_hd__a21o_1 _47975_ (.A1(_19039_),
    .A2(_19040_),
    .B1(_19088_),
    .X(_19089_));
 sky130_fd_sc_hd__nand3_1 _47976_ (.A(_19039_),
    .B(_19040_),
    .C(_19088_),
    .Y(_19090_));
 sky130_fd_sc_hd__a211oi_2 _47977_ (.A1(_19089_),
    .A2(_19090_),
    .B1(_18149_),
    .C1(_18148_),
    .Y(_19091_));
 sky130_fd_sc_hd__a21bo_1 _47978_ (.A1(_18136_),
    .A2(_18091_),
    .B1_N(_18090_),
    .X(_19092_));
 sky130_fd_sc_hd__inv_2 _47979_ (.A(_19092_),
    .Y(_19093_));
 sky130_fd_sc_hd__o211ai_2 _47980_ (.A1(_18149_),
    .A2(_18148_),
    .B1(_19089_),
    .C1(_19090_),
    .Y(_19094_));
 sky130_fd_sc_hd__o21ai_2 _47981_ (.A1(_19093_),
    .A2(_19091_),
    .B1(_19094_),
    .Y(_19095_));
 sky130_fd_sc_hd__inv_2 _47982_ (.A(_19094_),
    .Y(_19096_));
 sky130_fd_sc_hd__o21ai_1 _47983_ (.A1(_19096_),
    .A2(_19091_),
    .B1(_19092_),
    .Y(_19097_));
 sky130_fd_sc_hd__o21ai_1 _47984_ (.A1(_19091_),
    .A2(_19095_),
    .B1(_19097_),
    .Y(_19098_));
 sky130_fd_sc_hd__a31oi_2 _47985_ (.A1(_18022_),
    .A2(_18020_),
    .A3(_18021_),
    .B1(_18073_),
    .Y(_19099_));
 sky130_fd_sc_hd__nand3_2 _47986_ (.A(_19010_),
    .B(_18892_),
    .C(_19015_),
    .Y(_19100_));
 sky130_fd_sc_hd__a21o_1 _47987_ (.A1(_19010_),
    .A2(_19015_),
    .B1(_18892_),
    .X(_19101_));
 sky130_fd_sc_hd__o211ai_4 _47988_ (.A1(_18153_),
    .A2(_19099_),
    .B1(_19100_),
    .C1(_19101_),
    .Y(_19102_));
 sky130_fd_sc_hd__nand2_1 _47989_ (.A(_19098_),
    .B(_19102_),
    .Y(_19103_));
 sky130_fd_sc_hd__nand3_1 _47990_ (.A(_19017_),
    .B(_19018_),
    .C(_19019_),
    .Y(_19104_));
 sky130_fd_sc_hd__nand2_1 _47991_ (.A(_19104_),
    .B(_19102_),
    .Y(_19105_));
 sky130_fd_sc_hd__o21a_2 _47992_ (.A1(_19091_),
    .A2(_19095_),
    .B1(_19097_),
    .X(_19106_));
 sky130_fd_sc_hd__nand2_1 _47993_ (.A(_19105_),
    .B(_19106_),
    .Y(_19107_));
 sky130_fd_sc_hd__o221ai_4 _47994_ (.A1(_18841_),
    .A2(_18146_),
    .B1(_19020_),
    .B2(_19103_),
    .C1(_19107_),
    .Y(_19108_));
 sky130_fd_sc_hd__nand2_1 _47995_ (.A(_19098_),
    .B(_19105_),
    .Y(_19109_));
 sky130_fd_sc_hd__a21oi_1 _47996_ (.A1(_18160_),
    .A2(_18145_),
    .B1(_18841_),
    .Y(_19110_));
 sky130_fd_sc_hd__nand3_1 _47997_ (.A(_19106_),
    .B(_19104_),
    .C(_19102_),
    .Y(_19111_));
 sky130_fd_sc_hd__nand3_4 _47998_ (.A(_19109_),
    .B(_19110_),
    .C(_19111_),
    .Y(_19112_));
 sky130_fd_sc_hd__o21ai_1 _47999_ (.A1(_18199_),
    .A2(_18196_),
    .B1(_18197_),
    .Y(_19113_));
 sky130_fd_sc_hd__o2bb2a_1 _48000_ (.A1_N(_18171_),
    .A2_N(_18175_),
    .B1(_14361_),
    .B2(_18177_),
    .X(_19114_));
 sky130_fd_sc_hd__o21ai_1 _48001_ (.A1(_18181_),
    .A2(_19114_),
    .B1(_18176_),
    .Y(_19115_));
 sky130_fd_sc_hd__clkbuf_2 _48002_ (.A(_14317_),
    .X(_19116_));
 sky130_fd_sc_hd__clkbuf_2 _48003_ (.A(\delay_line[1][5] ),
    .X(_19117_));
 sky130_fd_sc_hd__clkbuf_2 _48004_ (.A(_19117_),
    .X(_19118_));
 sky130_fd_sc_hd__o21a_1 _48005_ (.A1(_19116_),
    .A2(_19118_),
    .B1(_14284_),
    .X(_19119_));
 sky130_fd_sc_hd__nor3_1 _48006_ (.A(_19116_),
    .B(_19118_),
    .C(_14284_),
    .Y(_19120_));
 sky130_fd_sc_hd__clkbuf_2 _48007_ (.A(\delay_line[1][6] ),
    .X(_19121_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48008_ (.A(\delay_line[1][6] ),
    .X(_19122_));
 sky130_fd_sc_hd__o21ai_1 _48009_ (.A1(_09305_),
    .A2(_19122_),
    .B1(\delay_line[2][6] ),
    .Y(_19123_));
 sky130_fd_sc_hd__a21o_1 _48010_ (.A1(_09305_),
    .A2(_19121_),
    .B1(_19123_),
    .X(_19124_));
 sky130_fd_sc_hd__and2_1 _48011_ (.A(_09305_),
    .B(_19122_),
    .X(_19125_));
 sky130_fd_sc_hd__nor2_1 _48012_ (.A(_09305_),
    .B(_19122_),
    .Y(_19126_));
 sky130_fd_sc_hd__o21bai_2 _48013_ (.A1(_19125_),
    .A2(_19126_),
    .B1_N(\delay_line[2][6] ),
    .Y(_19127_));
 sky130_fd_sc_hd__nand3b_2 _48014_ (.A_N(_18171_),
    .B(_19124_),
    .C(_19127_),
    .Y(_19128_));
 sky130_fd_sc_hd__or2_1 _48015_ (.A(_18169_),
    .B(_18173_),
    .X(_19129_));
 sky130_fd_sc_hd__o2bb2ai_1 _48016_ (.A1_N(_19124_),
    .A2_N(_19127_),
    .B1(_03678_),
    .B2(_19129_),
    .Y(_19130_));
 sky130_fd_sc_hd__o211ai_2 _48017_ (.A1(_19119_),
    .A2(_19120_),
    .B1(_19128_),
    .C1(_19130_),
    .Y(_19131_));
 sky130_fd_sc_hd__o21a_1 _48018_ (.A1(_19116_),
    .A2(_19118_),
    .B1(_09756_),
    .X(_19132_));
 sky130_fd_sc_hd__nor3_1 _48019_ (.A(_19116_),
    .B(_19118_),
    .C(_09800_),
    .Y(_19133_));
 sky130_fd_sc_hd__o2bb2ai_1 _48020_ (.A1_N(_19128_),
    .A2_N(_19130_),
    .B1(_19132_),
    .B2(_19133_),
    .Y(_19134_));
 sky130_fd_sc_hd__nand3_1 _48021_ (.A(_19115_),
    .B(_19131_),
    .C(_19134_),
    .Y(_19135_));
 sky130_fd_sc_hd__a21o_1 _48022_ (.A1(_19131_),
    .A2(_19134_),
    .B1(_19115_),
    .X(_19136_));
 sky130_fd_sc_hd__o21a_1 _48023_ (.A1(_09822_),
    .A2(_09800_),
    .B1(_14372_),
    .X(_19137_));
 sky130_fd_sc_hd__and3_1 _48024_ (.A(_19135_),
    .B(_19136_),
    .C(_19137_),
    .X(_19138_));
 sky130_fd_sc_hd__a21oi_1 _48025_ (.A1(_19135_),
    .A2(_19136_),
    .B1(_19137_),
    .Y(_19139_));
 sky130_fd_sc_hd__o21bai_1 _48026_ (.A1(_18132_),
    .A2(_18131_),
    .B1_N(_18129_),
    .Y(_19140_));
 sky130_fd_sc_hd__o21bai_1 _48027_ (.A1(_19138_),
    .A2(_19139_),
    .B1_N(_19140_),
    .Y(_19141_));
 sky130_fd_sc_hd__o2111ai_2 _48028_ (.A1(_09822_),
    .A2(_09800_),
    .B1(_14372_),
    .C1(_19135_),
    .D1(_19136_),
    .Y(_19142_));
 sky130_fd_sc_hd__a21o_1 _48029_ (.A1(_19135_),
    .A2(_19136_),
    .B1(_19137_),
    .X(_19143_));
 sky130_fd_sc_hd__nand3_1 _48030_ (.A(_19140_),
    .B(_19142_),
    .C(_19143_),
    .Y(_19144_));
 sky130_fd_sc_hd__o21ai_1 _48031_ (.A1(_18188_),
    .A2(_18189_),
    .B1(_18185_),
    .Y(_19145_));
 sky130_fd_sc_hd__a21oi_1 _48032_ (.A1(_19141_),
    .A2(_19144_),
    .B1(_19145_),
    .Y(_19146_));
 sky130_fd_sc_hd__and3_1 _48033_ (.A(_19145_),
    .B(_19141_),
    .C(_19144_),
    .X(_19147_));
 sky130_fd_sc_hd__or3_1 _48034_ (.A(_13735_),
    .B(net212),
    .C(_18114_),
    .X(_19148_));
 sky130_fd_sc_hd__o221ai_2 _48035_ (.A1(_18116_),
    .A2(_18135_),
    .B1(_19146_),
    .B2(_19147_),
    .C1(_19148_),
    .Y(_19149_));
 sky130_fd_sc_hd__nand3_1 _48036_ (.A(_18117_),
    .B(_18133_),
    .C(_18134_),
    .Y(_19150_));
 sky130_fd_sc_hd__a211o_1 _48037_ (.A1(_19148_),
    .A2(_19150_),
    .B1(_19146_),
    .C1(_19147_),
    .X(_19151_));
 sky130_fd_sc_hd__nand2_1 _48038_ (.A(_18191_),
    .B(_18194_),
    .Y(_19152_));
 sky130_fd_sc_hd__a21o_1 _48039_ (.A1(_19149_),
    .A2(_19151_),
    .B1(_19152_),
    .X(_19153_));
 sky130_fd_sc_hd__nand3_1 _48040_ (.A(_19152_),
    .B(_19149_),
    .C(_19151_),
    .Y(_19154_));
 sky130_fd_sc_hd__and3_1 _48041_ (.A(_19113_),
    .B(_19153_),
    .C(_19154_),
    .X(_19155_));
 sky130_fd_sc_hd__nand2_1 _48042_ (.A(_19153_),
    .B(_19154_),
    .Y(_19156_));
 sky130_fd_sc_hd__o211a_1 _48043_ (.A1(_18199_),
    .A2(_18196_),
    .B1(_18197_),
    .C1(_19156_),
    .X(_19157_));
 sky130_fd_sc_hd__o21a_1 _48044_ (.A1(_18140_),
    .A2(_18144_),
    .B1(_18141_),
    .X(_19158_));
 sky130_fd_sc_hd__o21ai_1 _48045_ (.A1(_19155_),
    .A2(_19157_),
    .B1(_19158_),
    .Y(_19159_));
 sky130_fd_sc_hd__nand2_1 _48046_ (.A(_19159_),
    .B(_18202_),
    .Y(_19160_));
 sky130_fd_sc_hd__inv_2 _48047_ (.A(_19160_),
    .Y(_19161_));
 sky130_fd_sc_hd__nor3_2 _48048_ (.A(_19158_),
    .B(_19155_),
    .C(_19157_),
    .Y(_19162_));
 sky130_fd_sc_hd__inv_2 _48049_ (.A(_19162_),
    .Y(_19163_));
 sky130_fd_sc_hd__nand2_1 _48050_ (.A(_19161_),
    .B(_19163_),
    .Y(_19164_));
 sky130_fd_sc_hd__and3_1 _48051_ (.A(_19164_),
    .B(_18201_),
    .C(_18203_),
    .X(_19165_));
 sky130_fd_sc_hd__and3_1 _48052_ (.A(_19163_),
    .B(_19159_),
    .C(_19160_),
    .X(_19166_));
 sky130_fd_sc_hd__o2bb2ai_1 _48053_ (.A1_N(_19108_),
    .A2_N(_19112_),
    .B1(_19165_),
    .B2(_19166_),
    .Y(_19167_));
 sky130_fd_sc_hd__a21boi_1 _48054_ (.A1(_18167_),
    .A2(_18210_),
    .B1_N(_18163_),
    .Y(_19168_));
 sky130_fd_sc_hd__inv_2 _48055_ (.A(_19164_),
    .Y(_19169_));
 sky130_fd_sc_hd__a21oi_1 _48056_ (.A1(_19163_),
    .A2(_19159_),
    .B1(_18202_),
    .Y(_19170_));
 sky130_fd_sc_hd__clkbuf_2 _48057_ (.A(_19108_),
    .X(_19171_));
 sky130_fd_sc_hd__o211ai_2 _48058_ (.A1(_19169_),
    .A2(_19170_),
    .B1(_19171_),
    .C1(_19112_),
    .Y(_19172_));
 sky130_fd_sc_hd__nand3_4 _48059_ (.A(_19167_),
    .B(_19168_),
    .C(_19172_),
    .Y(_19173_));
 sky130_fd_sc_hd__nor2_1 _48060_ (.A(_18215_),
    .B(net94),
    .Y(_19174_));
 sky130_fd_sc_hd__a21oi_2 _48061_ (.A1(_18158_),
    .A2(_18161_),
    .B1(_17908_),
    .Y(_19175_));
 sky130_fd_sc_hd__o21ai_2 _48062_ (.A1(_19174_),
    .A2(_19175_),
    .B1(_18163_),
    .Y(_19176_));
 sky130_fd_sc_hd__o211ai_2 _48063_ (.A1(_19165_),
    .A2(_19166_),
    .B1(_19171_),
    .C1(_19112_),
    .Y(_19177_));
 sky130_fd_sc_hd__o2bb2ai_2 _48064_ (.A1_N(_19171_),
    .A2_N(_19112_),
    .B1(_19169_),
    .B2(_19170_),
    .Y(_19178_));
 sky130_fd_sc_hd__nand3_4 _48065_ (.A(_19176_),
    .B(_19177_),
    .C(_19178_),
    .Y(_19179_));
 sky130_fd_sc_hd__o211ai_4 _48066_ (.A1(_18216_),
    .A2(_18840_),
    .B1(_19173_),
    .C1(_19179_),
    .Y(_19180_));
 sky130_fd_sc_hd__nor2_1 _48067_ (.A(_18216_),
    .B(_18840_),
    .Y(_19181_));
 sky130_fd_sc_hd__inv_2 _48068_ (.A(_19181_),
    .Y(_19182_));
 sky130_fd_sc_hd__a21o_1 _48069_ (.A1(_19179_),
    .A2(_19173_),
    .B1(_19182_),
    .X(_19183_));
 sky130_fd_sc_hd__nand3_2 _48070_ (.A(_18839_),
    .B(_19180_),
    .C(_19183_),
    .Y(_19184_));
 sky130_fd_sc_hd__inv_2 _48071_ (.A(_18230_),
    .Y(_19185_));
 sky130_fd_sc_hd__a21oi_2 _48072_ (.A1(_18231_),
    .A2(_18232_),
    .B1(_18229_),
    .Y(_19186_));
 sky130_fd_sc_hd__o211a_2 _48073_ (.A1(_18216_),
    .A2(_18840_),
    .B1(_19173_),
    .C1(_19179_),
    .X(_19187_));
 sky130_fd_sc_hd__a21oi_2 _48074_ (.A1(_19179_),
    .A2(_19173_),
    .B1(_19182_),
    .Y(_19188_));
 sky130_fd_sc_hd__o22ai_4 _48075_ (.A1(_19185_),
    .A2(_19186_),
    .B1(_19187_),
    .B2(_19188_),
    .Y(_19189_));
 sky130_fd_sc_hd__a31o_1 _48076_ (.A1(_18229_),
    .A2(_18230_),
    .A3(_18233_),
    .B1(_18226_),
    .X(_19190_));
 sky130_fd_sc_hd__a21oi_1 _48077_ (.A1(_18227_),
    .A2(_18224_),
    .B1(_19190_),
    .Y(_19191_));
 sky130_fd_sc_hd__a221oi_4 _48078_ (.A1(_17905_),
    .A2(_18238_),
    .B1(_19184_),
    .B2(_19189_),
    .C1(_19191_),
    .Y(_19192_));
 sky130_fd_sc_hd__nand2_2 _48079_ (.A(_19184_),
    .B(_19189_),
    .Y(_19193_));
 sky130_fd_sc_hd__a22oi_4 _48080_ (.A1(_18234_),
    .A2(_18235_),
    .B1(_17904_),
    .B2(_18237_),
    .Y(_19194_));
 sky130_fd_sc_hd__o21ai_2 _48081_ (.A1(_19193_),
    .A2(_19194_),
    .B1(\delay_line[23][6] ),
    .Y(_19195_));
 sky130_fd_sc_hd__nand2_1 _48082_ (.A(_19194_),
    .B(_19193_),
    .Y(_19196_));
 sky130_fd_sc_hd__inv_2 _48083_ (.A(_18235_),
    .Y(_19197_));
 sky130_fd_sc_hd__o2bb2ai_1 _48084_ (.A1_N(_17905_),
    .A2_N(_18237_),
    .B1(_19190_),
    .B2(_19197_),
    .Y(_19198_));
 sky130_fd_sc_hd__a31o_1 _48085_ (.A1(_18220_),
    .A2(_18221_),
    .A3(_18222_),
    .B1(_18227_),
    .X(_19199_));
 sky130_fd_sc_hd__a21oi_1 _48086_ (.A1(_18233_),
    .A2(_19199_),
    .B1(_19188_),
    .Y(_19200_));
 sky130_fd_sc_hd__a2bb2oi_2 _48087_ (.A1_N(_19185_),
    .A2_N(_19186_),
    .B1(_19180_),
    .B2(_19183_),
    .Y(_19201_));
 sky130_fd_sc_hd__a21oi_1 _48088_ (.A1(_19180_),
    .A2(_19200_),
    .B1(_19201_),
    .Y(_19202_));
 sky130_fd_sc_hd__nand2_1 _48089_ (.A(_19198_),
    .B(_19202_),
    .Y(_19203_));
 sky130_fd_sc_hd__clkbuf_2 _48090_ (.A(\delay_line[23][6] ),
    .X(_19204_));
 sky130_fd_sc_hd__a21o_1 _48091_ (.A1(_19196_),
    .A2(_19203_),
    .B1(_19204_),
    .X(_19205_));
 sky130_fd_sc_hd__o211ai_4 _48092_ (.A1(_19192_),
    .A2(_19195_),
    .B1(_18836_),
    .C1(_19205_),
    .Y(_19206_));
 sky130_fd_sc_hd__nor2_1 _48093_ (.A(_19192_),
    .B(_19195_),
    .Y(_19207_));
 sky130_fd_sc_hd__a21oi_1 _48094_ (.A1(_19196_),
    .A2(_19203_),
    .B1(_19204_),
    .Y(_19208_));
 sky130_fd_sc_hd__o21bai_4 _48095_ (.A1(_19207_),
    .A2(_19208_),
    .B1_N(_18836_),
    .Y(_19209_));
 sky130_fd_sc_hd__o211ai_4 _48096_ (.A1(_18621_),
    .A2(_18838_),
    .B1(_19206_),
    .C1(_19209_),
    .Y(_19210_));
 sky130_fd_sc_hd__a41o_1 _48097_ (.A1(_18600_),
    .A2(_18601_),
    .A3(_18619_),
    .A4(_18620_),
    .B1(_18838_),
    .X(_19211_));
 sky130_fd_sc_hd__a21o_1 _48098_ (.A1(_19206_),
    .A2(_19209_),
    .B1(_19211_),
    .X(_19212_));
 sky130_fd_sc_hd__o211ai_1 _48099_ (.A1(_17903_),
    .A2(_18837_),
    .B1(_19210_),
    .C1(_19212_),
    .Y(_19213_));
 sky130_fd_sc_hd__o211a_1 _48100_ (.A1(_18621_),
    .A2(_18838_),
    .B1(_19206_),
    .C1(_19209_),
    .X(_19214_));
 sky130_fd_sc_hd__a21oi_4 _48101_ (.A1(_19206_),
    .A2(_19209_),
    .B1(_19211_),
    .Y(_19215_));
 sky130_fd_sc_hd__buf_2 _48102_ (.A(_18836_),
    .X(_19216_));
 sky130_fd_sc_hd__nand2_2 _48103_ (.A(_18259_),
    .B(_19216_),
    .Y(_19217_));
 sky130_fd_sc_hd__o31a_2 _48104_ (.A1(_17901_),
    .A2(_18243_),
    .A3(_18244_),
    .B1(_19217_),
    .X(_19218_));
 sky130_fd_sc_hd__o21ai_1 _48105_ (.A1(_19214_),
    .A2(_19215_),
    .B1(_19218_),
    .Y(_19219_));
 sky130_fd_sc_hd__o211ai_1 _48106_ (.A1(_18583_),
    .A2(_18625_),
    .B1(_19213_),
    .C1(_19219_),
    .Y(_19220_));
 sky130_fd_sc_hd__buf_2 _48107_ (.A(_19220_),
    .X(_19221_));
 sky130_fd_sc_hd__o22ai_4 _48108_ (.A1(_17903_),
    .A2(_18837_),
    .B1(_19214_),
    .B2(_19215_),
    .Y(_19222_));
 sky130_fd_sc_hd__nor2_1 _48109_ (.A(_18583_),
    .B(_18625_),
    .Y(_19223_));
 sky130_fd_sc_hd__nand3_2 _48110_ (.A(_19212_),
    .B(_19218_),
    .C(_19210_),
    .Y(_19224_));
 sky130_fd_sc_hd__a21o_1 _48111_ (.A1(_18260_),
    .A2(_18258_),
    .B1(_18247_),
    .X(_19225_));
 sky130_fd_sc_hd__inv_2 _48112_ (.A(_19225_),
    .Y(_19226_));
 sky130_fd_sc_hd__a31oi_2 _48113_ (.A1(_19222_),
    .A2(_19223_),
    .A3(_19224_),
    .B1(_19226_),
    .Y(_19227_));
 sky130_fd_sc_hd__o31a_1 _48114_ (.A1(_15119_),
    .A2(_18274_),
    .A3(_18275_),
    .B1(_18266_),
    .X(_19228_));
 sky130_fd_sc_hd__inv_2 _48115_ (.A(_19228_),
    .Y(_19229_));
 sky130_fd_sc_hd__nand3_2 _48116_ (.A(_19222_),
    .B(_19223_),
    .C(_19224_),
    .Y(_19230_));
 sky130_fd_sc_hd__a21oi_4 _48117_ (.A1(_19221_),
    .A2(_19230_),
    .B1(_19225_),
    .Y(_19231_));
 sky130_fd_sc_hd__a211oi_2 _48118_ (.A1(_19221_),
    .A2(_19227_),
    .B1(_19229_),
    .C1(_19231_),
    .Y(_19232_));
 sky130_fd_sc_hd__nand2_2 _48119_ (.A(_19227_),
    .B(_19221_),
    .Y(_19233_));
 sky130_fd_sc_hd__a21o_1 _48120_ (.A1(_19221_),
    .A2(_19230_),
    .B1(_19225_),
    .X(_19234_));
 sky130_fd_sc_hd__a21oi_4 _48121_ (.A1(_19233_),
    .A2(_19234_),
    .B1(_19228_),
    .Y(_19235_));
 sky130_fd_sc_hd__clkbuf_2 _48122_ (.A(_18259_),
    .X(_19236_));
 sky130_fd_sc_hd__nor2_1 _48123_ (.A(_07909_),
    .B(_19236_),
    .Y(_19237_));
 sky130_fd_sc_hd__and2_1 _48124_ (.A(_00370_),
    .B(_18259_),
    .X(_19238_));
 sky130_fd_sc_hd__and4bb_2 _48125_ (.A_N(_19237_),
    .B_N(_19238_),
    .C(_17895_),
    .D(_17898_),
    .X(_19239_));
 sky130_fd_sc_hd__o2bb2a_2 _48126_ (.A1_N(_17895_),
    .A2_N(_17898_),
    .B1(_19237_),
    .B2(_19238_),
    .X(_19240_));
 sky130_fd_sc_hd__or2_1 _48127_ (.A(_19239_),
    .B(_19240_),
    .X(_19241_));
 sky130_fd_sc_hd__inv_2 _48128_ (.A(_19241_),
    .Y(_19242_));
 sky130_fd_sc_hd__o21ai_1 _48129_ (.A1(net60),
    .A2(_19235_),
    .B1(_19242_),
    .Y(_19243_));
 sky130_fd_sc_hd__a21oi_2 _48130_ (.A1(_16261_),
    .A2(_16305_),
    .B1(_18700_),
    .Y(_19244_));
 sky130_fd_sc_hd__a21oi_1 _48131_ (.A1(_18703_),
    .A2(_18701_),
    .B1(_19244_),
    .Y(_19245_));
 sky130_fd_sc_hd__o2111ai_4 _48132_ (.A1(_18267_),
    .A2(_18275_),
    .B1(_18266_),
    .C1(_19233_),
    .D1(_19234_),
    .Y(_19246_));
 sky130_fd_sc_hd__and3_2 _48133_ (.A(_19220_),
    .B(_19230_),
    .C(_19225_),
    .X(_19247_));
 sky130_fd_sc_hd__o21ai_2 _48134_ (.A1(_19247_),
    .A2(_19231_),
    .B1(_19229_),
    .Y(_19248_));
 sky130_fd_sc_hd__o211ai_1 _48135_ (.A1(_19239_),
    .A2(_19240_),
    .B1(_19246_),
    .C1(_19248_),
    .Y(_19249_));
 sky130_fd_sc_hd__nand3_1 _48136_ (.A(_19243_),
    .B(_19245_),
    .C(_19249_),
    .Y(_19250_));
 sky130_fd_sc_hd__clkbuf_2 _48137_ (.A(_19250_),
    .X(_19251_));
 sky130_fd_sc_hd__nand3_1 _48138_ (.A(_19248_),
    .B(_19242_),
    .C(_19246_),
    .Y(_19252_));
 sky130_fd_sc_hd__o22ai_4 _48139_ (.A1(_19239_),
    .A2(_19240_),
    .B1(net60),
    .B2(_19235_),
    .Y(_19253_));
 sky130_fd_sc_hd__o211ai_2 _48140_ (.A1(_19244_),
    .A2(_18705_),
    .B1(_19252_),
    .C1(_19253_),
    .Y(_19254_));
 sky130_fd_sc_hd__o21ai_2 _48141_ (.A1(_18284_),
    .A2(_18288_),
    .B1(_18297_),
    .Y(_19255_));
 sky130_fd_sc_hd__a21oi_1 _48142_ (.A1(_19251_),
    .A2(_19254_),
    .B1(_19255_),
    .Y(_19256_));
 sky130_fd_sc_hd__o221a_2 _48143_ (.A1(_18270_),
    .A2(_18272_),
    .B1(_15273_),
    .B2(_18295_),
    .C1(_18296_),
    .X(_19257_));
 sky130_fd_sc_hd__o21a_1 _48144_ (.A1(_17899_),
    .A2(_17900_),
    .B1(_18279_),
    .X(_19258_));
 sky130_fd_sc_hd__o211a_1 _48145_ (.A1(_19257_),
    .A2(_19258_),
    .B1(_19251_),
    .C1(_19254_),
    .X(_19259_));
 sky130_fd_sc_hd__a21o_1 _48146_ (.A1(_18544_),
    .A2(_18706_),
    .B1(_18543_),
    .X(_19260_));
 sky130_fd_sc_hd__o21bai_2 _48147_ (.A1(_18537_),
    .A2(_18538_),
    .B1_N(_18449_),
    .Y(_19261_));
 sky130_fd_sc_hd__o21a_1 _48148_ (.A1(_16481_),
    .A2(net173),
    .B1(_18339_),
    .X(_19262_));
 sky130_fd_sc_hd__and2_1 _48149_ (.A(_18485_),
    .B(_01161_),
    .X(_19263_));
 sky130_fd_sc_hd__clkbuf_2 _48150_ (.A(net338),
    .X(_19264_));
 sky130_fd_sc_hd__o21ai_1 _48151_ (.A1(_24314_),
    .A2(_01172_),
    .B1(_19264_),
    .Y(_19265_));
 sky130_fd_sc_hd__buf_1 _48152_ (.A(\delay_line[26][1] ),
    .X(_19266_));
 sky130_fd_sc_hd__nor2_1 _48153_ (.A(_24314_),
    .B(_19266_),
    .Y(_19267_));
 sky130_fd_sc_hd__o21bai_1 _48154_ (.A1(_19263_),
    .A2(_19267_),
    .B1_N(_19264_),
    .Y(_19268_));
 sky130_fd_sc_hd__o21a_1 _48155_ (.A1(_19263_),
    .A2(_19265_),
    .B1(_19268_),
    .X(_19269_));
 sky130_fd_sc_hd__nand2_1 _48156_ (.A(_18490_),
    .B(_19269_),
    .Y(_19270_));
 sky130_fd_sc_hd__clkbuf_2 _48157_ (.A(_18488_),
    .X(_19271_));
 sky130_fd_sc_hd__a21o_1 _48158_ (.A1(_24314_),
    .A2(_19271_),
    .B1(_19269_),
    .X(_19272_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48159_ (.A(\delay_line[27][6] ),
    .X(_19273_));
 sky130_fd_sc_hd__or2b_1 _48160_ (.A(_18492_),
    .B_N(_18493_),
    .X(_19274_));
 sky130_fd_sc_hd__nor2_1 _48161_ (.A(_16042_),
    .B(net332),
    .Y(_19275_));
 sky130_fd_sc_hd__nand2_1 _48162_ (.A(_16042_),
    .B(_19273_),
    .Y(_19276_));
 sky130_fd_sc_hd__nand3b_1 _48163_ (.A_N(_19275_),
    .B(_18495_),
    .C(_19276_),
    .Y(_19277_));
 sky130_fd_sc_hd__and2_1 _48164_ (.A(\delay_line[27][4] ),
    .B(net332),
    .X(_19278_));
 sky130_fd_sc_hd__buf_1 _48165_ (.A(_19278_),
    .X(_19279_));
 sky130_fd_sc_hd__o21ai_1 _48166_ (.A1(_19279_),
    .A2(_19275_),
    .B1(_18493_),
    .Y(_19280_));
 sky130_fd_sc_hd__a2bb2o_1 _48167_ (.A1_N(_18496_),
    .A2_N(_19274_),
    .B1(_19277_),
    .B2(_19280_),
    .X(_19281_));
 sky130_fd_sc_hd__o211ai_1 _48168_ (.A1(_19273_),
    .A2(_18494_),
    .B1(_22468_),
    .C1(_19281_),
    .Y(_19282_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48169_ (.A(_19282_),
    .X(_19283_));
 sky130_fd_sc_hd__nor2_1 _48170_ (.A(_19273_),
    .B(_18494_),
    .Y(_19284_));
 sky130_fd_sc_hd__nor3_1 _48171_ (.A(_19275_),
    .B(_18493_),
    .C(_19278_),
    .Y(_19285_));
 sky130_fd_sc_hd__o2bb2a_1 _48172_ (.A1_N(_06491_),
    .A2_N(_18491_),
    .B1(_19279_),
    .B2(_19275_),
    .X(_19286_));
 sky130_fd_sc_hd__o32a_1 _48173_ (.A1(_18496_),
    .A2(_18492_),
    .A3(_18495_),
    .B1(_19285_),
    .B2(_19286_),
    .X(_19287_));
 sky130_fd_sc_hd__o21bai_1 _48174_ (.A1(_19284_),
    .A2(_19287_),
    .B1_N(_22457_),
    .Y(_19288_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48175_ (.A(_19288_),
    .X(_19289_));
 sky130_fd_sc_hd__o2111a_1 _48176_ (.A1(_16108_),
    .A2(_18491_),
    .B1(_19283_),
    .C1(_18504_),
    .D1(_19289_),
    .X(_19290_));
 sky130_fd_sc_hd__a2111oi_1 _48177_ (.A1(_16097_),
    .A2(_18499_),
    .B1(_18500_),
    .C1(_16053_),
    .D1(_06579_),
    .Y(_19291_));
 sky130_fd_sc_hd__a2bb2oi_2 _48178_ (.A1_N(_18501_),
    .A2_N(net209),
    .B1(_19283_),
    .B2(_19289_),
    .Y(_19292_));
 sky130_fd_sc_hd__a211oi_2 _48179_ (.A1(_19270_),
    .A2(_19272_),
    .B1(_19290_),
    .C1(_19292_),
    .Y(_19293_));
 sky130_fd_sc_hd__o211a_1 _48180_ (.A1(_19290_),
    .A2(_19292_),
    .B1(_19270_),
    .C1(_19272_),
    .X(_19294_));
 sky130_fd_sc_hd__buf_1 _48181_ (.A(\delay_line[28][6] ),
    .X(_19295_));
 sky130_fd_sc_hd__nor2_1 _48182_ (.A(\delay_line[28][5] ),
    .B(_19295_),
    .Y(_19296_));
 sky130_fd_sc_hd__and2_1 _48183_ (.A(\delay_line[28][5] ),
    .B(_19295_),
    .X(_19297_));
 sky130_fd_sc_hd__nand2_1 _48184_ (.A(\delay_line[28][4] ),
    .B(_18510_),
    .Y(_19298_));
 sky130_fd_sc_hd__o21ai_2 _48185_ (.A1(_19296_),
    .A2(_19297_),
    .B1(_19298_),
    .Y(_19299_));
 sky130_fd_sc_hd__inv_2 _48186_ (.A(\delay_line[28][6] ),
    .Y(_19300_));
 sky130_fd_sc_hd__clkbuf_2 _48187_ (.A(_19300_),
    .X(_19301_));
 sky130_fd_sc_hd__nand2_1 _48188_ (.A(_18513_),
    .B(_19301_),
    .Y(_19302_));
 sky130_fd_sc_hd__a21oi_1 _48189_ (.A1(_19299_),
    .A2(_19302_),
    .B1(_01106_),
    .Y(_19303_));
 sky130_fd_sc_hd__clkbuf_2 _48190_ (.A(_19295_),
    .X(_19304_));
 sky130_fd_sc_hd__o211a_1 _48191_ (.A1(_19298_),
    .A2(_19304_),
    .B1(_01106_),
    .C1(_19299_),
    .X(_19305_));
 sky130_fd_sc_hd__a21boi_1 _48192_ (.A1(_18514_),
    .A2(_22248_),
    .B1_N(_18511_),
    .Y(_19306_));
 sky130_fd_sc_hd__o21bai_1 _48193_ (.A1(_19303_),
    .A2(_19305_),
    .B1_N(_19306_),
    .Y(_19307_));
 sky130_fd_sc_hd__a21o_1 _48194_ (.A1(_19299_),
    .A2(_19302_),
    .B1(_01106_),
    .X(_19308_));
 sky130_fd_sc_hd__nand3b_1 _48195_ (.A_N(_19305_),
    .B(_19306_),
    .C(_19308_),
    .Y(_19309_));
 sky130_fd_sc_hd__nand3_1 _48196_ (.A(_19307_),
    .B(_19309_),
    .C(_22259_),
    .Y(_19310_));
 sky130_fd_sc_hd__a21o_1 _48197_ (.A1(_19307_),
    .A2(_19309_),
    .B1(_22248_),
    .X(_19311_));
 sky130_fd_sc_hd__nand2_1 _48198_ (.A(_19310_),
    .B(_19311_),
    .Y(_19312_));
 sky130_fd_sc_hd__and3_1 _48199_ (.A(_18519_),
    .B(_18522_),
    .C(_19312_),
    .X(_19313_));
 sky130_fd_sc_hd__a21oi_1 _48200_ (.A1(_18519_),
    .A2(_18522_),
    .B1(_19312_),
    .Y(_19314_));
 sky130_fd_sc_hd__nor2_1 _48201_ (.A(_19313_),
    .B(_19314_),
    .Y(_19315_));
 sky130_fd_sc_hd__xor2_2 _48202_ (.A(_18520_),
    .B(_19315_),
    .X(_19316_));
 sky130_fd_sc_hd__or3b_2 _48203_ (.A(_19293_),
    .B(_19294_),
    .C_N(_19316_),
    .X(_19317_));
 sky130_fd_sc_hd__o21bai_2 _48204_ (.A1(_19293_),
    .A2(_19294_),
    .B1_N(_19316_),
    .Y(_19318_));
 sky130_fd_sc_hd__nand4_2 _48205_ (.A(_18507_),
    .B(_18526_),
    .C(_19317_),
    .D(_19318_),
    .Y(_19319_));
 sky130_fd_sc_hd__inv_2 _48206_ (.A(_19319_),
    .Y(_19320_));
 sky130_fd_sc_hd__a22oi_4 _48207_ (.A1(_18507_),
    .A2(_18526_),
    .B1(_19317_),
    .B2(_19318_),
    .Y(_19321_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48208_ (.A(\delay_line[29][4] ),
    .X(_19322_));
 sky130_fd_sc_hd__clkbuf_2 _48209_ (.A(_19322_),
    .X(_19323_));
 sky130_fd_sc_hd__nor2_1 _48210_ (.A(_01051_),
    .B(_19323_),
    .Y(_19324_));
 sky130_fd_sc_hd__and2_1 _48211_ (.A(_01051_),
    .B(_19323_),
    .X(_19325_));
 sky130_fd_sc_hd__nor2_1 _48212_ (.A(_18457_),
    .B(_18458_),
    .Y(_19326_));
 sky130_fd_sc_hd__inv_2 _48213_ (.A(_22281_),
    .Y(_19327_));
 sky130_fd_sc_hd__inv_2 _48214_ (.A(\delay_line[30][6] ),
    .Y(_19328_));
 sky130_fd_sc_hd__or2b_1 _48215_ (.A(net320),
    .B_N(_06293_),
    .X(_19329_));
 sky130_fd_sc_hd__or2b_1 _48216_ (.A(_06293_),
    .B_N(net320),
    .X(_19330_));
 sky130_fd_sc_hd__nand3_1 _48217_ (.A(_19328_),
    .B(_19329_),
    .C(_19330_),
    .Y(_19331_));
 sky130_fd_sc_hd__nor2b_2 _48218_ (.A(net320),
    .B_N(\delay_line[30][3] ),
    .Y(_19332_));
 sky130_fd_sc_hd__and2b_1 _48219_ (.A_N(\delay_line[30][3] ),
    .B(\delay_line[30][1] ),
    .X(_19333_));
 sky130_fd_sc_hd__clkbuf_2 _48220_ (.A(_19333_),
    .X(_19334_));
 sky130_fd_sc_hd__buf_1 _48221_ (.A(\delay_line[30][6] ),
    .X(_19335_));
 sky130_fd_sc_hd__buf_2 _48222_ (.A(_19335_),
    .X(_19336_));
 sky130_fd_sc_hd__o21ai_1 _48223_ (.A1(_19332_),
    .A2(_19334_),
    .B1(_19336_),
    .Y(_19337_));
 sky130_fd_sc_hd__o2111ai_1 _48224_ (.A1(_18455_),
    .A2(_18456_),
    .B1(_18452_),
    .C1(_19331_),
    .D1(_19337_),
    .Y(_19338_));
 sky130_fd_sc_hd__a21o_1 _48225_ (.A1(_19331_),
    .A2(_19337_),
    .B1(_18458_),
    .X(_19339_));
 sky130_fd_sc_hd__or4bb_1 _48226_ (.A(_19327_),
    .B(_01029_),
    .C_N(_19338_),
    .D_N(_19339_),
    .X(_19340_));
 sky130_fd_sc_hd__o2bb2a_1 _48227_ (.A1_N(_19338_),
    .A2_N(_19339_),
    .B1(_19327_),
    .B2(_01029_),
    .X(_19341_));
 sky130_fd_sc_hd__inv_2 _48228_ (.A(_19341_),
    .Y(_19342_));
 sky130_fd_sc_hd__a32o_1 _48229_ (.A1(_24622_),
    .A2(_15580_),
    .A3(_19326_),
    .B1(_19340_),
    .B2(_19342_),
    .X(_19343_));
 sky130_fd_sc_hd__nand4_1 _48230_ (.A(_19342_),
    .B(_19326_),
    .C(_15602_),
    .D(_19340_),
    .Y(_19344_));
 sky130_fd_sc_hd__nand4_1 _48231_ (.A(_19343_),
    .B(_19326_),
    .C(_15613_),
    .D(_19344_),
    .Y(_19345_));
 sky130_fd_sc_hd__buf_1 _48232_ (.A(_19345_),
    .X(_19346_));
 sky130_fd_sc_hd__buf_1 _48233_ (.A(_19344_),
    .X(_19347_));
 sky130_fd_sc_hd__a22o_1 _48234_ (.A1(_15624_),
    .A2(_19326_),
    .B1(_19347_),
    .B2(_19343_),
    .X(_19348_));
 sky130_fd_sc_hd__and4bb_4 _48235_ (.A_N(_19324_),
    .B_N(_19325_),
    .C(_19346_),
    .D(_19348_),
    .X(_19349_));
 sky130_fd_sc_hd__a2bb2oi_1 _48236_ (.A1_N(_19324_),
    .A2_N(_19325_),
    .B1(_19346_),
    .B2(_19348_),
    .Y(_19350_));
 sky130_fd_sc_hd__buf_1 _48237_ (.A(\delay_line[31][6] ),
    .X(_19351_));
 sky130_fd_sc_hd__nor2_1 _48238_ (.A(_18465_),
    .B(_19351_),
    .Y(_19352_));
 sky130_fd_sc_hd__nand2_1 _48239_ (.A(_18465_),
    .B(_19351_),
    .Y(_19353_));
 sky130_fd_sc_hd__nand3b_1 _48240_ (.A_N(_19352_),
    .B(_19353_),
    .C(_15789_),
    .Y(_19354_));
 sky130_fd_sc_hd__and2_1 _48241_ (.A(\delay_line[31][5] ),
    .B(_19351_),
    .X(_19355_));
 sky130_fd_sc_hd__inv_2 _48242_ (.A(\delay_line[31][4] ),
    .Y(_19356_));
 sky130_fd_sc_hd__o21ai_1 _48243_ (.A1(_19352_),
    .A2(_19355_),
    .B1(_19356_),
    .Y(_19357_));
 sky130_fd_sc_hd__o21ai_1 _48244_ (.A1(_06249_),
    .A2(_18466_),
    .B1(_18467_),
    .Y(_19358_));
 sky130_fd_sc_hd__a21o_1 _48245_ (.A1(_19354_),
    .A2(_19357_),
    .B1(_19358_),
    .X(_19359_));
 sky130_fd_sc_hd__nand3_1 _48246_ (.A(_19354_),
    .B(_19357_),
    .C(_19358_),
    .Y(_19360_));
 sky130_fd_sc_hd__nand3_1 _48247_ (.A(_19359_),
    .B(_18472_),
    .C(_19360_),
    .Y(_19361_));
 sky130_fd_sc_hd__o21a_1 _48248_ (.A1(_15701_),
    .A2(_15778_),
    .B1(_15800_),
    .X(_19362_));
 sky130_fd_sc_hd__a21oi_1 _48249_ (.A1(_19354_),
    .A2(_19357_),
    .B1(_19358_),
    .Y(_19363_));
 sky130_fd_sc_hd__and3_1 _48250_ (.A(_19354_),
    .B(_19357_),
    .C(_19358_),
    .X(_19364_));
 sky130_fd_sc_hd__o22ai_2 _48251_ (.A1(_19362_),
    .A2(_18473_),
    .B1(_19363_),
    .B2(_19364_),
    .Y(_19365_));
 sky130_fd_sc_hd__a21oi_1 _48252_ (.A1(_19361_),
    .A2(_19365_),
    .B1(_22215_),
    .Y(_19366_));
 sky130_fd_sc_hd__nand3_1 _48253_ (.A(_19365_),
    .B(\delay_line[31][0] ),
    .C(_19361_),
    .Y(_19367_));
 sky130_fd_sc_hd__nand4b_1 _48254_ (.A_N(_19366_),
    .B(_18475_),
    .C(_15855_),
    .D(_19367_),
    .Y(_19368_));
 sky130_fd_sc_hd__buf_1 _48255_ (.A(_19368_),
    .X(_19369_));
 sky130_fd_sc_hd__and3_1 _48256_ (.A(_19365_),
    .B(_22215_),
    .C(_19361_),
    .X(_19370_));
 sky130_fd_sc_hd__o2bb2ai_1 _48257_ (.A1_N(_15866_),
    .A2_N(_18475_),
    .B1(_19370_),
    .B2(_19366_),
    .Y(_19371_));
 sky130_fd_sc_hd__a32o_1 _48258_ (.A1(_15756_),
    .A2(_18476_),
    .A3(_18475_),
    .B1(_19369_),
    .B2(_19371_),
    .X(_19372_));
 sky130_fd_sc_hd__and3_1 _48259_ (.A(_15756_),
    .B(_18476_),
    .C(_18475_),
    .X(_19373_));
 sky130_fd_sc_hd__nand3_1 _48260_ (.A(_19371_),
    .B(_19373_),
    .C(_19368_),
    .Y(_19374_));
 sky130_fd_sc_hd__buf_1 _48261_ (.A(_19374_),
    .X(_19375_));
 sky130_fd_sc_hd__and3_1 _48262_ (.A(_19372_),
    .B(_19375_),
    .C(_18481_),
    .X(_19376_));
 sky130_fd_sc_hd__a21oi_1 _48263_ (.A1(_19372_),
    .A2(_19375_),
    .B1(_18481_),
    .Y(_19377_));
 sky130_fd_sc_hd__o22a_1 _48264_ (.A1(_19349_),
    .A2(_19350_),
    .B1(_19376_),
    .B2(_19377_),
    .X(_19378_));
 sky130_fd_sc_hd__nor4_2 _48265_ (.A(_19349_),
    .B(_19350_),
    .C(_19376_),
    .D(_19377_),
    .Y(_19379_));
 sky130_fd_sc_hd__nor4_2 _48266_ (.A(_19320_),
    .B(_19321_),
    .C(_19378_),
    .D(_19379_),
    .Y(_19380_));
 sky130_fd_sc_hd__o22a_1 _48267_ (.A1(_19320_),
    .A2(_19321_),
    .B1(_19378_),
    .B2(_19379_),
    .X(_19381_));
 sky130_fd_sc_hd__nor2_2 _48268_ (.A(_19380_),
    .B(_19381_),
    .Y(_19382_));
 sky130_fd_sc_hd__or3_1 _48269_ (.A(_19262_),
    .B(_18341_),
    .C(_19382_),
    .X(_19383_));
 sky130_fd_sc_hd__o21ai_2 _48270_ (.A1(_19262_),
    .A2(_18341_),
    .B1(_19382_),
    .Y(_19384_));
 sky130_fd_sc_hd__and2_1 _48271_ (.A(_19383_),
    .B(_19384_),
    .X(_19385_));
 sky130_fd_sc_hd__a31o_1 _48272_ (.A1(_18527_),
    .A2(_18525_),
    .A3(_18526_),
    .B1(_19385_),
    .X(_19386_));
 sky130_fd_sc_hd__o21ai_2 _48273_ (.A1(_18529_),
    .A2(net120),
    .B1(_19385_),
    .Y(_19387_));
 sky130_fd_sc_hd__o21a_2 _48274_ (.A1(net121),
    .A2(_19386_),
    .B1(_19387_),
    .X(_19388_));
 sky130_fd_sc_hd__a21boi_2 _48275_ (.A1(_18396_),
    .A2(_18438_),
    .B1_N(_18439_),
    .Y(_19389_));
 sky130_fd_sc_hd__clkbuf_2 _48276_ (.A(\delay_line[18][5] ),
    .X(_19390_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48277_ (.A(_19390_),
    .X(_19391_));
 sky130_fd_sc_hd__nor2_1 _48278_ (.A(_01666_),
    .B(_19391_),
    .Y(_19392_));
 sky130_fd_sc_hd__inv_2 _48279_ (.A(net375),
    .Y(_19393_));
 sky130_fd_sc_hd__inv_2 _48280_ (.A(\delay_line[18][5] ),
    .Y(_19394_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48281_ (.A(_19394_),
    .X(_19395_));
 sky130_fd_sc_hd__nor2_1 _48282_ (.A(_19393_),
    .B(_19395_),
    .Y(_19396_));
 sky130_fd_sc_hd__buf_1 _48283_ (.A(_19396_),
    .X(_19397_));
 sky130_fd_sc_hd__a2bb2o_1 _48284_ (.A1_N(_19392_),
    .A2_N(_19397_),
    .B1(_23863_),
    .B2(_18385_),
    .X(_19398_));
 sky130_fd_sc_hd__or4_2 _48285_ (.A(_23951_),
    .B(_18389_),
    .C(_19392_),
    .D(_19397_),
    .X(_19399_));
 sky130_fd_sc_hd__clkbuf_2 _48286_ (.A(_18370_),
    .X(_19400_));
 sky130_fd_sc_hd__and2_2 _48287_ (.A(net371),
    .B(\delay_line[19][5] ),
    .X(_19401_));
 sky130_fd_sc_hd__clkbuf_2 _48288_ (.A(\delay_line[19][5] ),
    .X(_19402_));
 sky130_fd_sc_hd__nor2_1 _48289_ (.A(_18374_),
    .B(_19402_),
    .Y(_19403_));
 sky130_fd_sc_hd__o2bb2ai_2 _48290_ (.A1_N(_18367_),
    .A2_N(_18374_),
    .B1(_19401_),
    .B2(_19403_),
    .Y(_19404_));
 sky130_fd_sc_hd__inv_2 _48291_ (.A(\delay_line[19][5] ),
    .Y(_19405_));
 sky130_fd_sc_hd__nand3_2 _48292_ (.A(_19405_),
    .B(_18374_),
    .C(_16382_),
    .Y(_19406_));
 sky130_fd_sc_hd__a21o_1 _48293_ (.A1(_19404_),
    .A2(_19406_),
    .B1(_23874_),
    .X(_19407_));
 sky130_fd_sc_hd__nand3_1 _48294_ (.A(_19404_),
    .B(_19406_),
    .C(_23874_),
    .Y(_19408_));
 sky130_fd_sc_hd__and4_1 _48295_ (.A(_19400_),
    .B(_19407_),
    .C(_19408_),
    .D(_18377_),
    .X(_19409_));
 sky130_fd_sc_hd__nand2_1 _48296_ (.A(_18367_),
    .B(_07393_),
    .Y(_19410_));
 sky130_fd_sc_hd__o2bb2a_1 _48297_ (.A1_N(_19407_),
    .A2_N(_19408_),
    .B1(_18376_),
    .B2(_19410_),
    .X(_19411_));
 sky130_fd_sc_hd__nor2_2 _48298_ (.A(_19409_),
    .B(_19411_),
    .Y(_19412_));
 sky130_fd_sc_hd__or3_2 _48299_ (.A(_18379_),
    .B(_18381_),
    .C(_19412_),
    .X(_19413_));
 sky130_fd_sc_hd__o21ai_2 _48300_ (.A1(_18379_),
    .A2(_18381_),
    .B1(_19412_),
    .Y(_19414_));
 sky130_fd_sc_hd__nand4_4 _48301_ (.A(_19398_),
    .B(_19399_),
    .C(_19413_),
    .D(_19414_),
    .Y(_19415_));
 sky130_fd_sc_hd__a22o_2 _48302_ (.A1(_19398_),
    .A2(_19399_),
    .B1(_19413_),
    .B2(_19414_),
    .X(_19416_));
 sky130_fd_sc_hd__buf_1 _48303_ (.A(\delay_line[21][5] ),
    .X(_19417_));
 sky130_fd_sc_hd__nor2_1 _48304_ (.A(net360),
    .B(_19417_),
    .Y(_19418_));
 sky130_fd_sc_hd__and2_1 _48305_ (.A(net360),
    .B(_19417_),
    .X(_19419_));
 sky130_fd_sc_hd__o2bb2ai_2 _48306_ (.A1_N(_18345_),
    .A2_N(_18347_),
    .B1(_19418_),
    .B2(_19419_),
    .Y(_19420_));
 sky130_fd_sc_hd__nand3b_2 _48307_ (.A_N(_19417_),
    .B(_18347_),
    .C(_18345_),
    .Y(_19421_));
 sky130_fd_sc_hd__a21o_1 _48308_ (.A1(_19420_),
    .A2(_19421_),
    .B1(_23995_),
    .X(_19422_));
 sky130_fd_sc_hd__nand3_1 _48309_ (.A(_19420_),
    .B(_19421_),
    .C(_23984_),
    .Y(_19423_));
 sky130_fd_sc_hd__or4bb_2 _48310_ (.A(_18349_),
    .B(_18360_),
    .C_N(_19422_),
    .D_N(_19423_),
    .X(_19424_));
 sky130_fd_sc_hd__a2bb2o_1 _48311_ (.A1_N(_18360_),
    .A2_N(_18349_),
    .B1(_19423_),
    .B2(_19422_),
    .X(_19425_));
 sky130_fd_sc_hd__a22oi_1 _48312_ (.A1(_18355_),
    .A2(_18366_),
    .B1(_19424_),
    .B2(_19425_),
    .Y(_19426_));
 sky130_fd_sc_hd__and4_1 _48313_ (.A(_18355_),
    .B(_18366_),
    .C(_19424_),
    .D(_19425_),
    .X(_19427_));
 sky130_fd_sc_hd__nor2_1 _48314_ (.A(_19426_),
    .B(_19427_),
    .Y(_19428_));
 sky130_fd_sc_hd__a21boi_1 _48315_ (.A1(_19415_),
    .A2(_19416_),
    .B1_N(_19428_),
    .Y(_19429_));
 sky130_fd_sc_hd__nand3b_4 _48316_ (.A_N(_19428_),
    .B(_19415_),
    .C(_19416_),
    .Y(_19430_));
 sky130_fd_sc_hd__inv_2 _48317_ (.A(_19430_),
    .Y(_19431_));
 sky130_fd_sc_hd__and2_1 _48318_ (.A(\delay_line[16][1] ),
    .B(\delay_line[16][2] ),
    .X(_19432_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48319_ (.A(_19432_),
    .X(_19433_));
 sky130_fd_sc_hd__o21ai_1 _48320_ (.A1(_01864_),
    .A2(_07206_),
    .B1(\delay_line[16][0] ),
    .Y(_19434_));
 sky130_fd_sc_hd__clkbuf_2 _48321_ (.A(\delay_line[16][5] ),
    .X(_19435_));
 sky130_fd_sc_hd__nor2_1 _48322_ (.A(\delay_line[16][1] ),
    .B(\delay_line[16][2] ),
    .Y(_19436_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48323_ (.A(_19436_),
    .X(_19437_));
 sky130_fd_sc_hd__o21ai_1 _48324_ (.A1(_19433_),
    .A2(_19437_),
    .B1(_16634_),
    .Y(_19438_));
 sky130_fd_sc_hd__o211a_1 _48325_ (.A1(_19433_),
    .A2(_19434_),
    .B1(_19435_),
    .C1(_19438_),
    .X(_19439_));
 sky130_fd_sc_hd__or3_1 _48326_ (.A(_19437_),
    .B(_16634_),
    .C(_19433_),
    .X(_19440_));
 sky130_fd_sc_hd__clkbuf_2 _48327_ (.A(_19435_),
    .X(_19441_));
 sky130_fd_sc_hd__a21oi_1 _48328_ (.A1(_19440_),
    .A2(_19438_),
    .B1(_19441_),
    .Y(_19442_));
 sky130_fd_sc_hd__a211oi_1 _48329_ (.A1(_18398_),
    .A2(_18401_),
    .B1(_19439_),
    .C1(_19442_),
    .Y(_19443_));
 sky130_fd_sc_hd__o211a_1 _48330_ (.A1(_19439_),
    .A2(_19442_),
    .B1(_18398_),
    .C1(_18401_),
    .X(_19444_));
 sky130_fd_sc_hd__nor3_2 _48331_ (.A(_19443_),
    .B(_18404_),
    .C(_19444_),
    .Y(_19445_));
 sky130_fd_sc_hd__clkbuf_2 _48332_ (.A(_19443_),
    .X(_19446_));
 sky130_fd_sc_hd__o21a_1 _48333_ (.A1(_19444_),
    .A2(_19446_),
    .B1(_18404_),
    .X(_19447_));
 sky130_fd_sc_hd__nor2_1 _48334_ (.A(\delay_line[14][0] ),
    .B(_01765_),
    .Y(_19448_));
 sky130_fd_sc_hd__and2_2 _48335_ (.A(net394),
    .B(net393),
    .X(_19449_));
 sky130_fd_sc_hd__buf_1 _48336_ (.A(\delay_line[14][5] ),
    .X(_19450_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48337_ (.A(_19450_),
    .X(_19451_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48338_ (.A(_19451_),
    .X(_19452_));
 sky130_fd_sc_hd__or3b_1 _48339_ (.A(_19448_),
    .B(_19449_),
    .C_N(_19452_),
    .X(_19453_));
 sky130_fd_sc_hd__o21bai_1 _48340_ (.A1(_19448_),
    .A2(_19449_),
    .B1_N(_19452_),
    .Y(_19454_));
 sky130_fd_sc_hd__nand4_2 _48341_ (.A(_19453_),
    .B(_19454_),
    .C(_24061_),
    .D(_18407_),
    .Y(_19455_));
 sky130_fd_sc_hd__a22o_1 _48342_ (.A1(_24072_),
    .A2(_18408_),
    .B1(_19453_),
    .B2(_19454_),
    .X(_19456_));
 sky130_fd_sc_hd__nand2_1 _48343_ (.A(_19455_),
    .B(_19456_),
    .Y(_19457_));
 sky130_fd_sc_hd__and2_1 _48344_ (.A(net387),
    .B(\delay_line[15][6] ),
    .X(_19458_));
 sky130_fd_sc_hd__nor2_1 _48345_ (.A(net387),
    .B(\delay_line[15][6] ),
    .Y(_19459_));
 sky130_fd_sc_hd__o21bai_2 _48346_ (.A1(_19458_),
    .A2(_19459_),
    .B1_N(_18415_),
    .Y(_19460_));
 sky130_fd_sc_hd__clkbuf_2 _48347_ (.A(\delay_line[15][6] ),
    .X(_19461_));
 sky130_fd_sc_hd__nand2_1 _48348_ (.A(\delay_line[15][4] ),
    .B(_19461_),
    .Y(_19462_));
 sky130_fd_sc_hd__nand3b_1 _48349_ (.A_N(_19459_),
    .B(_18415_),
    .C(_19462_),
    .Y(_19463_));
 sky130_fd_sc_hd__and3_1 _48350_ (.A(_19460_),
    .B(_24083_),
    .C(_19463_),
    .X(_19464_));
 sky130_fd_sc_hd__inv_2 _48351_ (.A(_19464_),
    .Y(_19465_));
 sky130_fd_sc_hd__a21o_1 _48352_ (.A1(_19463_),
    .A2(_19460_),
    .B1(_24083_),
    .X(_19466_));
 sky130_fd_sc_hd__clkbuf_2 _48353_ (.A(_18422_),
    .X(_19467_));
 sky130_fd_sc_hd__a21oi_2 _48354_ (.A1(_16788_),
    .A2(_19467_),
    .B1(_18417_),
    .Y(_19468_));
 sky130_fd_sc_hd__a211o_1 _48355_ (.A1(_19465_),
    .A2(_19466_),
    .B1(_19468_),
    .C1(_18421_),
    .X(_19469_));
 sky130_fd_sc_hd__o211ai_4 _48356_ (.A1(_19468_),
    .A2(_18421_),
    .B1(_19465_),
    .C1(_19466_),
    .Y(_19470_));
 sky130_fd_sc_hd__nand2_1 _48357_ (.A(_19469_),
    .B(_19470_),
    .Y(_19471_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48358_ (.A(_19471_),
    .X(_19472_));
 sky130_fd_sc_hd__o31a_1 _48359_ (.A1(_18413_),
    .A2(_07151_),
    .A3(_18426_),
    .B1(_18431_),
    .X(_19473_));
 sky130_fd_sc_hd__xnor2_1 _48360_ (.A(_19472_),
    .B(_19473_),
    .Y(_19474_));
 sky130_fd_sc_hd__nor2_2 _48361_ (.A(_19457_),
    .B(_19474_),
    .Y(_19475_));
 sky130_fd_sc_hd__and2_1 _48362_ (.A(_19457_),
    .B(_19474_),
    .X(_19476_));
 sky130_fd_sc_hd__nor2_1 _48363_ (.A(_19475_),
    .B(_19476_),
    .Y(_19477_));
 sky130_fd_sc_hd__nor3b_2 _48364_ (.A(_19445_),
    .B(_19447_),
    .C_N(_19477_),
    .Y(_19478_));
 sky130_fd_sc_hd__o21ba_1 _48365_ (.A1(_19445_),
    .A2(_19447_),
    .B1_N(_19477_),
    .X(_19479_));
 sky130_fd_sc_hd__nand4_1 _48366_ (.A(_18403_),
    .B(_18404_),
    .C(_18433_),
    .D(_18434_),
    .Y(_19480_));
 sky130_fd_sc_hd__o211a_2 _48367_ (.A1(_19478_),
    .A2(_19479_),
    .B1(_18433_),
    .C1(_19480_),
    .X(_19481_));
 sky130_fd_sc_hd__a211o_2 _48368_ (.A1(_18433_),
    .A2(_19480_),
    .B1(_19478_),
    .C1(_19479_),
    .X(_19482_));
 sky130_fd_sc_hd__inv_2 _48369_ (.A(_19482_),
    .Y(_19483_));
 sky130_fd_sc_hd__nor4_2 _48370_ (.A(_19429_),
    .B(_19431_),
    .C(_19481_),
    .D(_19483_),
    .Y(_19484_));
 sky130_fd_sc_hd__o22a_1 _48371_ (.A1(_19429_),
    .A2(_19431_),
    .B1(_19481_),
    .B2(_19483_),
    .X(_19485_));
 sky130_fd_sc_hd__nor3_4 _48372_ (.A(_19389_),
    .B(_19484_),
    .C(_19485_),
    .Y(_19486_));
 sky130_fd_sc_hd__and2_1 _48373_ (.A(\delay_line[25][4] ),
    .B(\delay_line[25][6] ),
    .X(_19487_));
 sky130_fd_sc_hd__clkbuf_2 _48374_ (.A(\delay_line[25][6] ),
    .X(_19488_));
 sky130_fd_sc_hd__nor2_1 _48375_ (.A(\delay_line[25][4] ),
    .B(_19488_),
    .Y(_19489_));
 sky130_fd_sc_hd__o21bai_2 _48376_ (.A1(_19487_),
    .A2(_19489_),
    .B1_N(_18326_),
    .Y(_19490_));
 sky130_fd_sc_hd__nand2_1 _48377_ (.A(_17204_),
    .B(_19488_),
    .Y(_19491_));
 sky130_fd_sc_hd__nand3b_2 _48378_ (.A_N(_19489_),
    .B(_18326_),
    .C(_19491_),
    .Y(_19492_));
 sky130_fd_sc_hd__and3_2 _48379_ (.A(_19490_),
    .B(_23731_),
    .C(_19492_),
    .X(_19493_));
 sky130_fd_sc_hd__a21oi_2 _48380_ (.A1(_19492_),
    .A2(_19490_),
    .B1(_23742_),
    .Y(_19494_));
 sky130_fd_sc_hd__o211ai_4 _48381_ (.A1(_19493_),
    .A2(_19494_),
    .B1(_18327_),
    .C1(_18331_),
    .Y(_19495_));
 sky130_fd_sc_hd__a211o_2 _48382_ (.A1(_18327_),
    .A2(_18330_),
    .B1(_19493_),
    .C1(_19494_),
    .X(_19496_));
 sky130_fd_sc_hd__nand2_4 _48383_ (.A(_19495_),
    .B(_19496_),
    .Y(_19497_));
 sky130_fd_sc_hd__and4b_1 _48384_ (.A_N(_17215_),
    .B(_18334_),
    .C(_18333_),
    .D(_17161_),
    .X(_19498_));
 sky130_fd_sc_hd__a41o_1 _48385_ (.A1(_17270_),
    .A2(_17193_),
    .A3(_18331_),
    .A4(_18329_),
    .B1(_19498_),
    .X(_19499_));
 sky130_fd_sc_hd__xor2_4 _48386_ (.A(_19497_),
    .B(_19499_),
    .X(_19500_));
 sky130_fd_sc_hd__buf_1 _48387_ (.A(\delay_line[22][5] ),
    .X(_19501_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48388_ (.A(_19501_),
    .X(_19502_));
 sky130_fd_sc_hd__nor2_1 _48389_ (.A(_01402_),
    .B(_19502_),
    .Y(_19503_));
 sky130_fd_sc_hd__and2_1 _48390_ (.A(_01402_),
    .B(_19502_),
    .X(_19504_));
 sky130_fd_sc_hd__o2bb2a_1 _48391_ (.A1_N(_23676_),
    .A2_N(_18318_),
    .B1(_19503_),
    .B2(_19504_),
    .X(_19505_));
 sky130_fd_sc_hd__and4bb_1 _48392_ (.A_N(_19503_),
    .B_N(_19504_),
    .C(_23666_),
    .D(_18316_),
    .X(_19506_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48393_ (.A(_19506_),
    .X(_19507_));
 sky130_fd_sc_hd__clkbuf_2 _48394_ (.A(_18306_),
    .X(_19508_));
 sky130_fd_sc_hd__and2_1 _48395_ (.A(net345),
    .B(net344),
    .X(_19509_));
 sky130_fd_sc_hd__clkbuf_2 _48396_ (.A(_19509_),
    .X(_19510_));
 sky130_fd_sc_hd__o21ai_2 _48397_ (.A1(net345),
    .A2(net344),
    .B1(net346),
    .Y(_19511_));
 sky130_fd_sc_hd__clkbuf_2 _48398_ (.A(\delay_line[24][5] ),
    .X(_19512_));
 sky130_fd_sc_hd__clkbuf_2 _48399_ (.A(_19512_),
    .X(_19513_));
 sky130_fd_sc_hd__nor2_2 _48400_ (.A(net345),
    .B(net344),
    .Y(_19514_));
 sky130_fd_sc_hd__o21ai_1 _48401_ (.A1(_19509_),
    .A2(_19514_),
    .B1(_18304_),
    .Y(_19515_));
 sky130_fd_sc_hd__o211a_1 _48402_ (.A1(_19510_),
    .A2(_19511_),
    .B1(_19513_),
    .C1(_19515_),
    .X(_19516_));
 sky130_fd_sc_hd__buf_2 _48403_ (.A(_19516_),
    .X(_19517_));
 sky130_fd_sc_hd__or3_1 _48404_ (.A(_19514_),
    .B(_18304_),
    .C(_19510_),
    .X(_19518_));
 sky130_fd_sc_hd__clkbuf_2 _48405_ (.A(_19513_),
    .X(_19519_));
 sky130_fd_sc_hd__a21oi_2 _48406_ (.A1(_19518_),
    .A2(_19515_),
    .B1(_19519_),
    .Y(_19520_));
 sky130_fd_sc_hd__o221ai_2 _48407_ (.A1(_18305_),
    .A2(_19508_),
    .B1(_19517_),
    .B2(_19520_),
    .C1(_18313_),
    .Y(_19521_));
 sky130_fd_sc_hd__a211o_1 _48408_ (.A1(_18308_),
    .A2(_18312_),
    .B1(_19517_),
    .C1(_19520_),
    .X(_19522_));
 sky130_fd_sc_hd__and3b_1 _48409_ (.A_N(_18314_),
    .B(_19521_),
    .C(_19522_),
    .X(_19523_));
 sky130_fd_sc_hd__buf_1 _48410_ (.A(_19523_),
    .X(_19524_));
 sky130_fd_sc_hd__a32o_1 _48411_ (.A1(_17062_),
    .A2(_18313_),
    .A3(_18311_),
    .B1(_19521_),
    .B2(_19522_),
    .X(_19525_));
 sky130_fd_sc_hd__or4b_1 _48412_ (.A(_19505_),
    .B(_19507_),
    .C(_19524_),
    .D_N(_19525_),
    .X(_19526_));
 sky130_fd_sc_hd__inv_2 _48413_ (.A(_19524_),
    .Y(_19527_));
 sky130_fd_sc_hd__a2bb2o_1 _48414_ (.A1_N(_19505_),
    .A2_N(_19507_),
    .B1(_19527_),
    .B2(_19525_),
    .X(_19528_));
 sky130_fd_sc_hd__nand2_1 _48415_ (.A(_19526_),
    .B(_19528_),
    .Y(_19529_));
 sky130_fd_sc_hd__xor2_2 _48416_ (.A(_19500_),
    .B(_19529_),
    .X(_19530_));
 sky130_fd_sc_hd__and3_1 _48417_ (.A(_19530_),
    .B(_18394_),
    .C(_18391_),
    .X(_19531_));
 sky130_fd_sc_hd__a21oi_1 _48418_ (.A1(_18391_),
    .A2(_18394_),
    .B1(_19530_),
    .Y(_19532_));
 sky130_fd_sc_hd__nor2_1 _48419_ (.A(_19531_),
    .B(_19532_),
    .Y(_19533_));
 sky130_fd_sc_hd__a31o_2 _48420_ (.A1(_18319_),
    .A2(_18314_),
    .A3(_18315_),
    .B1(_18337_),
    .X(_19534_));
 sky130_fd_sc_hd__xnor2_1 _48421_ (.A(_19533_),
    .B(_19534_),
    .Y(_19535_));
 sky130_fd_sc_hd__o21a_1 _48422_ (.A1(_19484_),
    .A2(_19485_),
    .B1(_19389_),
    .X(_19536_));
 sky130_fd_sc_hd__nor3_1 _48423_ (.A(_19486_),
    .B(_19535_),
    .C(_19536_),
    .Y(_19537_));
 sky130_fd_sc_hd__o21a_1 _48424_ (.A1(_19536_),
    .A2(_19486_),
    .B1(_19535_),
    .X(_19538_));
 sky130_fd_sc_hd__nor2_1 _48425_ (.A(_19537_),
    .B(_19538_),
    .Y(_19539_));
 sky130_fd_sc_hd__a211oi_1 _48426_ (.A1(_18343_),
    .A2(_18445_),
    .B1(_19539_),
    .C1(_18444_),
    .Y(_19540_));
 sky130_fd_sc_hd__o21a_1 _48427_ (.A1(_18444_),
    .A2(_18446_),
    .B1(_19539_),
    .X(_19541_));
 sky130_fd_sc_hd__nor2_1 _48428_ (.A(_19540_),
    .B(_19541_),
    .Y(_19542_));
 sky130_fd_sc_hd__xor2_2 _48429_ (.A(_19388_),
    .B(_19542_),
    .X(_19543_));
 sky130_fd_sc_hd__xor2_1 _48430_ (.A(_19261_),
    .B(_19543_),
    .X(_19544_));
 sky130_fd_sc_hd__a21boi_1 _48431_ (.A1(_18627_),
    .A2(_18699_),
    .B1_N(_18698_),
    .Y(_19545_));
 sky130_fd_sc_hd__a21o_1 _48432_ (.A1(_18629_),
    .A2(_18692_),
    .B1(_18695_),
    .X(_19546_));
 sky130_fd_sc_hd__nor2_1 _48433_ (.A(net138),
    .B(net118),
    .Y(_19547_));
 sky130_fd_sc_hd__buf_1 _48434_ (.A(\delay_line[34][4] ),
    .X(_19548_));
 sky130_fd_sc_hd__buf_1 _48435_ (.A(\delay_line[34][6] ),
    .X(_19549_));
 sky130_fd_sc_hd__nor2_1 _48436_ (.A(_19548_),
    .B(_19549_),
    .Y(_19550_));
 sky130_fd_sc_hd__and2_1 _48437_ (.A(_19548_),
    .B(_19549_),
    .X(_19551_));
 sky130_fd_sc_hd__o21ai_1 _48438_ (.A1(_19550_),
    .A2(_19551_),
    .B1(_18639_),
    .Y(_19552_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48439_ (.A(\delay_line[34][6] ),
    .X(_19553_));
 sky130_fd_sc_hd__nand2_1 _48440_ (.A(_17810_),
    .B(_19553_),
    .Y(_19554_));
 sky130_fd_sc_hd__nand3b_2 _48441_ (.A_N(_19550_),
    .B(_19554_),
    .C(_18632_),
    .Y(_19555_));
 sky130_fd_sc_hd__nor2_1 _48442_ (.A(net307),
    .B(_18630_),
    .Y(_19556_));
 sky130_fd_sc_hd__nand2_1 _48443_ (.A(net307),
    .B(_18630_),
    .Y(_19557_));
 sky130_fd_sc_hd__and2b_1 _48444_ (.A_N(_19556_),
    .B(_19557_),
    .X(_19558_));
 sky130_fd_sc_hd__a21oi_1 _48445_ (.A1(_19552_),
    .A2(_19555_),
    .B1(_19558_),
    .Y(_19559_));
 sky130_fd_sc_hd__and3_1 _48446_ (.A(_19558_),
    .B(_19552_),
    .C(_19555_),
    .X(_19560_));
 sky130_fd_sc_hd__o211ai_2 _48447_ (.A1(_19559_),
    .A2(_19560_),
    .B1(_18640_),
    .C1(_18641_),
    .Y(_19561_));
 sky130_fd_sc_hd__a211o_1 _48448_ (.A1(_18640_),
    .A2(_18641_),
    .B1(_19559_),
    .C1(_19560_),
    .X(_19562_));
 sky130_fd_sc_hd__nand3b_1 _48449_ (.A_N(_18637_),
    .B(_19561_),
    .C(_19562_),
    .Y(_19563_));
 sky130_fd_sc_hd__a21bo_1 _48450_ (.A1(_19561_),
    .A2(_19562_),
    .B1_N(_18637_),
    .X(_19564_));
 sky130_fd_sc_hd__nand4_1 _48451_ (.A(_18645_),
    .B(_18647_),
    .C(_19563_),
    .D(_19564_),
    .Y(_19565_));
 sky130_fd_sc_hd__a22o_1 _48452_ (.A1(_18645_),
    .A2(_18647_),
    .B1(_19563_),
    .B2(_19564_),
    .X(_19566_));
 sky130_fd_sc_hd__nand2_1 _48453_ (.A(_19565_),
    .B(_19566_),
    .Y(_19567_));
 sky130_fd_sc_hd__xor2_1 _48454_ (.A(_18648_),
    .B(_19567_),
    .X(_19568_));
 sky130_fd_sc_hd__inv_2 _48455_ (.A(_18657_),
    .Y(_19569_));
 sky130_fd_sc_hd__buf_1 _48456_ (.A(net314),
    .X(_19570_));
 sky130_fd_sc_hd__nor2_1 _48457_ (.A(_18652_),
    .B(_19570_),
    .Y(_19571_));
 sky130_fd_sc_hd__and2_1 _48458_ (.A(_18652_),
    .B(_02150_),
    .X(_19572_));
 sky130_fd_sc_hd__inv_2 _48459_ (.A(\delay_line[33][6] ),
    .Y(_19573_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48460_ (.A(_19573_),
    .X(_19574_));
 sky130_fd_sc_hd__o21ai_1 _48461_ (.A1(_19571_),
    .A2(_19572_),
    .B1(_19574_),
    .Y(_19575_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48462_ (.A(\delay_line[33][6] ),
    .X(_19576_));
 sky130_fd_sc_hd__o21ai_1 _48463_ (.A1(_18652_),
    .A2(net314),
    .B1(_19576_),
    .Y(_19577_));
 sky130_fd_sc_hd__a21o_1 _48464_ (.A1(_00557_),
    .A2(_02150_),
    .B1(_19577_),
    .X(_19578_));
 sky130_fd_sc_hd__and3_1 _48465_ (.A(_18656_),
    .B(_19575_),
    .C(_19578_),
    .X(_19579_));
 sky130_fd_sc_hd__a21o_1 _48466_ (.A1(_19575_),
    .A2(_19578_),
    .B1(_18656_),
    .X(_19580_));
 sky130_fd_sc_hd__and2b_1 _48467_ (.A_N(_19579_),
    .B(_19580_),
    .X(_19581_));
 sky130_fd_sc_hd__xor2_1 _48468_ (.A(_18653_),
    .B(_19581_),
    .X(_19582_));
 sky130_fd_sc_hd__nor2_1 _48469_ (.A(_19569_),
    .B(_19582_),
    .Y(_19583_));
 sky130_fd_sc_hd__and2_1 _48470_ (.A(_19569_),
    .B(_19582_),
    .X(_19584_));
 sky130_fd_sc_hd__nor2_1 _48471_ (.A(_19583_),
    .B(_19584_),
    .Y(_19585_));
 sky130_fd_sc_hd__nor2_2 _48472_ (.A(\delay_line[32][5] ),
    .B(\delay_line[32][6] ),
    .Y(_19586_));
 sky130_fd_sc_hd__and2_1 _48473_ (.A(\delay_line[32][5] ),
    .B(\delay_line[32][6] ),
    .X(_19587_));
 sky130_fd_sc_hd__o21ai_2 _48474_ (.A1(_19586_),
    .A2(_19587_),
    .B1(_18671_),
    .Y(_19588_));
 sky130_fd_sc_hd__buf_1 _48475_ (.A(\delay_line[32][6] ),
    .X(_19589_));
 sky130_fd_sc_hd__nand2_1 _48476_ (.A(_18663_),
    .B(_19589_),
    .Y(_19590_));
 sky130_fd_sc_hd__nand3b_2 _48477_ (.A_N(_19586_),
    .B(_19590_),
    .C(_17831_),
    .Y(_19591_));
 sky130_fd_sc_hd__o21ai_2 _48478_ (.A1(_05238_),
    .A2(_18664_),
    .B1(_18665_),
    .Y(_19592_));
 sky130_fd_sc_hd__a21oi_2 _48479_ (.A1(_19588_),
    .A2(_19591_),
    .B1(_19592_),
    .Y(_19593_));
 sky130_fd_sc_hd__inv_2 _48480_ (.A(_19593_),
    .Y(_19594_));
 sky130_fd_sc_hd__nand3_1 _48481_ (.A(_19592_),
    .B(_19588_),
    .C(_19591_),
    .Y(_19595_));
 sky130_fd_sc_hd__nand3_1 _48482_ (.A(_05271_),
    .B(_19594_),
    .C(_19595_),
    .Y(_19596_));
 sky130_fd_sc_hd__o21a_1 _48483_ (.A1(_05216_),
    .A2(_18674_),
    .B1(_18676_),
    .X(_19597_));
 sky130_fd_sc_hd__and3_1 _48484_ (.A(_19592_),
    .B(_19588_),
    .C(_19591_),
    .X(_19598_));
 sky130_fd_sc_hd__o21ai_1 _48485_ (.A1(_19593_),
    .A2(_19598_),
    .B1(_05315_),
    .Y(_19599_));
 sky130_fd_sc_hd__nand3_1 _48486_ (.A(_19596_),
    .B(_19597_),
    .C(_19599_),
    .Y(_19600_));
 sky130_fd_sc_hd__o21ai_1 _48487_ (.A1(_05216_),
    .A2(_18674_),
    .B1(_18676_),
    .Y(_19601_));
 sky130_fd_sc_hd__nand3_1 _48488_ (.A(_19594_),
    .B(_19595_),
    .C(_05315_),
    .Y(_19602_));
 sky130_fd_sc_hd__o21ai_1 _48489_ (.A1(_19593_),
    .A2(_19598_),
    .B1(_05260_),
    .Y(_19603_));
 sky130_fd_sc_hd__nand3_1 _48490_ (.A(_19601_),
    .B(_19602_),
    .C(_19603_),
    .Y(_19604_));
 sky130_fd_sc_hd__nand3_1 _48491_ (.A(_19600_),
    .B(_19604_),
    .C(_22556_),
    .Y(_19605_));
 sky130_fd_sc_hd__buf_1 _48492_ (.A(_19604_),
    .X(_19606_));
 sky130_fd_sc_hd__a21o_1 _48493_ (.A1(_19600_),
    .A2(_19606_),
    .B1(_22556_),
    .X(_19607_));
 sky130_fd_sc_hd__a2bb2o_2 _48494_ (.A1_N(_18679_),
    .A2_N(_18678_),
    .B1(_19605_),
    .B2(_19607_),
    .X(_19608_));
 sky130_fd_sc_hd__nor2_1 _48495_ (.A(_18685_),
    .B(_18682_),
    .Y(_19609_));
 sky130_fd_sc_hd__buf_2 _48496_ (.A(_19609_),
    .X(_19610_));
 sky130_fd_sc_hd__buf_2 _48497_ (.A(_18672_),
    .X(_19611_));
 sky130_fd_sc_hd__and4b_1 _48498_ (.A_N(_18661_),
    .B(_18680_),
    .C(_18681_),
    .D(_19611_),
    .X(_19612_));
 sky130_fd_sc_hd__inv_2 _48499_ (.A(_18681_),
    .Y(_19613_));
 sky130_fd_sc_hd__and3_1 _48500_ (.A(_19600_),
    .B(_19606_),
    .C(_22556_),
    .X(_19614_));
 sky130_fd_sc_hd__a21oi_1 _48501_ (.A1(_19600_),
    .A2(_19606_),
    .B1(_22556_),
    .Y(_19615_));
 sky130_fd_sc_hd__nor2_2 _48502_ (.A(_19614_),
    .B(_19615_),
    .Y(_19616_));
 sky130_fd_sc_hd__o21ai_2 _48503_ (.A1(_19613_),
    .A2(_19609_),
    .B1(_19616_),
    .Y(_19617_));
 sky130_fd_sc_hd__o211a_1 _48504_ (.A1(_19608_),
    .A2(_19610_),
    .B1(_19612_),
    .C1(_19617_),
    .X(_19618_));
 sky130_fd_sc_hd__o21ai_1 _48505_ (.A1(_19610_),
    .A2(_19608_),
    .B1(_19617_),
    .Y(_19619_));
 sky130_fd_sc_hd__o31a_1 _48506_ (.A1(_18660_),
    .A2(_18661_),
    .A3(_18683_),
    .B1(_19619_),
    .X(_19620_));
 sky130_fd_sc_hd__nor2_1 _48507_ (.A(_19618_),
    .B(_19620_),
    .Y(_19621_));
 sky130_fd_sc_hd__xnor2_1 _48508_ (.A(_19585_),
    .B(_19621_),
    .Y(_19622_));
 sky130_fd_sc_hd__or2_1 _48509_ (.A(_19568_),
    .B(_19622_),
    .X(_19623_));
 sky130_fd_sc_hd__nand2_1 _48510_ (.A(_19568_),
    .B(_19622_),
    .Y(_19624_));
 sky130_fd_sc_hd__and2_1 _48511_ (.A(_19623_),
    .B(_19624_),
    .X(_19625_));
 sky130_fd_sc_hd__or3_1 _48512_ (.A(_18462_),
    .B(_18483_),
    .C(_19625_),
    .X(_19626_));
 sky130_fd_sc_hd__o21ai_1 _48513_ (.A1(_18462_),
    .A2(_18483_),
    .B1(_19625_),
    .Y(_19627_));
 sky130_fd_sc_hd__nand2_1 _48514_ (.A(_19626_),
    .B(_19627_),
    .Y(_19628_));
 sky130_fd_sc_hd__or2_1 _48515_ (.A(_19547_),
    .B(_19628_),
    .X(_19629_));
 sky130_fd_sc_hd__or3b_1 _48516_ (.A(net138),
    .B(net118),
    .C_N(_19628_),
    .X(_19630_));
 sky130_fd_sc_hd__and2_1 _48517_ (.A(_19629_),
    .B(_19630_),
    .X(_19631_));
 sky130_fd_sc_hd__xnor2_1 _48518_ (.A(_19546_),
    .B(_19631_),
    .Y(_19632_));
 sky130_fd_sc_hd__buf_1 _48519_ (.A(_18585_),
    .X(_19633_));
 sky130_fd_sc_hd__and3_1 _48520_ (.A(_19633_),
    .B(_05689_),
    .C(_17769_),
    .X(_19634_));
 sky130_fd_sc_hd__a31o_2 _48521_ (.A1(_18586_),
    .A2(_24776_),
    .A3(_18587_),
    .B1(_19634_),
    .X(_19635_));
 sky130_fd_sc_hd__buf_1 _48522_ (.A(\delay_line[40][6] ),
    .X(_19636_));
 sky130_fd_sc_hd__or3b_2 _48523_ (.A(\delay_line[40][6] ),
    .B(_18585_),
    .C_N(\delay_line[40][4] ),
    .X(_19637_));
 sky130_fd_sc_hd__or3b_1 _48524_ (.A(\delay_line[40][4] ),
    .B(_18585_),
    .C_N(_19636_),
    .X(_19638_));
 sky130_fd_sc_hd__o211a_1 _48525_ (.A1(\delay_line[40][5] ),
    .A2(_19636_),
    .B1(_19637_),
    .C1(_19638_),
    .X(_19639_));
 sky130_fd_sc_hd__nand2_1 _48526_ (.A(_04173_),
    .B(_19639_),
    .Y(_19640_));
 sky130_fd_sc_hd__or2_1 _48527_ (.A(\delay_line[40][2] ),
    .B(_19639_),
    .X(_19641_));
 sky130_fd_sc_hd__and2_2 _48528_ (.A(_19640_),
    .B(_19641_),
    .X(_19642_));
 sky130_fd_sc_hd__xnor2_4 _48529_ (.A(_19635_),
    .B(_19642_),
    .Y(_19643_));
 sky130_fd_sc_hd__a21boi_4 _48530_ (.A1(_18591_),
    .A2(_18593_),
    .B1_N(_18592_),
    .Y(_19644_));
 sky130_fd_sc_hd__xnor2_4 _48531_ (.A(_19643_),
    .B(_19644_),
    .Y(_19645_));
 sky130_fd_sc_hd__and3_1 _48532_ (.A(_00458_),
    .B(net288),
    .C(_18598_),
    .X(_19646_));
 sky130_fd_sc_hd__xor2_2 _48533_ (.A(net289),
    .B(\delay_line[38][6] ),
    .X(_19647_));
 sky130_fd_sc_hd__o21ai_1 _48534_ (.A1(_18596_),
    .A2(_19646_),
    .B1(_19647_),
    .Y(_19648_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48535_ (.A(net288),
    .X(_19649_));
 sky130_fd_sc_hd__a311o_1 _48536_ (.A1(_00458_),
    .A2(_19649_),
    .A3(_18599_),
    .B1(_19647_),
    .C1(_18596_),
    .X(_19650_));
 sky130_fd_sc_hd__and4bb_1 _48537_ (.A_N(_17778_),
    .B_N(_17779_),
    .C(_18599_),
    .D(_05590_),
    .X(_19651_));
 sky130_fd_sc_hd__and3_1 _48538_ (.A(_19648_),
    .B(_19650_),
    .C(_19651_),
    .X(_19652_));
 sky130_fd_sc_hd__a21oi_1 _48539_ (.A1(_19648_),
    .A2(_19650_),
    .B1(_19651_),
    .Y(_19653_));
 sky130_fd_sc_hd__or2_1 _48540_ (.A(_19652_),
    .B(_19653_),
    .X(_19654_));
 sky130_fd_sc_hd__and3b_1 _48541_ (.A_N(_18605_),
    .B(_18607_),
    .C(_05612_),
    .X(_19655_));
 sky130_fd_sc_hd__inv_2 _48542_ (.A(_17788_),
    .Y(_19656_));
 sky130_fd_sc_hd__nor2_1 _48543_ (.A(_18606_),
    .B(net283),
    .Y(_19657_));
 sky130_fd_sc_hd__nand2_1 _48544_ (.A(_18606_),
    .B(net283),
    .Y(_19658_));
 sky130_fd_sc_hd__or3b_2 _48545_ (.A(_19656_),
    .B(_19657_),
    .C_N(_19658_),
    .X(_19659_));
 sky130_fd_sc_hd__inv_2 _48546_ (.A(\delay_line[39][5] ),
    .Y(_19660_));
 sky130_fd_sc_hd__inv_2 _48547_ (.A(net283),
    .Y(_19661_));
 sky130_fd_sc_hd__clkbuf_2 _48548_ (.A(_19661_),
    .X(_19662_));
 sky130_fd_sc_hd__nand2_1 _48549_ (.A(_19660_),
    .B(_19662_),
    .Y(_19663_));
 sky130_fd_sc_hd__a21o_1 _48550_ (.A1(_19663_),
    .A2(_19658_),
    .B1(_18603_),
    .X(_19664_));
 sky130_fd_sc_hd__o211a_1 _48551_ (.A1(_18609_),
    .A2(_19655_),
    .B1(_19659_),
    .C1(_19664_),
    .X(_19665_));
 sky130_fd_sc_hd__a221oi_1 _48552_ (.A1(_18603_),
    .A2(_18606_),
    .B1(_19659_),
    .B2(_19664_),
    .C1(_19655_),
    .Y(_19666_));
 sky130_fd_sc_hd__or3b_2 _48553_ (.A(_19665_),
    .B(_19666_),
    .C_N(_05623_),
    .X(_19667_));
 sky130_fd_sc_hd__o21bai_1 _48554_ (.A1(_19665_),
    .A2(_19666_),
    .B1_N(_05634_),
    .Y(_19668_));
 sky130_fd_sc_hd__inv_2 _48555_ (.A(_18613_),
    .Y(_19669_));
 sky130_fd_sc_hd__a211oi_1 _48556_ (.A1(_19667_),
    .A2(_19668_),
    .B1(_18611_),
    .C1(_19669_),
    .Y(_19670_));
 sky130_fd_sc_hd__o211a_1 _48557_ (.A1(_18611_),
    .A2(_19669_),
    .B1(_19667_),
    .C1(_19668_),
    .X(_19671_));
 sky130_fd_sc_hd__a211oi_2 _48558_ (.A1(_18617_),
    .A2(_18619_),
    .B1(_19670_),
    .C1(_19671_),
    .Y(_19672_));
 sky130_fd_sc_hd__o211a_1 _48559_ (.A1(_19670_),
    .A2(_19671_),
    .B1(_18617_),
    .C1(_18619_),
    .X(_19673_));
 sky130_fd_sc_hd__nor2_1 _48560_ (.A(_19672_),
    .B(_19673_),
    .Y(_19674_));
 sky130_fd_sc_hd__xor2_2 _48561_ (.A(_19654_),
    .B(_19674_),
    .X(_19675_));
 sky130_fd_sc_hd__xor2_4 _48562_ (.A(_19645_),
    .B(_19675_),
    .X(_19676_));
 sky130_fd_sc_hd__and3b_1 _48563_ (.A_N(_04294_),
    .B(_18576_),
    .C(_18572_),
    .X(_19677_));
 sky130_fd_sc_hd__and2b_1 _48564_ (.A_N(_18576_),
    .B(\delay_line[37][6] ),
    .X(_19678_));
 sky130_fd_sc_hd__buf_1 _48565_ (.A(\delay_line[37][6] ),
    .X(_19679_));
 sky130_fd_sc_hd__and2b_1 _48566_ (.A_N(_19679_),
    .B(_18576_),
    .X(_19680_));
 sky130_fd_sc_hd__nor2_1 _48567_ (.A(_19678_),
    .B(_19680_),
    .Y(_19681_));
 sky130_fd_sc_hd__o21a_1 _48568_ (.A1(_18569_),
    .A2(_19677_),
    .B1(_19681_),
    .X(_19682_));
 sky130_fd_sc_hd__a211oi_1 _48569_ (.A1(_17521_),
    .A2(_18572_),
    .B1(_19681_),
    .C1(_18569_),
    .Y(_19683_));
 sky130_fd_sc_hd__nand3_1 _48570_ (.A(_18570_),
    .B(_18573_),
    .C(_17543_),
    .Y(_19684_));
 sky130_fd_sc_hd__o211a_1 _48571_ (.A1(_19682_),
    .A2(_19683_),
    .B1(_18579_),
    .C1(_19684_),
    .X(_19685_));
 sky130_fd_sc_hd__a211oi_1 _48572_ (.A1(_18579_),
    .A2(_19684_),
    .B1(_19682_),
    .C1(_19683_),
    .Y(_19686_));
 sky130_fd_sc_hd__nor2_1 _48573_ (.A(_19685_),
    .B(_19686_),
    .Y(_19687_));
 sky130_fd_sc_hd__nand2_1 _48574_ (.A(_18557_),
    .B(_18558_),
    .Y(_19688_));
 sky130_fd_sc_hd__nand2_1 _48575_ (.A(_18552_),
    .B(_18554_),
    .Y(_19689_));
 sky130_fd_sc_hd__buf_1 _48576_ (.A(\delay_line[35][6] ),
    .X(_19690_));
 sky130_fd_sc_hd__or2_1 _48577_ (.A(_18554_),
    .B(_19690_),
    .X(_19691_));
 sky130_fd_sc_hd__nand2_1 _48578_ (.A(_18550_),
    .B(_19690_),
    .Y(_19692_));
 sky130_fd_sc_hd__nand4_1 _48579_ (.A(_19689_),
    .B(_18555_),
    .C(_19691_),
    .D(_19692_),
    .Y(_19693_));
 sky130_fd_sc_hd__nor2_1 _48580_ (.A(_18554_),
    .B(_19690_),
    .Y(_19694_));
 sky130_fd_sc_hd__and2_1 _48581_ (.A(_18554_),
    .B(\delay_line[35][6] ),
    .X(_19695_));
 sky130_fd_sc_hd__o2bb2ai_2 _48582_ (.A1_N(_19689_),
    .A2_N(_18555_),
    .B1(_19694_),
    .B2(_19695_),
    .Y(_19696_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48583_ (.A(_18552_),
    .X(_19697_));
 sky130_fd_sc_hd__a21oi_1 _48584_ (.A1(_19693_),
    .A2(_19696_),
    .B1(_19697_),
    .Y(_19698_));
 sky130_fd_sc_hd__and3_1 _48585_ (.A(_19693_),
    .B(_19696_),
    .C(_18552_),
    .X(_19699_));
 sky130_fd_sc_hd__nor3_1 _48586_ (.A(_19688_),
    .B(_19698_),
    .C(_19699_),
    .Y(_19700_));
 sky130_fd_sc_hd__o21a_1 _48587_ (.A1(_19698_),
    .A2(_19699_),
    .B1(_19688_),
    .X(_19701_));
 sky130_fd_sc_hd__o21ai_1 _48588_ (.A1(_19700_),
    .A2(_19701_),
    .B1(net302),
    .Y(_19702_));
 sky130_fd_sc_hd__nor2_1 _48589_ (.A(_17673_),
    .B(_18559_),
    .Y(_19703_));
 sky130_fd_sc_hd__nand3_1 _48590_ (.A(_19693_),
    .B(_19696_),
    .C(_19697_),
    .Y(_19704_));
 sky130_fd_sc_hd__nand4b_1 _48591_ (.A_N(_19698_),
    .B(_18557_),
    .C(_18558_),
    .D(_19704_),
    .Y(_19705_));
 sky130_fd_sc_hd__o21ai_1 _48592_ (.A1(_19698_),
    .A2(_19699_),
    .B1(_19688_),
    .Y(_19706_));
 sky130_fd_sc_hd__nand3b_1 _48593_ (.A_N(net302),
    .B(_19705_),
    .C(_19706_),
    .Y(_19707_));
 sky130_fd_sc_hd__nand3_1 _48594_ (.A(_19702_),
    .B(_19703_),
    .C(_19707_),
    .Y(_19708_));
 sky130_fd_sc_hd__o2bb2ai_1 _48595_ (.A1_N(_19707_),
    .A2_N(_19702_),
    .B1(_17673_),
    .B2(_18562_),
    .Y(_19709_));
 sky130_fd_sc_hd__o2bb2a_1 _48596_ (.A1_N(_19708_),
    .A2_N(_19709_),
    .B1(_18562_),
    .B2(_18560_),
    .X(_19710_));
 sky130_fd_sc_hd__or4bb_1 _48597_ (.A(_18562_),
    .B(_18560_),
    .C_N(_19708_),
    .D_N(_19709_),
    .X(_19711_));
 sky130_fd_sc_hd__or3b_1 _48598_ (.A(_19710_),
    .B(_18565_),
    .C_N(_19711_),
    .X(_19712_));
 sky130_fd_sc_hd__a2bb2o_1 _48599_ (.A1_N(_18562_),
    .A2_N(_18560_),
    .B1(_19708_),
    .B2(_19709_),
    .X(_19713_));
 sky130_fd_sc_hd__a21bo_1 _48600_ (.A1(_19711_),
    .A2(_19713_),
    .B1_N(_18565_),
    .X(_19714_));
 sky130_fd_sc_hd__clkbuf_2 _48601_ (.A(\delay_line[36][3] ),
    .X(_19715_));
 sky130_fd_sc_hd__xnor2_2 _48602_ (.A(net298),
    .B(_19715_),
    .Y(_19716_));
 sky130_fd_sc_hd__or3b_1 _48603_ (.A(_18546_),
    .B(_19716_),
    .C_N(_05931_),
    .X(_19717_));
 sky130_fd_sc_hd__inv_2 _48604_ (.A(_19716_),
    .Y(_19718_));
 sky130_fd_sc_hd__or2_1 _48605_ (.A(_18547_),
    .B(_19718_),
    .X(_19719_));
 sky130_fd_sc_hd__and4_1 _48606_ (.A(_19712_),
    .B(_19714_),
    .C(_19717_),
    .D(_19719_),
    .X(_19720_));
 sky130_fd_sc_hd__a22o_1 _48607_ (.A1(_19712_),
    .A2(_19714_),
    .B1(_19717_),
    .B2(_19719_),
    .X(_19721_));
 sky130_fd_sc_hd__and2b_1 _48608_ (.A_N(_19720_),
    .B(_19721_),
    .X(_19722_));
 sky130_fd_sc_hd__xor2_1 _48609_ (.A(_19687_),
    .B(_19722_),
    .X(_19723_));
 sky130_fd_sc_hd__a311o_1 _48610_ (.A1(_18579_),
    .A2(_18568_),
    .A3(_18578_),
    .B1(_18566_),
    .C1(_19723_),
    .X(_19724_));
 sky130_fd_sc_hd__o21ai_1 _48611_ (.A1(_18566_),
    .A2(_18580_),
    .B1(_19723_),
    .Y(_19725_));
 sky130_fd_sc_hd__and2_2 _48612_ (.A(_19724_),
    .B(_19725_),
    .X(_19726_));
 sky130_fd_sc_hd__xnor2_4 _48613_ (.A(_19676_),
    .B(_19726_),
    .Y(_19727_));
 sky130_fd_sc_hd__nor2_1 _48614_ (.A(_19632_),
    .B(_19727_),
    .Y(_19728_));
 sky130_fd_sc_hd__and2_1 _48615_ (.A(_19632_),
    .B(_19727_),
    .X(_19729_));
 sky130_fd_sc_hd__nand2_1 _48616_ (.A(_18535_),
    .B(net119),
    .Y(_19730_));
 sky130_fd_sc_hd__o211a_1 _48617_ (.A1(_19728_),
    .A2(_19729_),
    .B1(_18534_),
    .C1(_19730_),
    .X(_19731_));
 sky130_fd_sc_hd__a211o_1 _48618_ (.A1(_18534_),
    .A2(_19730_),
    .B1(_19728_),
    .C1(_19729_),
    .X(_19732_));
 sky130_fd_sc_hd__or2b_1 _48619_ (.A(_19731_),
    .B_N(_19732_),
    .X(_19733_));
 sky130_fd_sc_hd__xor2_1 _48620_ (.A(_19545_),
    .B(_19733_),
    .X(_19734_));
 sky130_fd_sc_hd__nand2_1 _48621_ (.A(_19544_),
    .B(_19734_),
    .Y(_19735_));
 sky130_fd_sc_hd__or2_1 _48622_ (.A(_19544_),
    .B(_19734_),
    .X(_19736_));
 sky130_fd_sc_hd__and3_1 _48623_ (.A(_19260_),
    .B(_19735_),
    .C(_19736_),
    .X(_19737_));
 sky130_fd_sc_hd__a21oi_1 _48624_ (.A1(_19735_),
    .A2(_19736_),
    .B1(_19260_),
    .Y(_19738_));
 sky130_fd_sc_hd__or2_1 _48625_ (.A(_19737_),
    .B(_19738_),
    .X(_19739_));
 sky130_fd_sc_hd__o21bai_1 _48626_ (.A1(_19256_),
    .A2(_19259_),
    .B1_N(_19739_),
    .Y(_19740_));
 sky130_fd_sc_hd__a21o_1 _48627_ (.A1(_19251_),
    .A2(_19254_),
    .B1(_19255_),
    .X(_19741_));
 sky130_fd_sc_hd__and3_1 _48628_ (.A(_19248_),
    .B(_19242_),
    .C(_19246_),
    .X(_19742_));
 sky130_fd_sc_hd__o21ai_2 _48629_ (.A1(_19244_),
    .A2(_18705_),
    .B1(_19253_),
    .Y(_19743_));
 sky130_fd_sc_hd__o221ai_2 _48630_ (.A1(_19257_),
    .A2(_19258_),
    .B1(_19742_),
    .B2(_19743_),
    .C1(_19251_),
    .Y(_19744_));
 sky130_fd_sc_hd__o211ai_1 _48631_ (.A1(_19737_),
    .A2(_19738_),
    .B1(_19741_),
    .C1(_19744_),
    .Y(_19745_));
 sky130_fd_sc_hd__nand3b_2 _48632_ (.A_N(_18835_),
    .B(_19740_),
    .C(_19745_),
    .Y(_19746_));
 sky130_fd_sc_hd__o22ai_1 _48633_ (.A1(_19737_),
    .A2(_19738_),
    .B1(_19256_),
    .B2(_19259_),
    .Y(_19747_));
 sky130_fd_sc_hd__nand3b_1 _48634_ (.A_N(_19739_),
    .B(_19741_),
    .C(_19744_),
    .Y(_19748_));
 sky130_fd_sc_hd__nand3_2 _48635_ (.A(_18835_),
    .B(_19747_),
    .C(_19748_),
    .Y(_19749_));
 sky130_fd_sc_hd__nand3_2 _48636_ (.A(_18834_),
    .B(_19746_),
    .C(_19749_),
    .Y(_19750_));
 sky130_fd_sc_hd__a21bo_1 _48637_ (.A1(_19746_),
    .A2(_19749_),
    .B1_N(_18833_),
    .X(_19751_));
 sky130_fd_sc_hd__o21a_1 _48638_ (.A1(_18766_),
    .A2(_18768_),
    .B1(_18770_),
    .X(_19752_));
 sky130_fd_sc_hd__o2bb2ai_2 _48639_ (.A1_N(_19750_),
    .A2_N(_19751_),
    .B1(_19752_),
    .B2(_18718_),
    .Y(_19753_));
 sky130_fd_sc_hd__a21oi_1 _48640_ (.A1(_18762_),
    .A2(_18770_),
    .B1(_18718_),
    .Y(_19754_));
 sky130_fd_sc_hd__nand3_2 _48641_ (.A(_19750_),
    .B(_19751_),
    .C(_19754_),
    .Y(_19755_));
 sky130_fd_sc_hd__a21bo_1 _48642_ (.A1(_05161_),
    .A2(_18765_),
    .B1_N(_18782_),
    .X(_19756_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48643_ (.A(_18722_),
    .X(_19757_));
 sky130_fd_sc_hd__and3_1 _48644_ (.A(_05172_),
    .B(_19757_),
    .C(_11361_),
    .X(_19758_));
 sky130_fd_sc_hd__o21ba_1 _48645_ (.A1(_04953_),
    .A2(_18724_),
    .B1_N(_19758_),
    .X(_19759_));
 sky130_fd_sc_hd__or3_1 _48646_ (.A(_18728_),
    .B(_18735_),
    .C(_19759_),
    .X(_19760_));
 sky130_fd_sc_hd__o21ai_1 _48647_ (.A1(_18728_),
    .A2(net210),
    .B1(_19759_),
    .Y(_19761_));
 sky130_fd_sc_hd__and2_1 _48648_ (.A(_19760_),
    .B(_19761_),
    .X(_19762_));
 sky130_fd_sc_hd__xnor2_2 _48649_ (.A(_19756_),
    .B(_19762_),
    .Y(_19763_));
 sky130_fd_sc_hd__a21oi_2 _48650_ (.A1(_18756_),
    .A2(_18761_),
    .B1(_19763_),
    .Y(_19764_));
 sky130_fd_sc_hd__and3_1 _48651_ (.A(_18756_),
    .B(_18761_),
    .C(_19763_),
    .X(_19765_));
 sky130_fd_sc_hd__nor2_1 _48652_ (.A(_19764_),
    .B(_19765_),
    .Y(_19766_));
 sky130_fd_sc_hd__a32oi_4 _48653_ (.A1(_18773_),
    .A2(_18774_),
    .A3(_18775_),
    .B1(_18772_),
    .B2(_18788_),
    .Y(_19767_));
 sky130_fd_sc_hd__a31oi_2 _48654_ (.A1(_19753_),
    .A2(_19755_),
    .A3(_19766_),
    .B1(_19767_),
    .Y(_19768_));
 sky130_fd_sc_hd__a21o_1 _48655_ (.A1(_19753_),
    .A2(_19755_),
    .B1(_19766_),
    .X(_19769_));
 sky130_fd_sc_hd__or2_1 _48656_ (.A(_19764_),
    .B(_19765_),
    .X(_19770_));
 sky130_fd_sc_hd__a21oi_1 _48657_ (.A1(_19753_),
    .A2(_19755_),
    .B1(_19770_),
    .Y(_19771_));
 sky130_fd_sc_hd__nand3_1 _48658_ (.A(_19753_),
    .B(_19755_),
    .C(_19770_),
    .Y(_19772_));
 sky130_fd_sc_hd__nand2_1 _48659_ (.A(_19772_),
    .B(_19767_),
    .Y(_19773_));
 sky130_fd_sc_hd__o2bb2ai_1 _48660_ (.A1_N(_19768_),
    .A2_N(_19769_),
    .B1(_19771_),
    .B2(_19773_),
    .Y(_19774_));
 sky130_fd_sc_hd__nand2_1 _48661_ (.A(_19774_),
    .B(_18785_),
    .Y(_19775_));
 sky130_fd_sc_hd__o21ai_1 _48662_ (.A1(_11251_),
    .A2(_18791_),
    .B1(_18792_),
    .Y(_19776_));
 sky130_fd_sc_hd__inv_2 _48663_ (.A(_19776_),
    .Y(_19777_));
 sky130_fd_sc_hd__o21ai_1 _48664_ (.A1(_18778_),
    .A2(_11614_),
    .B1(_18784_),
    .Y(_19778_));
 sky130_fd_sc_hd__nand2_1 _48665_ (.A(_19769_),
    .B(_19768_),
    .Y(_19779_));
 sky130_fd_sc_hd__o211ai_1 _48666_ (.A1(_19773_),
    .A2(_19771_),
    .B1(_19778_),
    .C1(_19779_),
    .Y(_19780_));
 sky130_fd_sc_hd__nand3_2 _48667_ (.A(_19775_),
    .B(_19777_),
    .C(_19780_),
    .Y(_19781_));
 sky130_fd_sc_hd__o21ai_1 _48668_ (.A1(_19771_),
    .A2(_19773_),
    .B1(_18785_),
    .Y(_19782_));
 sky130_fd_sc_hd__a21o_1 _48669_ (.A1(_19769_),
    .A2(_19768_),
    .B1(_19782_),
    .X(_19783_));
 sky130_fd_sc_hd__a211o_1 _48670_ (.A1(_11240_),
    .A2(_11119_),
    .B1(_10877_),
    .C1(_18791_),
    .X(_19784_));
 sky130_fd_sc_hd__a22oi_2 _48671_ (.A1(_18792_),
    .A2(_19784_),
    .B1(_19774_),
    .B2(_19778_),
    .Y(_19785_));
 sky130_fd_sc_hd__a22oi_4 _48672_ (.A1(_19783_),
    .A2(_19785_),
    .B1(_18795_),
    .B2(_19781_),
    .Y(_19786_));
 sky130_fd_sc_hd__o21a_1 _48673_ (.A1(_18795_),
    .A2(_19781_),
    .B1(_19786_),
    .X(_00037_));
 sky130_fd_sc_hd__a21bo_1 _48674_ (.A1(_19753_),
    .A2(_19766_),
    .B1_N(_19755_),
    .X(_19787_));
 sky130_fd_sc_hd__a21bo_1 _48675_ (.A1(_18834_),
    .A2(_19746_),
    .B1_N(_19749_),
    .X(_19788_));
 sky130_fd_sc_hd__or4bb_2 _48676_ (.A(_19237_),
    .B(_19238_),
    .C_N(_23502_),
    .D_N(_17897_),
    .X(_19789_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48677_ (.A(net365),
    .X(_19790_));
 sky130_fd_sc_hd__and2_1 _48678_ (.A(net365),
    .B(\delay_line[20][7] ),
    .X(_19791_));
 sky130_fd_sc_hd__buf_1 _48679_ (.A(\delay_line[20][7] ),
    .X(_19792_));
 sky130_fd_sc_hd__nor2_1 _48680_ (.A(net365),
    .B(_19792_),
    .Y(_19793_));
 sky130_fd_sc_hd__o2bb2a_1 _48681_ (.A1_N(_18740_),
    .A2_N(_19790_),
    .B1(_19791_),
    .B2(_19793_),
    .X(_19794_));
 sky130_fd_sc_hd__clkbuf_2 _48682_ (.A(_19792_),
    .X(_19795_));
 sky130_fd_sc_hd__nand2_1 _48683_ (.A(\delay_line[20][5] ),
    .B(net365),
    .Y(_19796_));
 sky130_fd_sc_hd__nor2_1 _48684_ (.A(_19795_),
    .B(_19796_),
    .Y(_19797_));
 sky130_fd_sc_hd__nor2_1 _48685_ (.A(_18737_),
    .B(_18738_),
    .Y(_19798_));
 sky130_fd_sc_hd__xnor2_2 _48686_ (.A(_10888_),
    .B(_19798_),
    .Y(_19799_));
 sky130_fd_sc_hd__clkbuf_2 _48687_ (.A(_19799_),
    .X(_19800_));
 sky130_fd_sc_hd__nor3_1 _48688_ (.A(_19794_),
    .B(_19797_),
    .C(_19800_),
    .Y(_19801_));
 sky130_fd_sc_hd__o21a_1 _48689_ (.A1(_19794_),
    .A2(_19797_),
    .B1(_19800_),
    .X(_19802_));
 sky130_fd_sc_hd__a211oi_2 _48690_ (.A1(_18801_),
    .A2(_18803_),
    .B1(_19801_),
    .C1(_19802_),
    .Y(_19803_));
 sky130_fd_sc_hd__o211a_1 _48691_ (.A1(_19801_),
    .A2(_19802_),
    .B1(_18801_),
    .C1(_18803_),
    .X(_19804_));
 sky130_fd_sc_hd__or2_1 _48692_ (.A(_19803_),
    .B(_19804_),
    .X(_19805_));
 sky130_fd_sc_hd__xor2_1 _48693_ (.A(_19789_),
    .B(_19805_),
    .X(_19806_));
 sky130_fd_sc_hd__o21a_1 _48694_ (.A1(_18749_),
    .A2(_18808_),
    .B1(_18807_),
    .X(_19807_));
 sky130_fd_sc_hd__xnor2_1 _48695_ (.A(_19806_),
    .B(_19807_),
    .Y(_19808_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48696_ (.A(\delay_line[17][7] ),
    .X(_19809_));
 sky130_fd_sc_hd__and2_1 _48697_ (.A(\delay_line[17][6] ),
    .B(_19809_),
    .X(_19810_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48698_ (.A(\delay_line[17][6] ),
    .X(_19811_));
 sky130_fd_sc_hd__nor2_1 _48699_ (.A(_19811_),
    .B(_19809_),
    .Y(_19812_));
 sky130_fd_sc_hd__clkbuf_2 _48700_ (.A(_18814_),
    .X(_19813_));
 sky130_fd_sc_hd__a21oi_2 _48701_ (.A1(_10932_),
    .A2(_11438_),
    .B1(_11405_),
    .Y(_19814_));
 sky130_fd_sc_hd__clkbuf_2 _48702_ (.A(_19814_),
    .X(_19815_));
 sky130_fd_sc_hd__nor2_1 _48703_ (.A(_19815_),
    .B(_10767_),
    .Y(_19816_));
 sky130_fd_sc_hd__a221oi_4 _48704_ (.A1(_18729_),
    .A2(_11438_),
    .B1(_04854_),
    .B2(_04832_),
    .C1(_11405_),
    .Y(_19817_));
 sky130_fd_sc_hd__nor3_1 _48705_ (.A(_19813_),
    .B(_19816_),
    .C(_19817_),
    .Y(_19818_));
 sky130_fd_sc_hd__clkbuf_2 _48706_ (.A(_10998_),
    .X(_19819_));
 sky130_fd_sc_hd__o221a_1 _48707_ (.A1(_10987_),
    .A2(_19813_),
    .B1(_19816_),
    .B2(_19817_),
    .C1(_19819_),
    .X(_19820_));
 sky130_fd_sc_hd__nor4_1 _48708_ (.A(_19810_),
    .B(_19812_),
    .C(net181),
    .D(_19820_),
    .Y(_19821_));
 sky130_fd_sc_hd__o22a_1 _48709_ (.A1(_19810_),
    .A2(_19812_),
    .B1(_19818_),
    .B2(_19820_),
    .X(_19822_));
 sky130_fd_sc_hd__a211o_2 _48710_ (.A1(_18818_),
    .A2(_18819_),
    .B1(net172),
    .C1(_19822_),
    .X(_19823_));
 sky130_fd_sc_hd__o211ai_2 _48711_ (.A1(net172),
    .A2(_19822_),
    .B1(_18818_),
    .C1(_18819_),
    .Y(_19824_));
 sky130_fd_sc_hd__buf_1 _48712_ (.A(_18811_),
    .X(_19825_));
 sky130_fd_sc_hd__or2b_1 _48713_ (.A(_19811_),
    .B_N(_19825_),
    .X(_19826_));
 sky130_fd_sc_hd__buf_1 _48714_ (.A(_19811_),
    .X(_19827_));
 sky130_fd_sc_hd__nor2_1 _48715_ (.A(_19827_),
    .B(_18726_),
    .Y(_19828_));
 sky130_fd_sc_hd__a21oi_1 _48716_ (.A1(_18726_),
    .A2(_19826_),
    .B1(_19828_),
    .Y(_19829_));
 sky130_fd_sc_hd__nand3_2 _48717_ (.A(_19823_),
    .B(_19824_),
    .C(_19829_),
    .Y(_19830_));
 sky130_fd_sc_hd__a21o_1 _48718_ (.A1(_19823_),
    .A2(_19824_),
    .B1(_19829_),
    .X(_19831_));
 sky130_fd_sc_hd__nand2_1 _48719_ (.A(_19830_),
    .B(_19831_),
    .Y(_19832_));
 sky130_fd_sc_hd__xor2_1 _48720_ (.A(_19808_),
    .B(_19832_),
    .X(_19833_));
 sky130_fd_sc_hd__inv_2 _48721_ (.A(_19833_),
    .Y(_19834_));
 sky130_fd_sc_hd__a21oi_1 _48722_ (.A1(_19255_),
    .A2(_19251_),
    .B1(_19834_),
    .Y(_19835_));
 sky130_fd_sc_hd__o21ai_1 _48723_ (.A1(_19742_),
    .A2(_19743_),
    .B1(_19835_),
    .Y(_19836_));
 sky130_fd_sc_hd__o2bb2ai_1 _48724_ (.A1_N(_19255_),
    .A2_N(_19250_),
    .B1(_19743_),
    .B2(_19742_),
    .Y(_19837_));
 sky130_fd_sc_hd__nand2_1 _48725_ (.A(_19837_),
    .B(_19834_),
    .Y(_19838_));
 sky130_fd_sc_hd__clkbuf_2 _48726_ (.A(_19838_),
    .X(_19839_));
 sky130_fd_sc_hd__o32ai_2 _48727_ (.A1(_11548_),
    .A2(_18750_),
    .A3(_18808_),
    .B1(_18810_),
    .B2(_18828_),
    .Y(_19840_));
 sky130_fd_sc_hd__a21oi_1 _48728_ (.A1(_19836_),
    .A2(_19839_),
    .B1(_19840_),
    .Y(_19841_));
 sky130_fd_sc_hd__and3_1 _48729_ (.A(_19840_),
    .B(_19836_),
    .C(_19838_),
    .X(_19842_));
 sky130_fd_sc_hd__inv_2 _48730_ (.A(_19737_),
    .Y(_19843_));
 sky130_fd_sc_hd__nand2_1 _48731_ (.A(_19843_),
    .B(_19748_),
    .Y(_19844_));
 sky130_fd_sc_hd__nor2_1 _48732_ (.A(_15383_),
    .B(_19216_),
    .Y(_19845_));
 sky130_fd_sc_hd__and2_1 _48733_ (.A(_15383_),
    .B(_18836_),
    .X(_19846_));
 sky130_fd_sc_hd__and4bb_1 _48734_ (.A_N(_19845_),
    .B_N(_19846_),
    .C(_00370_),
    .D(_19236_),
    .X(_19847_));
 sky130_fd_sc_hd__buf_1 _48735_ (.A(_19236_),
    .X(_19848_));
 sky130_fd_sc_hd__clkbuf_2 _48736_ (.A(_19848_),
    .X(_19849_));
 sky130_fd_sc_hd__o2bb2a_1 _48737_ (.A1_N(_10635_),
    .A2_N(_19849_),
    .B1(_19845_),
    .B2(_19846_),
    .X(_19850_));
 sky130_fd_sc_hd__o32a_2 _48738_ (.A1(_19654_),
    .A2(_19672_),
    .A3(_19673_),
    .B1(_19675_),
    .B2(_19645_),
    .X(_19851_));
 sky130_fd_sc_hd__inv_2 _48739_ (.A(_19102_),
    .Y(_19852_));
 sky130_fd_sc_hd__nor2_1 _48740_ (.A(_19106_),
    .B(_19020_),
    .Y(_19853_));
 sky130_fd_sc_hd__a21boi_2 _48741_ (.A1(_18842_),
    .A2(_18889_),
    .B1_N(_18888_),
    .Y(_19854_));
 sky130_fd_sc_hd__nand2_1 _48742_ (.A(_19035_),
    .B(_19038_),
    .Y(_19855_));
 sky130_fd_sc_hd__nor2_1 _48743_ (.A(_19024_),
    .B(_19025_),
    .Y(_19856_));
 sky130_fd_sc_hd__buf_1 _48744_ (.A(\delay_line[7][2] ),
    .X(_19857_));
 sky130_fd_sc_hd__and2_1 _48745_ (.A(_19857_),
    .B(\delay_line[7][3] ),
    .X(_19858_));
 sky130_fd_sc_hd__nor2_1 _48746_ (.A(_19857_),
    .B(_08954_),
    .Y(_19859_));
 sky130_fd_sc_hd__o21bai_1 _48747_ (.A1(_19858_),
    .A2(_19859_),
    .B1_N(\delay_line[7][7] ),
    .Y(_19860_));
 sky130_fd_sc_hd__o21ai_1 _48748_ (.A1(_19857_),
    .A2(\delay_line[7][3] ),
    .B1(\delay_line[7][7] ),
    .Y(_19861_));
 sky130_fd_sc_hd__a21o_1 _48749_ (.A1(_19857_),
    .A2(_08954_),
    .B1(_19861_),
    .X(_19862_));
 sky130_fd_sc_hd__and3_1 _48750_ (.A(_19860_),
    .B(_19023_),
    .C(_19862_),
    .X(_19863_));
 sky130_fd_sc_hd__a21o_1 _48751_ (.A1(_19862_),
    .A2(_19860_),
    .B1(_19024_),
    .X(_19864_));
 sky130_fd_sc_hd__nand4b_2 _48752_ (.A_N(_19863_),
    .B(_03447_),
    .C(_03139_),
    .D(_19864_),
    .Y(_19865_));
 sky130_fd_sc_hd__a21oi_1 _48753_ (.A1(_19862_),
    .A2(_19860_),
    .B1(_19024_),
    .Y(_19866_));
 sky130_fd_sc_hd__o21ai_2 _48754_ (.A1(_19863_),
    .A2(_19866_),
    .B1(_19021_),
    .Y(_19867_));
 sky130_fd_sc_hd__a22o_1 _48755_ (.A1(_23040_),
    .A2(_18036_),
    .B1(_19865_),
    .B2(_19867_),
    .X(_19868_));
 sky130_fd_sc_hd__nand4_4 _48756_ (.A(_19865_),
    .B(_19867_),
    .C(_23040_),
    .D(_18036_),
    .Y(_19869_));
 sky130_fd_sc_hd__a32o_1 _48757_ (.A1(_23029_),
    .A2(_00073_),
    .A3(_19856_),
    .B1(_19868_),
    .B2(_19869_),
    .X(_19870_));
 sky130_fd_sc_hd__nor2_1 _48758_ (.A(_03458_),
    .B(_22974_),
    .Y(_19871_));
 sky130_fd_sc_hd__nand4_2 _48759_ (.A(_19868_),
    .B(_19869_),
    .C(_19871_),
    .D(_19856_),
    .Y(_19872_));
 sky130_fd_sc_hd__nand2_1 _48760_ (.A(_19870_),
    .B(_19872_),
    .Y(_19873_));
 sky130_fd_sc_hd__a21oi_2 _48761_ (.A1(_18861_),
    .A2(_18864_),
    .B1(_19873_),
    .Y(_19874_));
 sky130_fd_sc_hd__inv_2 _48762_ (.A(_19874_),
    .Y(_19875_));
 sky130_fd_sc_hd__o211a_1 _48763_ (.A1(_18042_),
    .A2(_18862_),
    .B1(_18864_),
    .C1(_19873_),
    .X(_19876_));
 sky130_fd_sc_hd__a21oi_2 _48764_ (.A1(_19028_),
    .A2(_19030_),
    .B1(_19876_),
    .Y(_19877_));
 sky130_fd_sc_hd__nor2_1 _48765_ (.A(_19874_),
    .B(_19876_),
    .Y(_19878_));
 sky130_fd_sc_hd__nand2_1 _48766_ (.A(_19028_),
    .B(_19030_),
    .Y(_19879_));
 sky130_fd_sc_hd__o2bb2ai_2 _48767_ (.A1_N(_19875_),
    .A2_N(_19877_),
    .B1(_19878_),
    .B2(_19879_),
    .Y(_19880_));
 sky130_fd_sc_hd__xnor2_2 _48768_ (.A(_19855_),
    .B(_19880_),
    .Y(_19881_));
 sky130_fd_sc_hd__buf_2 _48769_ (.A(_19070_),
    .X(_19882_));
 sky130_fd_sc_hd__clkbuf_2 _48770_ (.A(_19882_),
    .X(_19883_));
 sky130_fd_sc_hd__and4_1 _48771_ (.A(_19044_),
    .B(_19883_),
    .C(_19045_),
    .D(_18098_),
    .X(_19884_));
 sky130_fd_sc_hd__buf_1 _48772_ (.A(\delay_line[3][7] ),
    .X(_19885_));
 sky130_fd_sc_hd__or2b_1 _48773_ (.A(\delay_line[3][5] ),
    .B_N(_19885_),
    .X(_19886_));
 sky130_fd_sc_hd__or2b_1 _48774_ (.A(\delay_line[3][7] ),
    .B_N(\delay_line[3][5] ),
    .X(_19887_));
 sky130_fd_sc_hd__and2b_1 _48775_ (.A_N(_13592_),
    .B(_19047_),
    .X(_19888_));
 sky130_fd_sc_hd__a21o_1 _48776_ (.A1(_19886_),
    .A2(_19887_),
    .B1(_19888_),
    .X(_19889_));
 sky130_fd_sc_hd__nand3_1 _48777_ (.A(_19886_),
    .B(_19887_),
    .C(_19888_),
    .Y(_19890_));
 sky130_fd_sc_hd__nand3_2 _48778_ (.A(_19889_),
    .B(_19073_),
    .C(_19890_),
    .Y(_19891_));
 sky130_fd_sc_hd__a21o_1 _48779_ (.A1(_19890_),
    .A2(_19889_),
    .B1(_19073_),
    .X(_19892_));
 sky130_fd_sc_hd__nand3b_2 _48780_ (.A_N(_19052_),
    .B(_19891_),
    .C(_19892_),
    .Y(_19893_));
 sky130_fd_sc_hd__a32o_1 _48781_ (.A1(_18123_),
    .A2(_19048_),
    .A3(_19049_),
    .B1(_19891_),
    .B2(_19892_),
    .X(_19894_));
 sky130_fd_sc_hd__o211a_1 _48782_ (.A1(net237),
    .A2(_19884_),
    .B1(_19893_),
    .C1(_19894_),
    .X(_19895_));
 sky130_fd_sc_hd__a211oi_1 _48783_ (.A1(_19893_),
    .A2(_19894_),
    .B1(net237),
    .C1(_19884_),
    .Y(_19896_));
 sky130_fd_sc_hd__and2_1 _48784_ (.A(_19053_),
    .B(_19055_),
    .X(_19897_));
 sky130_fd_sc_hd__or3_1 _48785_ (.A(_19895_),
    .B(_19896_),
    .C(_19897_),
    .X(_19898_));
 sky130_fd_sc_hd__o21ai_1 _48786_ (.A1(_19895_),
    .A2(_19896_),
    .B1(_19897_),
    .Y(_19899_));
 sky130_fd_sc_hd__nand2_1 _48787_ (.A(_19898_),
    .B(_19899_),
    .Y(_19900_));
 sky130_fd_sc_hd__nor2_1 _48788_ (.A(_13449_),
    .B(\delay_line[6][3] ),
    .Y(_19901_));
 sky130_fd_sc_hd__nor2_1 _48789_ (.A(_13460_),
    .B(_09217_),
    .Y(_19902_));
 sky130_fd_sc_hd__nor2_1 _48790_ (.A(net429),
    .B(\delay_line[6][7] ),
    .Y(_19903_));
 sky130_fd_sc_hd__buf_2 _48791_ (.A(\delay_line[6][7] ),
    .X(_19904_));
 sky130_fd_sc_hd__nand2_2 _48792_ (.A(net429),
    .B(_19904_),
    .Y(_19905_));
 sky130_fd_sc_hd__nand3b_2 _48793_ (.A_N(_19903_),
    .B(_19066_),
    .C(_19905_),
    .Y(_19906_));
 sky130_fd_sc_hd__and2_1 _48794_ (.A(net429),
    .B(\delay_line[6][7] ),
    .X(_19907_));
 sky130_fd_sc_hd__o21bai_1 _48795_ (.A1(_19907_),
    .A2(_19903_),
    .B1_N(_19065_),
    .Y(_19908_));
 sky130_fd_sc_hd__a2bb2o_1 _48796_ (.A1_N(_19901_),
    .A2_N(_19902_),
    .B1(_19906_),
    .B2(_19908_),
    .X(_19909_));
 sky130_fd_sc_hd__nor2_1 _48797_ (.A(_19901_),
    .B(_19902_),
    .Y(_19910_));
 sky130_fd_sc_hd__nand3_1 _48798_ (.A(_19910_),
    .B(_19906_),
    .C(_19908_),
    .Y(_19911_));
 sky130_fd_sc_hd__nand4_2 _48799_ (.A(_19909_),
    .B(_19911_),
    .C(_23018_),
    .D(_03447_),
    .Y(_19912_));
 sky130_fd_sc_hd__a21oi_1 _48800_ (.A1(_19906_),
    .A2(_19908_),
    .B1(_19910_),
    .Y(_19913_));
 sky130_fd_sc_hd__and3_1 _48801_ (.A(_19910_),
    .B(_19906_),
    .C(_19908_),
    .X(_19914_));
 sky130_fd_sc_hd__o22ai_4 _48802_ (.A1(_22974_),
    .A2(_00062_),
    .B1(_19913_),
    .B2(_19914_),
    .Y(_19915_));
 sky130_fd_sc_hd__nor2_1 _48803_ (.A(_19064_),
    .B(_19066_),
    .Y(_19916_));
 sky130_fd_sc_hd__o22a_1 _48804_ (.A1(_03403_),
    .A2(_18094_),
    .B1(_19916_),
    .B2(_09437_),
    .X(_19917_));
 sky130_fd_sc_hd__and3_1 _48805_ (.A(_19912_),
    .B(_19915_),
    .C(_19917_),
    .X(_19918_));
 sky130_fd_sc_hd__a21oi_1 _48806_ (.A1(_19912_),
    .A2(_19915_),
    .B1(_19917_),
    .Y(_19919_));
 sky130_fd_sc_hd__nand2_1 _48807_ (.A(_18103_),
    .B(_18104_),
    .Y(_19920_));
 sky130_fd_sc_hd__nand2_1 _48808_ (.A(_19044_),
    .B(_19070_),
    .Y(_19921_));
 sky130_fd_sc_hd__or2b_1 _48809_ (.A(\delay_line[5][6] ),
    .B_N(\delay_line[5][5] ),
    .X(_19922_));
 sky130_fd_sc_hd__nand3_1 _48810_ (.A(_19920_),
    .B(_19921_),
    .C(_19922_),
    .Y(_19923_));
 sky130_fd_sc_hd__or3b_1 _48811_ (.A(_19070_),
    .B(_19043_),
    .C_N(_13559_),
    .X(_19924_));
 sky130_fd_sc_hd__a21oi_1 _48812_ (.A1(_19923_),
    .A2(_19924_),
    .B1(_03590_),
    .Y(_19925_));
 sky130_fd_sc_hd__and3_1 _48813_ (.A(_19924_),
    .B(_03590_),
    .C(_19923_),
    .X(_19926_));
 sky130_fd_sc_hd__inv_2 _48814_ (.A(\delay_line[5][7] ),
    .Y(_19927_));
 sky130_fd_sc_hd__nor2_2 _48815_ (.A(\delay_line[6][0] ),
    .B(_19927_),
    .Y(_19928_));
 sky130_fd_sc_hd__nand2_1 _48816_ (.A(_19927_),
    .B(_22897_),
    .Y(_19929_));
 sky130_fd_sc_hd__and4b_1 _48817_ (.A_N(_19928_),
    .B(_19929_),
    .C(_19062_),
    .D(\delay_line[6][3] ),
    .X(_19930_));
 sky130_fd_sc_hd__nor2_1 _48818_ (.A(\delay_line[5][7] ),
    .B(_18096_),
    .Y(_19931_));
 sky130_fd_sc_hd__a2bb2o_1 _48819_ (.A1_N(_19928_),
    .A2_N(_19931_),
    .B1(_19062_),
    .B2(_18094_),
    .X(_19932_));
 sky130_fd_sc_hd__nand4b_1 _48820_ (.A_N(_19930_),
    .B(_19932_),
    .C(_19882_),
    .D(_18107_),
    .Y(_19933_));
 sky130_fd_sc_hd__o2bb2a_1 _48821_ (.A1_N(_03403_),
    .A2_N(_18094_),
    .B1(_19928_),
    .B2(_19931_),
    .X(_19934_));
 sky130_fd_sc_hd__o2bb2ai_1 _48822_ (.A1_N(_19882_),
    .A2_N(_18107_),
    .B1(_19930_),
    .B2(_19934_),
    .Y(_19935_));
 sky130_fd_sc_hd__o211a_1 _48823_ (.A1(_19925_),
    .A2(_19926_),
    .B1(_19933_),
    .C1(_19935_),
    .X(_19936_));
 sky130_fd_sc_hd__a211oi_1 _48824_ (.A1(_19933_),
    .A2(_19935_),
    .B1(_19925_),
    .C1(_19926_),
    .Y(_19937_));
 sky130_fd_sc_hd__nor2_1 _48825_ (.A(_19918_),
    .B(_19919_),
    .Y(_19938_));
 sky130_fd_sc_hd__nor2_1 _48826_ (.A(_19936_),
    .B(_19937_),
    .Y(_19939_));
 sky130_fd_sc_hd__or2_1 _48827_ (.A(_19938_),
    .B(_19939_),
    .X(_19940_));
 sky130_fd_sc_hd__o41ai_1 _48828_ (.A1(_19918_),
    .A2(_19919_),
    .A3(_19936_),
    .A4(_19937_),
    .B1(_19940_),
    .Y(_19941_));
 sky130_fd_sc_hd__a21o_1 _48829_ (.A1(_19079_),
    .A2(_19080_),
    .B1(net147),
    .X(_19942_));
 sky130_fd_sc_hd__nand3_1 _48830_ (.A(_19079_),
    .B(_19080_),
    .C(net147),
    .Y(_19943_));
 sky130_fd_sc_hd__nand2_1 _48831_ (.A(_19942_),
    .B(_19943_),
    .Y(_19944_));
 sky130_fd_sc_hd__xor2_2 _48832_ (.A(_19900_),
    .B(_19944_),
    .X(_19945_));
 sky130_fd_sc_hd__nand2_1 _48833_ (.A(_19881_),
    .B(_19945_),
    .Y(_19946_));
 sky130_fd_sc_hd__a21oi_2 _48834_ (.A1(_19035_),
    .A2(_19038_),
    .B1(_19880_),
    .Y(_19947_));
 sky130_fd_sc_hd__and3_1 _48835_ (.A(_19035_),
    .B(_19038_),
    .C(_19880_),
    .X(_19948_));
 sky130_fd_sc_hd__o21bai_2 _48836_ (.A1(_19947_),
    .A2(_19948_),
    .B1_N(_19945_),
    .Y(_19949_));
 sky130_fd_sc_hd__and3b_2 _48837_ (.A_N(_19854_),
    .B(_19946_),
    .C(_19949_),
    .X(_19950_));
 sky130_fd_sc_hd__a21bo_1 _48838_ (.A1(_19039_),
    .A2(_19088_),
    .B1_N(_19040_),
    .X(_19951_));
 sky130_fd_sc_hd__a21bo_1 _48839_ (.A1(_19946_),
    .A2(_19949_),
    .B1_N(_19854_),
    .X(_19952_));
 sky130_fd_sc_hd__nand2_1 _48840_ (.A(_19951_),
    .B(_19952_),
    .Y(_19953_));
 sky130_fd_sc_hd__a21boi_2 _48841_ (.A1(_19946_),
    .A2(_19949_),
    .B1_N(_19854_),
    .Y(_19954_));
 sky130_fd_sc_hd__o21bai_2 _48842_ (.A1(_19950_),
    .A2(_19954_),
    .B1_N(_19951_),
    .Y(_19955_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48843_ (.A(\delay_line[10][7] ),
    .X(_19956_));
 sky130_fd_sc_hd__nor2_1 _48844_ (.A(net414),
    .B(net413),
    .Y(_19957_));
 sky130_fd_sc_hd__and2_1 _48845_ (.A(net414),
    .B(\delay_line[10][4] ),
    .X(_19958_));
 sky130_fd_sc_hd__nor2_1 _48846_ (.A(_19957_),
    .B(_19958_),
    .Y(_19959_));
 sky130_fd_sc_hd__or2_1 _48847_ (.A(_19956_),
    .B(_19959_),
    .X(_19960_));
 sky130_fd_sc_hd__buf_1 _48848_ (.A(_19958_),
    .X(_19961_));
 sky130_fd_sc_hd__or3b_1 _48849_ (.A(_19957_),
    .B(_19961_),
    .C_N(_19956_),
    .X(_19962_));
 sky130_fd_sc_hd__a21o_1 _48850_ (.A1(_19960_),
    .A2(_19962_),
    .B1(_18904_),
    .X(_19963_));
 sky130_fd_sc_hd__clkbuf_2 _48851_ (.A(\delay_line[10][6] ),
    .X(_19964_));
 sky130_fd_sc_hd__o2111ai_2 _48852_ (.A1(_18901_),
    .A2(_18902_),
    .B1(_19962_),
    .C1(_19964_),
    .D1(_19960_),
    .Y(_19965_));
 sky130_fd_sc_hd__nand3_1 _48853_ (.A(_19963_),
    .B(_18901_),
    .C(_19965_),
    .Y(_19966_));
 sky130_fd_sc_hd__a21o_1 _48854_ (.A1(_19965_),
    .A2(_19963_),
    .B1(_18901_),
    .X(_19967_));
 sky130_fd_sc_hd__nand2_2 _48855_ (.A(_19966_),
    .B(_19967_),
    .Y(_19968_));
 sky130_fd_sc_hd__and4bb_1 _48856_ (.A_N(_18986_),
    .B_N(_02799_),
    .C(_12130_),
    .D(_18988_),
    .X(_19969_));
 sky130_fd_sc_hd__o21a_1 _48857_ (.A1(_18986_),
    .A2(_17995_),
    .B1(_02799_),
    .X(_19970_));
 sky130_fd_sc_hd__nor3_1 _48858_ (.A(_19969_),
    .B(_19970_),
    .C(_18896_),
    .Y(_19971_));
 sky130_fd_sc_hd__a2bb2o_1 _48859_ (.A1_N(_17992_),
    .A2_N(_18988_),
    .B1(_23238_),
    .B2(_17999_),
    .X(_19972_));
 sky130_fd_sc_hd__o2bb2a_1 _48860_ (.A1_N(_25314_),
    .A2_N(_19972_),
    .B1(_19969_),
    .B2(_19970_),
    .X(_19973_));
 sky130_fd_sc_hd__nor2_1 _48861_ (.A(_19971_),
    .B(_19973_),
    .Y(_19974_));
 sky130_fd_sc_hd__xor2_2 _48862_ (.A(_19968_),
    .B(_19974_),
    .X(_19975_));
 sky130_fd_sc_hd__nand4_1 _48863_ (.A(_18895_),
    .B(_18896_),
    .C(_17921_),
    .D(_12163_),
    .Y(_19976_));
 sky130_fd_sc_hd__o21ai_1 _48864_ (.A1(_18906_),
    .A2(_18898_),
    .B1(_19976_),
    .Y(_19977_));
 sky130_fd_sc_hd__nor2_1 _48865_ (.A(_19975_),
    .B(_19977_),
    .Y(_19978_));
 sky130_fd_sc_hd__and2_1 _48866_ (.A(_19975_),
    .B(_19977_),
    .X(_19979_));
 sky130_fd_sc_hd__a32o_1 _48867_ (.A1(_18971_),
    .A2(_18972_),
    .A3(_18973_),
    .B1(_18970_),
    .B2(_18977_),
    .X(_19980_));
 sky130_fd_sc_hd__a2bb2o_2 _48868_ (.A1_N(_18951_),
    .A2_N(_18955_),
    .B1(_18965_),
    .B2(_18960_),
    .X(_19981_));
 sky130_fd_sc_hd__buf_2 _48869_ (.A(_17950_),
    .X(_19982_));
 sky130_fd_sc_hd__buf_2 _48870_ (.A(_18948_),
    .X(_19983_));
 sky130_fd_sc_hd__and3_2 _48871_ (.A(_12570_),
    .B(_19982_),
    .C(_19983_),
    .X(_19984_));
 sky130_fd_sc_hd__a21oi_2 _48872_ (.A1(_19982_),
    .A2(_19983_),
    .B1(_12570_),
    .Y(_19985_));
 sky130_fd_sc_hd__buf_2 _48873_ (.A(\delay_line[0][7] ),
    .X(_19986_));
 sky130_fd_sc_hd__nor2_1 _48874_ (.A(_18948_),
    .B(_19986_),
    .Y(_19987_));
 sky130_fd_sc_hd__and2_2 _48875_ (.A(_18948_),
    .B(\delay_line[0][7] ),
    .X(_19988_));
 sky130_fd_sc_hd__nand4_1 _48876_ (.A(_08140_),
    .B(_17941_),
    .C(_18930_),
    .D(_18931_),
    .Y(_19989_));
 sky130_fd_sc_hd__inv_2 _48877_ (.A(\delay_line[4][3] ),
    .Y(_19990_));
 sky130_fd_sc_hd__a21oi_1 _48878_ (.A1(_19990_),
    .A2(_12240_),
    .B1(_17940_),
    .Y(_19991_));
 sky130_fd_sc_hd__or2b_2 _48879_ (.A(net434),
    .B_N(\delay_line[4][2] ),
    .X(_19992_));
 sky130_fd_sc_hd__clkbuf_2 _48880_ (.A(net434),
    .X(_19993_));
 sky130_fd_sc_hd__buf_2 _48881_ (.A(_19993_),
    .X(_19994_));
 sky130_fd_sc_hd__nand2_1 _48882_ (.A(_17941_),
    .B(_19994_),
    .Y(_19995_));
 sky130_fd_sc_hd__clkbuf_2 _48883_ (.A(_19995_),
    .X(_19996_));
 sky130_fd_sc_hd__nand2_1 _48884_ (.A(_19992_),
    .B(_19996_),
    .Y(_19997_));
 sky130_fd_sc_hd__o21ai_1 _48885_ (.A1(_18925_),
    .A2(_19991_),
    .B1(_19997_),
    .Y(_19998_));
 sky130_fd_sc_hd__o21ai_1 _48886_ (.A1(_18923_),
    .A2(_12339_),
    .B1(_17946_),
    .Y(_19999_));
 sky130_fd_sc_hd__o2111ai_1 _48887_ (.A1(_12251_),
    .A2(_19990_),
    .B1(_19992_),
    .C1(_19996_),
    .D1(_19999_),
    .Y(_20000_));
 sky130_fd_sc_hd__and3_1 _48888_ (.A(_19989_),
    .B(_19998_),
    .C(_20000_),
    .X(_20001_));
 sky130_fd_sc_hd__clkbuf_2 _48889_ (.A(\delay_line[11][4] ),
    .X(_20002_));
 sky130_fd_sc_hd__clkbuf_2 _48890_ (.A(\delay_line[11][5] ),
    .X(_20003_));
 sky130_fd_sc_hd__nor2_1 _48891_ (.A(_20002_),
    .B(_20003_),
    .Y(_20004_));
 sky130_fd_sc_hd__clkbuf_2 _48892_ (.A(\delay_line[11][5] ),
    .X(_20005_));
 sky130_fd_sc_hd__and2_1 _48893_ (.A(_18933_),
    .B(_20005_),
    .X(_20006_));
 sky130_fd_sc_hd__o21ai_2 _48894_ (.A1(_20004_),
    .A2(_20006_),
    .B1(_07986_),
    .Y(_20007_));
 sky130_fd_sc_hd__o21ba_1 _48895_ (.A1(_20002_),
    .A2(_20005_),
    .B1_N(_07986_),
    .X(_20008_));
 sky130_fd_sc_hd__nand2_1 _48896_ (.A(_20002_),
    .B(_20005_),
    .Y(_20009_));
 sky130_fd_sc_hd__nand2_1 _48897_ (.A(_20008_),
    .B(_20009_),
    .Y(_20010_));
 sky130_fd_sc_hd__nand3_2 _48898_ (.A(_20007_),
    .B(_18935_),
    .C(_20010_),
    .Y(_20011_));
 sky130_fd_sc_hd__clkbuf_2 _48899_ (.A(_20011_),
    .X(_20012_));
 sky130_fd_sc_hd__a2bb2o_1 _48900_ (.A1_N(_02513_),
    .A2_N(_18934_),
    .B1(_20010_),
    .B2(_20007_),
    .X(_20013_));
 sky130_fd_sc_hd__nand4b_2 _48901_ (.A_N(_19993_),
    .B(_18929_),
    .C(_18931_),
    .D(_17935_),
    .Y(_20014_));
 sky130_fd_sc_hd__clkbuf_2 _48902_ (.A(_20014_),
    .X(_20015_));
 sky130_fd_sc_hd__clkbuf_2 _48903_ (.A(_20015_),
    .X(_20016_));
 sky130_fd_sc_hd__nand3_1 _48904_ (.A(_20012_),
    .B(_20013_),
    .C(_20016_),
    .Y(_20017_));
 sky130_fd_sc_hd__clkbuf_2 _48905_ (.A(_20011_),
    .X(_20018_));
 sky130_fd_sc_hd__inv_2 _48906_ (.A(_20018_),
    .Y(_20019_));
 sky130_fd_sc_hd__a21oi_1 _48907_ (.A1(_20010_),
    .A2(_20007_),
    .B1(_18936_),
    .Y(_20020_));
 sky130_fd_sc_hd__nand3_1 _48908_ (.A(_19989_),
    .B(_19998_),
    .C(_20000_),
    .Y(_20021_));
 sky130_fd_sc_hd__nand2_1 _48909_ (.A(_20016_),
    .B(_20021_),
    .Y(_20022_));
 sky130_fd_sc_hd__o21ai_1 _48910_ (.A1(_20019_),
    .A2(_20020_),
    .B1(_20022_),
    .Y(_20023_));
 sky130_fd_sc_hd__o211a_1 _48911_ (.A1(_20001_),
    .A2(_20017_),
    .B1(_18941_),
    .C1(_20023_),
    .X(_20024_));
 sky130_fd_sc_hd__clkbuf_2 _48912_ (.A(_20023_),
    .X(_20025_));
 sky130_fd_sc_hd__nand4_2 _48913_ (.A(_20012_),
    .B(_20013_),
    .C(_20016_),
    .D(_20021_),
    .Y(_20026_));
 sky130_fd_sc_hd__a21oi_4 _48914_ (.A1(_20025_),
    .A2(_20026_),
    .B1(_18941_),
    .Y(_20027_));
 sky130_fd_sc_hd__o22ai_4 _48915_ (.A1(_19987_),
    .A2(_19988_),
    .B1(_20024_),
    .B2(_20027_),
    .Y(_20028_));
 sky130_fd_sc_hd__a21o_1 _48916_ (.A1(_20025_),
    .A2(_20026_),
    .B1(_18941_),
    .X(_20029_));
 sky130_fd_sc_hd__nor2_1 _48917_ (.A(_19987_),
    .B(_19988_),
    .Y(_20030_));
 sky130_fd_sc_hd__o211ai_2 _48918_ (.A1(_20001_),
    .A2(_20017_),
    .B1(_18941_),
    .C1(_20025_),
    .Y(_20031_));
 sky130_fd_sc_hd__nand3_1 _48919_ (.A(_20029_),
    .B(_20030_),
    .C(_20031_),
    .Y(_20032_));
 sky130_fd_sc_hd__a21bo_2 _48920_ (.A1(_18950_),
    .A2(_18946_),
    .B1_N(_18942_),
    .X(_20033_));
 sky130_fd_sc_hd__a21oi_2 _48921_ (.A1(_20028_),
    .A2(_20032_),
    .B1(_20033_),
    .Y(_20034_));
 sky130_fd_sc_hd__nand2_1 _48922_ (.A(_20031_),
    .B(_20030_),
    .Y(_20035_));
 sky130_fd_sc_hd__o211a_1 _48923_ (.A1(_20035_),
    .A2(_20027_),
    .B1(_20033_),
    .C1(_20028_),
    .X(_20036_));
 sky130_fd_sc_hd__o22ai_4 _48924_ (.A1(_19984_),
    .A2(_19985_),
    .B1(_20034_),
    .B2(_20036_),
    .Y(_20037_));
 sky130_fd_sc_hd__a21o_1 _48925_ (.A1(_20028_),
    .A2(_20032_),
    .B1(_20033_),
    .X(_20038_));
 sky130_fd_sc_hd__o211ai_4 _48926_ (.A1(_20035_),
    .A2(_20027_),
    .B1(_20033_),
    .C1(_20028_),
    .Y(_20039_));
 sky130_fd_sc_hd__nor2_1 _48927_ (.A(_19984_),
    .B(_19985_),
    .Y(_20040_));
 sky130_fd_sc_hd__nand3_2 _48928_ (.A(_20038_),
    .B(_20039_),
    .C(_20040_),
    .Y(_20041_));
 sky130_fd_sc_hd__nand3_2 _48929_ (.A(_19981_),
    .B(_20037_),
    .C(_20041_),
    .Y(_20042_));
 sky130_fd_sc_hd__o21ai_1 _48930_ (.A1(_20034_),
    .A2(_20036_),
    .B1(_20040_),
    .Y(_20043_));
 sky130_fd_sc_hd__o211ai_2 _48931_ (.A1(_19984_),
    .A2(_19985_),
    .B1(_20038_),
    .C1(_20039_),
    .Y(_20044_));
 sky130_fd_sc_hd__nand3b_4 _48932_ (.A_N(_19981_),
    .B(_20043_),
    .C(_20044_),
    .Y(_20045_));
 sky130_fd_sc_hd__clkbuf_4 _48933_ (.A(\delay_line[13][7] ),
    .X(_20046_));
 sky130_fd_sc_hd__nor2_1 _48934_ (.A(net397),
    .B(_20046_),
    .Y(_20047_));
 sky130_fd_sc_hd__and2_1 _48935_ (.A(net397),
    .B(\delay_line[13][7] ),
    .X(_20048_));
 sky130_fd_sc_hd__or3_1 _48936_ (.A(_18914_),
    .B(_20047_),
    .C(_20048_),
    .X(_20049_));
 sky130_fd_sc_hd__a2bb2o_1 _48937_ (.A1_N(_20047_),
    .A2_N(_20048_),
    .B1(_12207_),
    .B2(_18913_),
    .X(_20050_));
 sky130_fd_sc_hd__and3_1 _48938_ (.A(_20049_),
    .B(_20050_),
    .C(_18964_),
    .X(_20051_));
 sky130_fd_sc_hd__clkbuf_2 _48939_ (.A(_20051_),
    .X(_20052_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48940_ (.A(_20049_),
    .X(_20053_));
 sky130_fd_sc_hd__a21oi_1 _48941_ (.A1(_20053_),
    .A2(_20050_),
    .B1(_18967_),
    .Y(_20054_));
 sky130_fd_sc_hd__o2bb2ai_2 _48942_ (.A1_N(_20042_),
    .A2_N(_20045_),
    .B1(_20052_),
    .B2(_20054_),
    .Y(_20055_));
 sky130_fd_sc_hd__and3b_1 _48943_ (.A_N(_18967_),
    .B(_20053_),
    .C(_20050_),
    .X(_20056_));
 sky130_fd_sc_hd__a21boi_2 _48944_ (.A1(_20053_),
    .A2(_20050_),
    .B1_N(_18967_),
    .Y(_20057_));
 sky130_fd_sc_hd__o211ai_4 _48945_ (.A1(_20056_),
    .A2(_20057_),
    .B1(_20042_),
    .C1(_20045_),
    .Y(_20058_));
 sky130_fd_sc_hd__clkbuf_2 _48946_ (.A(_02689_),
    .X(_20059_));
 sky130_fd_sc_hd__clkbuf_2 _48947_ (.A(net405),
    .X(_20060_));
 sky130_fd_sc_hd__nand2_2 _48948_ (.A(\delay_line[12][6] ),
    .B(_20060_),
    .Y(_20061_));
 sky130_fd_sc_hd__buf_2 _48949_ (.A(_20060_),
    .X(_20062_));
 sky130_fd_sc_hd__and2b_1 _48950_ (.A_N(\delay_line[12][5] ),
    .B(_18984_),
    .X(_20063_));
 sky130_fd_sc_hd__o22ai_4 _48951_ (.A1(_20061_),
    .A2(_18987_),
    .B1(_20062_),
    .B2(_20063_),
    .Y(_20064_));
 sky130_fd_sc_hd__xor2_2 _48952_ (.A(_08393_),
    .B(_20064_),
    .X(_20065_));
 sky130_fd_sc_hd__xnor2_2 _48953_ (.A(_18920_),
    .B(_20065_),
    .Y(_20066_));
 sky130_fd_sc_hd__nor3_2 _48954_ (.A(_20059_),
    .B(_18991_),
    .C(_20066_),
    .Y(_20067_));
 sky130_fd_sc_hd__o21a_1 _48955_ (.A1(_20059_),
    .A2(_18991_),
    .B1(_20066_),
    .X(_20068_));
 sky130_fd_sc_hd__nor2_1 _48956_ (.A(_20067_),
    .B(_20068_),
    .Y(_20069_));
 sky130_fd_sc_hd__a31oi_1 _48957_ (.A1(_19980_),
    .A2(_20055_),
    .A3(_20058_),
    .B1(_20069_),
    .Y(_20070_));
 sky130_fd_sc_hd__o2bb2ai_1 _48958_ (.A1_N(_20042_),
    .A2_N(_20045_),
    .B1(_20056_),
    .B2(_20057_),
    .Y(_20071_));
 sky130_fd_sc_hd__inv_2 _48959_ (.A(_19980_),
    .Y(_20072_));
 sky130_fd_sc_hd__o211ai_1 _48960_ (.A1(_20052_),
    .A2(_20054_),
    .B1(_20042_),
    .C1(_20045_),
    .Y(_20073_));
 sky130_fd_sc_hd__nand3_1 _48961_ (.A(_20071_),
    .B(_20072_),
    .C(_20073_),
    .Y(_20074_));
 sky130_fd_sc_hd__clkbuf_2 _48962_ (.A(_20074_),
    .X(_20075_));
 sky130_fd_sc_hd__a31o_1 _48963_ (.A1(_18912_),
    .A2(_18976_),
    .A3(_18978_),
    .B1(_19002_),
    .X(_20076_));
 sky130_fd_sc_hd__and3b_1 _48964_ (.A_N(_18991_),
    .B(_20066_),
    .C(_08525_),
    .X(_20077_));
 sky130_fd_sc_hd__o21ba_1 _48965_ (.A1(_20059_),
    .A2(_18991_),
    .B1_N(_20066_),
    .X(_20078_));
 sky130_fd_sc_hd__nand3_2 _48966_ (.A(_19980_),
    .B(_20055_),
    .C(_20058_),
    .Y(_20079_));
 sky130_fd_sc_hd__a2bb2oi_1 _48967_ (.A1_N(_20077_),
    .A2_N(_20078_),
    .B1(_20075_),
    .B2(_20079_),
    .Y(_20080_));
 sky130_fd_sc_hd__a211oi_2 _48968_ (.A1(_20070_),
    .A2(_20075_),
    .B1(_20076_),
    .C1(_20080_),
    .Y(_20081_));
 sky130_fd_sc_hd__and3_1 _48969_ (.A(_18912_),
    .B(_18976_),
    .C(_18978_),
    .X(_20082_));
 sky130_fd_sc_hd__o211ai_2 _48970_ (.A1(_20067_),
    .A2(_20068_),
    .B1(_20075_),
    .C1(_20079_),
    .Y(_20083_));
 sky130_fd_sc_hd__nand2_1 _48971_ (.A(_20075_),
    .B(_20079_),
    .Y(_20084_));
 sky130_fd_sc_hd__nand2_1 _48972_ (.A(_20084_),
    .B(_20069_),
    .Y(_20085_));
 sky130_fd_sc_hd__a2bb2oi_2 _48973_ (.A1_N(_20082_),
    .A2_N(_19002_),
    .B1(_20083_),
    .B2(_20085_),
    .Y(_20086_));
 sky130_fd_sc_hd__o22ai_1 _48974_ (.A1(_19978_),
    .A2(_19979_),
    .B1(_20081_),
    .B2(_20086_),
    .Y(_20087_));
 sky130_fd_sc_hd__nor2_1 _48975_ (.A(_18908_),
    .B(_18909_),
    .Y(_20088_));
 sky130_fd_sc_hd__and3_1 _48976_ (.A(_18911_),
    .B(_18994_),
    .C(_18996_),
    .X(_20089_));
 sky130_fd_sc_hd__o21a_1 _48977_ (.A1(_20088_),
    .A2(_20089_),
    .B1(_19004_),
    .X(_20090_));
 sky130_fd_sc_hd__nor2b_2 _48978_ (.A(_19975_),
    .B_N(_19977_),
    .Y(_20091_));
 sky130_fd_sc_hd__o211a_1 _48979_ (.A1(_18906_),
    .A2(_18898_),
    .B1(_19976_),
    .C1(_19975_),
    .X(_20092_));
 sky130_fd_sc_hd__a21oi_1 _48980_ (.A1(_18983_),
    .A2(_19000_),
    .B1(_20082_),
    .Y(_20093_));
 sky130_fd_sc_hd__nand3_1 _48981_ (.A(_20085_),
    .B(_20093_),
    .C(_20083_),
    .Y(_20094_));
 sky130_fd_sc_hd__o211a_1 _48982_ (.A1(_20067_),
    .A2(_20068_),
    .B1(_20075_),
    .C1(_20079_),
    .X(_20095_));
 sky130_fd_sc_hd__o21ai_1 _48983_ (.A1(_20095_),
    .A2(_20080_),
    .B1(_20076_),
    .Y(_20096_));
 sky130_fd_sc_hd__o211ai_1 _48984_ (.A1(_20091_),
    .A2(_20092_),
    .B1(_20094_),
    .C1(_20096_),
    .Y(_20097_));
 sky130_fd_sc_hd__nand3_2 _48985_ (.A(_20087_),
    .B(_20090_),
    .C(_20097_),
    .Y(_20098_));
 sky130_fd_sc_hd__clkbuf_2 _48986_ (.A(\delay_line[8][6] ),
    .X(_20099_));
 sky130_fd_sc_hd__nor3_2 _48987_ (.A(_18040_),
    .B(_20099_),
    .C(\delay_line[8][7] ),
    .Y(_20100_));
 sky130_fd_sc_hd__nand2_1 _48988_ (.A(_18845_),
    .B(\delay_line[8][7] ),
    .Y(_20101_));
 sky130_fd_sc_hd__o21ai_1 _48989_ (.A1(_18845_),
    .A2(\delay_line[8][7] ),
    .B1(_18039_),
    .Y(_20102_));
 sky130_fd_sc_hd__nand2_2 _48990_ (.A(_20101_),
    .B(_20102_),
    .Y(_20103_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _48991_ (.A(\delay_line[8][7] ),
    .X(_20104_));
 sky130_fd_sc_hd__nand2_1 _48992_ (.A(_20104_),
    .B(_18849_),
    .Y(_20105_));
 sky130_fd_sc_hd__o21ai_1 _48993_ (.A1(_20100_),
    .A2(_20103_),
    .B1(_20105_),
    .Y(_20106_));
 sky130_fd_sc_hd__o21ai_2 _48994_ (.A1(_18849_),
    .A2(_18846_),
    .B1(_20106_),
    .Y(_20107_));
 sky130_fd_sc_hd__o221ai_2 _48995_ (.A1(_11822_),
    .A2(_18850_),
    .B1(_20100_),
    .B2(_20103_),
    .C1(_18847_),
    .Y(_20108_));
 sky130_fd_sc_hd__a21o_1 _48996_ (.A1(_20107_),
    .A2(_20108_),
    .B1(_18030_),
    .X(_20109_));
 sky130_fd_sc_hd__nand3_1 _48997_ (.A(_20107_),
    .B(_20108_),
    .C(_18030_),
    .Y(_20110_));
 sky130_fd_sc_hd__and3_1 _48998_ (.A(_20109_),
    .B(_20110_),
    .C(_02876_),
    .X(_20111_));
 sky130_fd_sc_hd__a21oi_1 _48999_ (.A1(_20109_),
    .A2(_20110_),
    .B1(_08877_),
    .Y(_20112_));
 sky130_fd_sc_hd__o21ai_1 _49000_ (.A1(_20111_),
    .A2(_20112_),
    .B1(_18859_),
    .Y(_20113_));
 sky130_fd_sc_hd__or3_2 _49001_ (.A(_20112_),
    .B(_18859_),
    .C(_20111_),
    .X(_20114_));
 sky130_fd_sc_hd__nand2_1 _49002_ (.A(_18857_),
    .B(_18858_),
    .Y(_20115_));
 sky130_fd_sc_hd__xor2_2 _49003_ (.A(_11943_),
    .B(_20115_),
    .X(_20116_));
 sky130_fd_sc_hd__a21oi_1 _49004_ (.A1(_20113_),
    .A2(_20114_),
    .B1(_20116_),
    .Y(_20117_));
 sky130_fd_sc_hd__nand3_2 _49005_ (.A(_20114_),
    .B(_20116_),
    .C(_20113_),
    .Y(_20118_));
 sky130_fd_sc_hd__inv_2 _49006_ (.A(_20118_),
    .Y(_20119_));
 sky130_fd_sc_hd__o21bai_1 _49007_ (.A1(_18876_),
    .A2(_18875_),
    .B1_N(_18877_),
    .Y(_20120_));
 sky130_fd_sc_hd__or3b_1 _49008_ (.A(_18869_),
    .B(_18870_),
    .C_N(_18053_),
    .X(_20121_));
 sky130_fd_sc_hd__clkbuf_4 _49009_ (.A(net421),
    .X(_20122_));
 sky130_fd_sc_hd__buf_2 _49010_ (.A(_20122_),
    .X(_20123_));
 sky130_fd_sc_hd__a21o_1 _49011_ (.A1(_17913_),
    .A2(_20122_),
    .B1(_12976_),
    .X(_20124_));
 sky130_fd_sc_hd__buf_2 _49012_ (.A(net420),
    .X(_20125_));
 sky130_fd_sc_hd__a21boi_1 _49013_ (.A1(_18867_),
    .A2(net420),
    .B1_N(\delay_line[9][5] ),
    .Y(_20126_));
 sky130_fd_sc_hd__o21ai_2 _49014_ (.A1(_18867_),
    .A2(_20125_),
    .B1(_20126_),
    .Y(_20127_));
 sky130_fd_sc_hd__nor2_2 _49015_ (.A(\delay_line[9][6] ),
    .B(net420),
    .Y(_20128_));
 sky130_fd_sc_hd__and2_1 _49016_ (.A(net421),
    .B(net420),
    .X(_20129_));
 sky130_fd_sc_hd__o21bai_2 _49017_ (.A1(_20128_),
    .A2(_20129_),
    .B1_N(_17912_),
    .Y(_20130_));
 sky130_fd_sc_hd__o2111ai_4 _49018_ (.A1(_17913_),
    .A2(_20123_),
    .B1(_20124_),
    .C1(_20127_),
    .D1(_20130_),
    .Y(_20131_));
 sky130_fd_sc_hd__a21oi_1 _49019_ (.A1(_17913_),
    .A2(_20122_),
    .B1(_12976_),
    .Y(_20132_));
 sky130_fd_sc_hd__a2bb2o_1 _49020_ (.A1_N(_18869_),
    .A2_N(_20132_),
    .B1(_20127_),
    .B2(_20130_),
    .X(_20133_));
 sky130_fd_sc_hd__o211a_1 _49021_ (.A1(_18869_),
    .A2(_18870_),
    .B1(_12976_),
    .C1(net422),
    .X(_20134_));
 sky130_fd_sc_hd__a21o_1 _49022_ (.A1(_20131_),
    .A2(_20133_),
    .B1(_20134_),
    .X(_20135_));
 sky130_fd_sc_hd__o21a_1 _49023_ (.A1(_02832_),
    .A2(_18905_),
    .B1(_23106_),
    .X(_20136_));
 sky130_fd_sc_hd__nand3_1 _49024_ (.A(_20134_),
    .B(_20131_),
    .C(_20133_),
    .Y(_20137_));
 sky130_fd_sc_hd__and3_1 _49025_ (.A(_20135_),
    .B(_20136_),
    .C(_20137_),
    .X(_20138_));
 sky130_fd_sc_hd__a21oi_1 _49026_ (.A1(_20137_),
    .A2(_20135_),
    .B1(_20136_),
    .Y(_20139_));
 sky130_fd_sc_hd__nor2_1 _49027_ (.A(_18055_),
    .B(_20121_),
    .Y(_20140_));
 sky130_fd_sc_hd__o21bai_1 _49028_ (.A1(_20138_),
    .A2(_20139_),
    .B1_N(_20140_),
    .Y(_20141_));
 sky130_fd_sc_hd__o41a_1 _49029_ (.A1(_18055_),
    .A2(_20121_),
    .A3(_20138_),
    .A4(_20139_),
    .B1(_20141_),
    .X(_20142_));
 sky130_fd_sc_hd__xor2_1 _49030_ (.A(_20120_),
    .B(_20142_),
    .X(_20143_));
 sky130_fd_sc_hd__o21ba_1 _49031_ (.A1(_20117_),
    .A2(_20119_),
    .B1_N(_20143_),
    .X(_20144_));
 sky130_fd_sc_hd__and3b_1 _49032_ (.A_N(_20117_),
    .B(_20143_),
    .C(_20118_),
    .X(_20145_));
 sky130_fd_sc_hd__o21bai_1 _49033_ (.A1(_20144_),
    .A2(_20145_),
    .B1_N(_19006_),
    .Y(_20146_));
 sky130_fd_sc_hd__o21bai_1 _49034_ (.A1(_20117_),
    .A2(_20119_),
    .B1_N(_20143_),
    .Y(_20147_));
 sky130_fd_sc_hd__nand3b_1 _49035_ (.A_N(_20145_),
    .B(_19006_),
    .C(_20147_),
    .Y(_20148_));
 sky130_fd_sc_hd__a31o_1 _49036_ (.A1(_18883_),
    .A2(_18864_),
    .A3(_18865_),
    .B1(_18882_),
    .X(_20149_));
 sky130_fd_sc_hd__a21oi_1 _49037_ (.A1(_20146_),
    .A2(_20148_),
    .B1(_20149_),
    .Y(_20150_));
 sky130_fd_sc_hd__nand3_1 _49038_ (.A(_20149_),
    .B(_20146_),
    .C(_20148_),
    .Y(_20151_));
 sky130_fd_sc_hd__or2b_1 _49039_ (.A(_20150_),
    .B_N(_20151_),
    .X(_20152_));
 sky130_fd_sc_hd__inv_2 _49040_ (.A(_20152_),
    .Y(_20153_));
 sky130_fd_sc_hd__nand2_1 _49041_ (.A(_20098_),
    .B(_20153_),
    .Y(_20154_));
 sky130_fd_sc_hd__nor2_1 _49042_ (.A(_19978_),
    .B(_19979_),
    .Y(_20155_));
 sky130_fd_sc_hd__a31o_1 _49043_ (.A1(_20085_),
    .A2(_20093_),
    .A3(_20083_),
    .B1(_20155_),
    .X(_20156_));
 sky130_fd_sc_hd__inv_2 _49044_ (.A(_20090_),
    .Y(_20157_));
 sky130_fd_sc_hd__o22ai_2 _49045_ (.A1(_20091_),
    .A2(_20092_),
    .B1(_20081_),
    .B2(_20086_),
    .Y(_20158_));
 sky130_fd_sc_hd__o211a_1 _49046_ (.A1(_20156_),
    .A2(_20086_),
    .B1(_20157_),
    .C1(_20158_),
    .X(_20159_));
 sky130_fd_sc_hd__nand2_1 _49047_ (.A(_19010_),
    .B(_19100_),
    .Y(_20160_));
 sky130_fd_sc_hd__o211ai_2 _49048_ (.A1(_20156_),
    .A2(_20086_),
    .B1(_20157_),
    .C1(_20158_),
    .Y(_20161_));
 sky130_fd_sc_hd__a21o_1 _49049_ (.A1(_20161_),
    .A2(_20098_),
    .B1(_20153_),
    .X(_20162_));
 sky130_fd_sc_hd__o211ai_4 _49050_ (.A1(_20154_),
    .A2(_20159_),
    .B1(_20160_),
    .C1(_20162_),
    .Y(_20163_));
 sky130_fd_sc_hd__nand2_1 _49051_ (.A(_20161_),
    .B(_20098_),
    .Y(_20164_));
 sky130_fd_sc_hd__o2bb2ai_1 _49052_ (.A1_N(_20152_),
    .A2_N(_20164_),
    .B1(_20154_),
    .B2(_20159_),
    .Y(_20165_));
 sky130_fd_sc_hd__inv_2 _49053_ (.A(_20160_),
    .Y(_20166_));
 sky130_fd_sc_hd__nand2_2 _49054_ (.A(_20165_),
    .B(_20166_),
    .Y(_20167_));
 sky130_fd_sc_hd__o2111ai_4 _49055_ (.A1(_19950_),
    .A2(_19953_),
    .B1(_19955_),
    .C1(_20163_),
    .D1(_20167_),
    .Y(_20168_));
 sky130_fd_sc_hd__or2_1 _49056_ (.A(_19950_),
    .B(_19953_),
    .X(_20169_));
 sky130_fd_sc_hd__inv_2 _49057_ (.A(_20169_),
    .Y(_20170_));
 sky130_fd_sc_hd__inv_2 _49058_ (.A(_19955_),
    .Y(_20171_));
 sky130_fd_sc_hd__o2bb2ai_1 _49059_ (.A1_N(_20167_),
    .A2_N(_20163_),
    .B1(_20170_),
    .B2(_20171_),
    .Y(_20172_));
 sky130_fd_sc_hd__o211ai_2 _49060_ (.A1(_19852_),
    .A2(_19853_),
    .B1(_20168_),
    .C1(_20172_),
    .Y(_20173_));
 sky130_fd_sc_hd__o21a_1 _49061_ (.A1(_19950_),
    .A2(_19954_),
    .B1(_19951_),
    .X(_20174_));
 sky130_fd_sc_hd__a21o_1 _49062_ (.A1(_19951_),
    .A2(_19952_),
    .B1(_19950_),
    .X(_20175_));
 sky130_fd_sc_hd__nor2_1 _49063_ (.A(_19954_),
    .B(_20175_),
    .Y(_20176_));
 sky130_fd_sc_hd__o2bb2ai_1 _49064_ (.A1_N(_20167_),
    .A2_N(_20163_),
    .B1(_20174_),
    .B2(_20176_),
    .Y(_20177_));
 sky130_fd_sc_hd__o21ai_2 _49065_ (.A1(_19106_),
    .A2(_19020_),
    .B1(_19102_),
    .Y(_20178_));
 sky130_fd_sc_hd__inv_2 _49066_ (.A(_20178_),
    .Y(_20179_));
 sky130_fd_sc_hd__o211ai_1 _49067_ (.A1(_20170_),
    .A2(_20171_),
    .B1(_20167_),
    .C1(_20163_),
    .Y(_20180_));
 sky130_fd_sc_hd__nand3_1 _49068_ (.A(_20177_),
    .B(_20179_),
    .C(_20180_),
    .Y(_20181_));
 sky130_fd_sc_hd__buf_1 _49069_ (.A(_20181_),
    .X(_20182_));
 sky130_fd_sc_hd__nand2_1 _49070_ (.A(_20173_),
    .B(_20182_),
    .Y(_20183_));
 sky130_fd_sc_hd__a31o_2 _49071_ (.A1(_19140_),
    .A2(_19142_),
    .A3(_19143_),
    .B1(_19147_),
    .X(_20184_));
 sky130_fd_sc_hd__o21ai_2 _49072_ (.A1(_14317_),
    .A2(_19118_),
    .B1(_14273_),
    .Y(_20185_));
 sky130_fd_sc_hd__clkbuf_2 _49073_ (.A(_19122_),
    .X(_20186_));
 sky130_fd_sc_hd__o211ai_1 _49074_ (.A1(_18172_),
    .A2(_18174_),
    .B1(_09316_),
    .C1(_20186_),
    .Y(_20187_));
 sky130_fd_sc_hd__a211o_1 _49075_ (.A1(_09316_),
    .A2(_19121_),
    .B1(_18172_),
    .C1(_18174_),
    .X(_20188_));
 sky130_fd_sc_hd__a22o_2 _49076_ (.A1(_18170_),
    .A2(_20185_),
    .B1(_20187_),
    .B2(_20188_),
    .X(_20189_));
 sky130_fd_sc_hd__nand4_1 _49077_ (.A(_18170_),
    .B(_20185_),
    .C(_20187_),
    .D(_20188_),
    .Y(_20190_));
 sky130_fd_sc_hd__buf_1 _49078_ (.A(\delay_line[1][7] ),
    .X(_20191_));
 sky130_fd_sc_hd__nor2_1 _49079_ (.A(net444),
    .B(_20191_),
    .Y(_20192_));
 sky130_fd_sc_hd__clkbuf_2 _49080_ (.A(\delay_line[2][7] ),
    .X(_20193_));
 sky130_fd_sc_hd__nand2_1 _49081_ (.A(net444),
    .B(_20191_),
    .Y(_20194_));
 sky130_fd_sc_hd__nand3b_2 _49082_ (.A_N(_20192_),
    .B(_20193_),
    .C(_20194_),
    .Y(_20195_));
 sky130_fd_sc_hd__and2_1 _49083_ (.A(net444),
    .B(_20191_),
    .X(_20196_));
 sky130_fd_sc_hd__o21bai_1 _49084_ (.A1(_20196_),
    .A2(_20192_),
    .B1_N(\delay_line[2][7] ),
    .Y(_20197_));
 sky130_fd_sc_hd__nand3b_1 _49085_ (.A_N(_19124_),
    .B(_20195_),
    .C(_20197_),
    .Y(_20198_));
 sky130_fd_sc_hd__a2bb2o_1 _49086_ (.A1_N(_19125_),
    .A2_N(_19123_),
    .B1(_20195_),
    .B2(_20197_),
    .X(_20199_));
 sky130_fd_sc_hd__a22o_1 _49087_ (.A1(_20189_),
    .A2(_20190_),
    .B1(_20198_),
    .B2(_20199_),
    .X(_20200_));
 sky130_fd_sc_hd__nand4_2 _49088_ (.A(_20189_),
    .B(_20190_),
    .C(_20198_),
    .D(_20199_),
    .Y(_20201_));
 sky130_fd_sc_hd__nand2_1 _49089_ (.A(_19128_),
    .B(_19131_),
    .Y(_20202_));
 sky130_fd_sc_hd__a21o_1 _49090_ (.A1(_20200_),
    .A2(_20201_),
    .B1(_20202_),
    .X(_20203_));
 sky130_fd_sc_hd__nand3_1 _49091_ (.A(_20202_),
    .B(_20200_),
    .C(_20201_),
    .Y(_20204_));
 sky130_fd_sc_hd__a21o_1 _49092_ (.A1(_03909_),
    .A2(_18172_),
    .B1(_18174_),
    .X(_20205_));
 sky130_fd_sc_hd__and2_1 _49093_ (.A(_20205_),
    .B(_14273_),
    .X(_20206_));
 sky130_fd_sc_hd__nand3_1 _49094_ (.A(_20203_),
    .B(_20204_),
    .C(_20206_),
    .Y(_20207_));
 sky130_fd_sc_hd__a21o_1 _49095_ (.A1(_20203_),
    .A2(_20204_),
    .B1(_20206_),
    .X(_20208_));
 sky130_fd_sc_hd__a21oi_1 _49096_ (.A1(_19042_),
    .A2(_19046_),
    .B1(_19057_),
    .Y(_20209_));
 sky130_fd_sc_hd__a211o_1 _49097_ (.A1(_20207_),
    .A2(_20208_),
    .B1(_20209_),
    .C1(_19060_),
    .X(_20210_));
 sky130_fd_sc_hd__o211ai_2 _49098_ (.A1(_20209_),
    .A2(_19060_),
    .B1(_20207_),
    .C1(_20208_),
    .Y(_20211_));
 sky130_fd_sc_hd__a31o_1 _49099_ (.A1(_19115_),
    .A2(_19131_),
    .A3(_19134_),
    .B1(_19138_),
    .X(_20212_));
 sky130_fd_sc_hd__a21o_1 _49100_ (.A1(_20210_),
    .A2(_20211_),
    .B1(_20212_),
    .X(_20213_));
 sky130_fd_sc_hd__nand3_1 _49101_ (.A(_20212_),
    .B(_20210_),
    .C(_20211_),
    .Y(_20214_));
 sky130_fd_sc_hd__a31o_1 _49102_ (.A1(net211),
    .A2(_19080_),
    .A3(_19083_),
    .B1(_19087_),
    .X(_20215_));
 sky130_fd_sc_hd__a21oi_1 _49103_ (.A1(_20213_),
    .A2(_20214_),
    .B1(_20215_),
    .Y(_20216_));
 sky130_fd_sc_hd__and3_1 _49104_ (.A(_20215_),
    .B(_20213_),
    .C(_20214_),
    .X(_20217_));
 sky130_fd_sc_hd__nor2_1 _49105_ (.A(_20216_),
    .B(_20217_),
    .Y(_20218_));
 sky130_fd_sc_hd__xnor2_2 _49106_ (.A(_20184_),
    .B(_20218_),
    .Y(_20219_));
 sky130_fd_sc_hd__a21o_1 _49107_ (.A1(_19151_),
    .A2(_19154_),
    .B1(_20219_),
    .X(_20220_));
 sky130_fd_sc_hd__and2_1 _49108_ (.A(_19151_),
    .B(_19154_),
    .X(_20221_));
 sky130_fd_sc_hd__nand2_1 _49109_ (.A(_20219_),
    .B(_20221_),
    .Y(_20222_));
 sky130_fd_sc_hd__and3_1 _49110_ (.A(_19095_),
    .B(_20220_),
    .C(_20222_),
    .X(_20223_));
 sky130_fd_sc_hd__a21oi_1 _49111_ (.A1(_20220_),
    .A2(_20222_),
    .B1(_19095_),
    .Y(_20224_));
 sky130_fd_sc_hd__o21ba_1 _49112_ (.A1(_20223_),
    .A2(_20224_),
    .B1_N(_19155_),
    .X(_20225_));
 sky130_fd_sc_hd__nor4b_1 _49113_ (.A(_19156_),
    .B(_20223_),
    .C(_20224_),
    .D_N(_19113_),
    .Y(_20226_));
 sky130_fd_sc_hd__nor2_1 _49114_ (.A(_20225_),
    .B(_20226_),
    .Y(_20227_));
 sky130_fd_sc_hd__buf_1 _49115_ (.A(_20227_),
    .X(_20228_));
 sky130_fd_sc_hd__nand2_1 _49116_ (.A(_20183_),
    .B(_20228_),
    .Y(_20229_));
 sky130_fd_sc_hd__nand3b_1 _49117_ (.A_N(_20227_),
    .B(_20173_),
    .C(_20182_),
    .Y(_20230_));
 sky130_fd_sc_hd__o21ai_1 _49118_ (.A1(_19165_),
    .A2(_19166_),
    .B1(_19112_),
    .Y(_20231_));
 sky130_fd_sc_hd__and2_1 _49119_ (.A(_19171_),
    .B(_20231_),
    .X(_20232_));
 sky130_fd_sc_hd__nand3_2 _49120_ (.A(_20229_),
    .B(_20230_),
    .C(_20232_),
    .Y(_20233_));
 sky130_fd_sc_hd__nand2_1 _49121_ (.A(_20182_),
    .B(_20228_),
    .Y(_20234_));
 sky130_fd_sc_hd__and3_1 _49122_ (.A(_20178_),
    .B(_20168_),
    .C(_20172_),
    .X(_20235_));
 sky130_fd_sc_hd__nand2_1 _49123_ (.A(_19171_),
    .B(_20231_),
    .Y(_20236_));
 sky130_fd_sc_hd__a21o_1 _49124_ (.A1(_20173_),
    .A2(_20181_),
    .B1(_20228_),
    .X(_20237_));
 sky130_fd_sc_hd__o211ai_2 _49125_ (.A1(_20234_),
    .A2(_20235_),
    .B1(_20236_),
    .C1(_20237_),
    .Y(_20238_));
 sky130_fd_sc_hd__o31a_1 _49126_ (.A1(_19158_),
    .A2(_19155_),
    .A3(_19157_),
    .B1(_19160_),
    .X(_20239_));
 sky130_fd_sc_hd__inv_2 _49127_ (.A(_20239_),
    .Y(_20240_));
 sky130_fd_sc_hd__a21oi_4 _49128_ (.A1(_20233_),
    .A2(_20238_),
    .B1(_20240_),
    .Y(_20241_));
 sky130_fd_sc_hd__inv_2 _49129_ (.A(_19179_),
    .Y(_20242_));
 sky130_fd_sc_hd__o21a_1 _49130_ (.A1(_18216_),
    .A2(_18840_),
    .B1(_19173_),
    .X(_20243_));
 sky130_fd_sc_hd__clkbuf_2 _49131_ (.A(_20233_),
    .X(_20244_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49132_ (.A(_20238_),
    .X(_20245_));
 sky130_fd_sc_hd__o211ai_2 _49133_ (.A1(_19162_),
    .A2(_19161_),
    .B1(_20244_),
    .C1(_20245_),
    .Y(_20246_));
 sky130_fd_sc_hd__o21ai_4 _49134_ (.A1(_20242_),
    .A2(_20243_),
    .B1(_20246_),
    .Y(_20247_));
 sky130_fd_sc_hd__nor2_1 _49135_ (.A(_20241_),
    .B(_20247_),
    .Y(_20248_));
 sky130_fd_sc_hd__a21o_1 _49136_ (.A1(_20244_),
    .A2(_20245_),
    .B1(_20240_),
    .X(_20249_));
 sky130_fd_sc_hd__a31o_1 _49137_ (.A1(_19176_),
    .A2(_19177_),
    .A3(_19178_),
    .B1(_20243_),
    .X(_20250_));
 sky130_fd_sc_hd__a21oi_1 _49138_ (.A1(_20249_),
    .A2(_20246_),
    .B1(_20250_),
    .Y(_20251_));
 sky130_fd_sc_hd__a211o_1 _49139_ (.A1(_18233_),
    .A2(_18227_),
    .B1(_19185_),
    .C1(_19188_),
    .X(_20252_));
 sky130_fd_sc_hd__o22a_1 _49140_ (.A1(_19187_),
    .A2(_20252_),
    .B1(_19201_),
    .B2(_19194_),
    .X(_20253_));
 sky130_fd_sc_hd__o21ai_4 _49141_ (.A1(_20248_),
    .A2(_20251_),
    .B1(_20253_),
    .Y(_20254_));
 sky130_fd_sc_hd__o211a_1 _49142_ (.A1(_19162_),
    .A2(_19161_),
    .B1(_20244_),
    .C1(_20245_),
    .X(_20255_));
 sky130_fd_sc_hd__o21bai_4 _49143_ (.A1(_20241_),
    .A2(_20255_),
    .B1_N(_20250_),
    .Y(_20256_));
 sky130_fd_sc_hd__o22ai_4 _49144_ (.A1(_19187_),
    .A2(_20252_),
    .B1(_19201_),
    .B2(_19194_),
    .Y(_20257_));
 sky130_fd_sc_hd__o211ai_4 _49145_ (.A1(_20241_),
    .A2(_20247_),
    .B1(_20256_),
    .C1(_20257_),
    .Y(_20258_));
 sky130_fd_sc_hd__and2_1 _49146_ (.A(\delay_line[23][6] ),
    .B(net349),
    .X(_20259_));
 sky130_fd_sc_hd__nor2_1 _49147_ (.A(_19204_),
    .B(\delay_line[23][7] ),
    .Y(_20260_));
 sky130_fd_sc_hd__nor2_1 _49148_ (.A(_20259_),
    .B(_20260_),
    .Y(_20261_));
 sky130_fd_sc_hd__a21o_1 _49149_ (.A1(_20254_),
    .A2(_20258_),
    .B1(_20261_),
    .X(_20262_));
 sky130_fd_sc_hd__nand3_1 _49150_ (.A(_20254_),
    .B(_20258_),
    .C(_20261_),
    .Y(_20263_));
 sky130_fd_sc_hd__nand3b_1 _49151_ (.A_N(_19851_),
    .B(_20262_),
    .C(_20263_),
    .Y(_20264_));
 sky130_fd_sc_hd__a21bo_1 _49152_ (.A1(_20254_),
    .A2(_20258_),
    .B1_N(_20261_),
    .X(_20265_));
 sky130_fd_sc_hd__clkbuf_2 _49153_ (.A(_20259_),
    .X(_20266_));
 sky130_fd_sc_hd__o211ai_2 _49154_ (.A1(_20266_),
    .A2(_20260_),
    .B1(_20254_),
    .C1(_20258_),
    .Y(_20267_));
 sky130_fd_sc_hd__nand3_2 _49155_ (.A(_20265_),
    .B(_20267_),
    .C(_19851_),
    .Y(_20268_));
 sky130_fd_sc_hd__a2bb2o_1 _49156_ (.A1_N(_19192_),
    .A2_N(_19195_),
    .B1(_19216_),
    .B2(_19205_),
    .X(_20269_));
 sky130_fd_sc_hd__a21o_1 _49157_ (.A1(_20264_),
    .A2(_20268_),
    .B1(_20269_),
    .X(_20270_));
 sky130_fd_sc_hd__nand3_2 _49158_ (.A(_20269_),
    .B(_20264_),
    .C(_20268_),
    .Y(_20271_));
 sky130_fd_sc_hd__a21bo_2 _49159_ (.A1(_19676_),
    .A2(_19726_),
    .B1_N(_19725_),
    .X(_20272_));
 sky130_fd_sc_hd__a21oi_4 _49160_ (.A1(_20270_),
    .A2(_20271_),
    .B1(_20272_),
    .Y(_20273_));
 sky130_fd_sc_hd__nand2_1 _49161_ (.A(_20269_),
    .B(_20268_),
    .Y(_20274_));
 sky130_fd_sc_hd__a21oi_1 _49162_ (.A1(_20265_),
    .A2(_20267_),
    .B1(_19851_),
    .Y(_20275_));
 sky130_fd_sc_hd__o211a_2 _49163_ (.A1(_20274_),
    .A2(_20275_),
    .B1(_20272_),
    .C1(_20270_),
    .X(_20276_));
 sky130_fd_sc_hd__o21ai_4 _49164_ (.A1(_19218_),
    .A2(_19215_),
    .B1(_19210_),
    .Y(_20277_));
 sky130_fd_sc_hd__o21bai_4 _49165_ (.A1(_20273_),
    .A2(_20276_),
    .B1_N(_20277_),
    .Y(_20278_));
 sky130_fd_sc_hd__a21o_1 _49166_ (.A1(_20270_),
    .A2(_20271_),
    .B1(_20272_),
    .X(_20279_));
 sky130_fd_sc_hd__o211ai_1 _49167_ (.A1(_20274_),
    .A2(_20275_),
    .B1(_20272_),
    .C1(_20270_),
    .Y(_20280_));
 sky130_fd_sc_hd__nand3_1 _49168_ (.A(_20277_),
    .B(_20279_),
    .C(_20280_),
    .Y(_20281_));
 sky130_fd_sc_hd__a31o_1 _49169_ (.A1(_19222_),
    .A2(_19223_),
    .A3(_19224_),
    .B1(_19226_),
    .X(_20282_));
 sky130_fd_sc_hd__nand2_2 _49170_ (.A(_19221_),
    .B(_20282_),
    .Y(_20283_));
 sky130_fd_sc_hd__a21o_2 _49171_ (.A1(_20278_),
    .A2(_20281_),
    .B1(_20283_),
    .X(_20284_));
 sky130_fd_sc_hd__nand2_1 _49172_ (.A(_20277_),
    .B(_20280_),
    .Y(_20285_));
 sky130_fd_sc_hd__o211ai_4 _49173_ (.A1(_20285_),
    .A2(_20273_),
    .B1(_20283_),
    .C1(_20278_),
    .Y(_20286_));
 sky130_fd_sc_hd__o211ai_2 _49174_ (.A1(_19847_),
    .A2(_19850_),
    .B1(_20284_),
    .C1(_20286_),
    .Y(_20287_));
 sky130_fd_sc_hd__a21oi_2 _49175_ (.A1(_20278_),
    .A2(_20281_),
    .B1(_20283_),
    .Y(_20288_));
 sky130_fd_sc_hd__o211a_2 _49176_ (.A1(_20285_),
    .A2(_20273_),
    .B1(_20283_),
    .C1(_20278_),
    .X(_20289_));
 sky130_fd_sc_hd__or3b_1 _49177_ (.A(_19845_),
    .B(_19846_),
    .C_N(_19238_),
    .X(_20290_));
 sky130_fd_sc_hd__buf_1 _49178_ (.A(_20290_),
    .X(_20291_));
 sky130_fd_sc_hd__a2bb2o_1 _49179_ (.A1_N(_19845_),
    .A2_N(_19846_),
    .B1(_10635_),
    .B2(_19849_),
    .X(_20292_));
 sky130_fd_sc_hd__nand2_1 _49180_ (.A(_20291_),
    .B(_20292_),
    .Y(_20293_));
 sky130_fd_sc_hd__o21bai_2 _49181_ (.A1(_20288_),
    .A2(_20289_),
    .B1_N(_20293_),
    .Y(_20294_));
 sky130_fd_sc_hd__o21a_2 _49182_ (.A1(_19545_),
    .A2(_19731_),
    .B1(_19732_),
    .X(_20295_));
 sky130_fd_sc_hd__a21oi_2 _49183_ (.A1(_20287_),
    .A2(_20294_),
    .B1(_20295_),
    .Y(_20296_));
 sky130_fd_sc_hd__nand3_2 _49184_ (.A(_20294_),
    .B(_20295_),
    .C(_20287_),
    .Y(_20297_));
 sky130_fd_sc_hd__a21oi_1 _49185_ (.A1(_19241_),
    .A2(_19246_),
    .B1(_19235_),
    .Y(_20298_));
 sky130_fd_sc_hd__nand2_1 _49186_ (.A(_20297_),
    .B(_20298_),
    .Y(_20299_));
 sky130_fd_sc_hd__a21boi_2 _49187_ (.A1(_19261_),
    .A2(_19543_),
    .B1_N(_19735_),
    .Y(_20300_));
 sky130_fd_sc_hd__a21oi_1 _49188_ (.A1(_19533_),
    .A2(_19534_),
    .B1(_19531_),
    .Y(_20301_));
 sky130_fd_sc_hd__buf_1 _49189_ (.A(\delay_line[31][6] ),
    .X(_20302_));
 sky130_fd_sc_hd__buf_1 _49190_ (.A(net317),
    .X(_20303_));
 sky130_fd_sc_hd__and2_1 _49191_ (.A(_20302_),
    .B(_20303_),
    .X(_20304_));
 sky130_fd_sc_hd__o21ai_4 _49192_ (.A1(\delay_line[31][6] ),
    .A2(net317),
    .B1(\delay_line[31][5] ),
    .Y(_20305_));
 sky130_fd_sc_hd__o21ai_2 _49193_ (.A1(_19356_),
    .A2(_19352_),
    .B1(_19353_),
    .Y(_20306_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49194_ (.A(\delay_line[31][5] ),
    .X(_20307_));
 sky130_fd_sc_hd__inv_2 _49195_ (.A(net317),
    .Y(_20308_));
 sky130_fd_sc_hd__nand2_1 _49196_ (.A(_20308_),
    .B(_20302_),
    .Y(_20309_));
 sky130_fd_sc_hd__or2b_1 _49197_ (.A(_19351_),
    .B_N(net317),
    .X(_20310_));
 sky130_fd_sc_hd__nand3b_1 _49198_ (.A_N(_20307_),
    .B(_20309_),
    .C(_20310_),
    .Y(_20311_));
 sky130_fd_sc_hd__o211a_1 _49199_ (.A1(_20304_),
    .A2(_20305_),
    .B1(_20306_),
    .C1(_20311_),
    .X(_20312_));
 sky130_fd_sc_hd__buf_2 _49200_ (.A(_20303_),
    .X(_20313_));
 sky130_fd_sc_hd__a21o_1 _49201_ (.A1(_20302_),
    .A2(_20313_),
    .B1(_20305_),
    .X(_20314_));
 sky130_fd_sc_hd__a21oi_1 _49202_ (.A1(_20311_),
    .A2(_20314_),
    .B1(_20306_),
    .Y(_20315_));
 sky130_fd_sc_hd__o21ai_1 _49203_ (.A1(_20312_),
    .A2(_20315_),
    .B1(_19360_),
    .Y(_20316_));
 sky130_fd_sc_hd__buf_1 _49204_ (.A(\delay_line[31][1] ),
    .X(_20317_));
 sky130_fd_sc_hd__o211ai_2 _49205_ (.A1(_20304_),
    .A2(_20305_),
    .B1(_20306_),
    .C1(_20311_),
    .Y(_20318_));
 sky130_fd_sc_hd__nand3b_1 _49206_ (.A_N(_20315_),
    .B(_19364_),
    .C(_20318_),
    .Y(_20319_));
 sky130_fd_sc_hd__nand3_1 _49207_ (.A(_20316_),
    .B(_20317_),
    .C(_20319_),
    .Y(_20320_));
 sky130_fd_sc_hd__a21o_1 _49208_ (.A1(_20319_),
    .A2(_20316_),
    .B1(_20317_),
    .X(_20321_));
 sky130_fd_sc_hd__nand2_1 _49209_ (.A(_19361_),
    .B(_19367_),
    .Y(_20322_));
 sky130_fd_sc_hd__nand3_1 _49210_ (.A(_20320_),
    .B(_20321_),
    .C(_20322_),
    .Y(_20323_));
 sky130_fd_sc_hd__a21o_1 _49211_ (.A1(_20320_),
    .A2(_20321_),
    .B1(_20322_),
    .X(_20324_));
 sky130_fd_sc_hd__nand4_1 _49212_ (.A(_19369_),
    .B(_19375_),
    .C(_20323_),
    .D(_20324_),
    .Y(_20325_));
 sky130_fd_sc_hd__nand2_1 _49213_ (.A(_20323_),
    .B(_20324_),
    .Y(_20326_));
 sky130_fd_sc_hd__nand2_1 _49214_ (.A(_19369_),
    .B(_19374_),
    .Y(_20327_));
 sky130_fd_sc_hd__nand2_1 _49215_ (.A(_20326_),
    .B(_20327_),
    .Y(_20328_));
 sky130_fd_sc_hd__nand2_1 _49216_ (.A(_20325_),
    .B(_20328_),
    .Y(_20329_));
 sky130_fd_sc_hd__nand2_1 _49217_ (.A(_20329_),
    .B(_19376_),
    .Y(_20330_));
 sky130_fd_sc_hd__inv_2 _49218_ (.A(_20330_),
    .Y(_20331_));
 sky130_fd_sc_hd__clkbuf_2 _49219_ (.A(\delay_line[29][5] ),
    .X(_20332_));
 sky130_fd_sc_hd__nor2_1 _49220_ (.A(_19322_),
    .B(_20332_),
    .Y(_20333_));
 sky130_fd_sc_hd__and2_1 _49221_ (.A(\delay_line[29][4] ),
    .B(\delay_line[29][5] ),
    .X(_20334_));
 sky130_fd_sc_hd__nor3_2 _49222_ (.A(net323),
    .B(_20333_),
    .C(_20334_),
    .Y(_20335_));
 sky130_fd_sc_hd__o21a_1 _49223_ (.A1(_20333_),
    .A2(_20334_),
    .B1(net323),
    .X(_20336_));
 sky130_fd_sc_hd__or4_2 _49224_ (.A(\delay_line[29][0] ),
    .B(_19322_),
    .C(_20335_),
    .D(_20336_),
    .X(_20337_));
 sky130_fd_sc_hd__o22ai_2 _49225_ (.A1(_01051_),
    .A2(_19323_),
    .B1(_20335_),
    .B2(_20336_),
    .Y(_20338_));
 sky130_fd_sc_hd__inv_2 _49226_ (.A(\delay_line[30][7] ),
    .Y(_20339_));
 sky130_fd_sc_hd__buf_1 _49227_ (.A(\delay_line[30][4] ),
    .X(_20340_));
 sky130_fd_sc_hd__or2b_1 _49228_ (.A(_18454_),
    .B_N(_20340_),
    .X(_20341_));
 sky130_fd_sc_hd__inv_2 _49229_ (.A(\delay_line[30][4] ),
    .Y(_20342_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49230_ (.A(_20342_),
    .X(_20343_));
 sky130_fd_sc_hd__nand2_2 _49231_ (.A(_20343_),
    .B(_18454_),
    .Y(_20344_));
 sky130_fd_sc_hd__nand3_2 _49232_ (.A(_20339_),
    .B(_20341_),
    .C(_20344_),
    .Y(_20345_));
 sky130_fd_sc_hd__nor2b_4 _49233_ (.A(_01007_),
    .B_N(_20340_),
    .Y(_20346_));
 sky130_fd_sc_hd__and2b_1 _49234_ (.A_N(_20340_),
    .B(_18454_),
    .X(_20347_));
 sky130_fd_sc_hd__clkbuf_2 _49235_ (.A(\delay_line[30][7] ),
    .X(_20348_));
 sky130_fd_sc_hd__o21ai_2 _49236_ (.A1(_20346_),
    .A2(_20347_),
    .B1(_20348_),
    .Y(_20349_));
 sky130_fd_sc_hd__clkbuf_2 _49237_ (.A(_19328_),
    .X(_20350_));
 sky130_fd_sc_hd__nor2_1 _49238_ (.A(_19332_),
    .B(_19334_),
    .Y(_20351_));
 sky130_fd_sc_hd__o2bb2ai_1 _49239_ (.A1_N(_20345_),
    .A2_N(_20349_),
    .B1(_20350_),
    .B2(_20351_),
    .Y(_20352_));
 sky130_fd_sc_hd__o2111ai_4 _49240_ (.A1(_19332_),
    .A2(_19334_),
    .B1(_19336_),
    .C1(_20345_),
    .D1(_20349_),
    .Y(_20353_));
 sky130_fd_sc_hd__nand3_1 _49241_ (.A(_20352_),
    .B(_19334_),
    .C(_20353_),
    .Y(_20354_));
 sky130_fd_sc_hd__a21o_1 _49242_ (.A1(_20353_),
    .A2(_20352_),
    .B1(_19334_),
    .X(_20355_));
 sky130_fd_sc_hd__a21bo_1 _49243_ (.A1(_19339_),
    .A2(_18455_),
    .B1_N(_19338_),
    .X(_20356_));
 sky130_fd_sc_hd__a21o_1 _49244_ (.A1(_20354_),
    .A2(_20355_),
    .B1(_20356_),
    .X(_20357_));
 sky130_fd_sc_hd__nand3_1 _49245_ (.A(_20356_),
    .B(_20354_),
    .C(_20355_),
    .Y(_20358_));
 sky130_fd_sc_hd__a22oi_1 _49246_ (.A1(_22292_),
    .A2(_01029_),
    .B1(_20357_),
    .B2(_20358_),
    .Y(_20359_));
 sky130_fd_sc_hd__a31o_1 _49247_ (.A1(_22292_),
    .A2(_01040_),
    .A3(_20357_),
    .B1(_20359_),
    .X(_20360_));
 sky130_fd_sc_hd__buf_1 _49248_ (.A(_20360_),
    .X(_20361_));
 sky130_fd_sc_hd__a21bo_1 _49249_ (.A1(_19347_),
    .A2(_19346_),
    .B1_N(_20361_),
    .X(_20362_));
 sky130_fd_sc_hd__nand3b_1 _49250_ (.A_N(_20361_),
    .B(_19346_),
    .C(_19347_),
    .Y(_20363_));
 sky130_fd_sc_hd__nand2_1 _49251_ (.A(_20362_),
    .B(_20363_),
    .Y(_20364_));
 sky130_fd_sc_hd__a21o_1 _49252_ (.A1(_20337_),
    .A2(_20338_),
    .B1(_20364_),
    .X(_20365_));
 sky130_fd_sc_hd__nand3_4 _49253_ (.A(_20337_),
    .B(_20338_),
    .C(_20364_),
    .Y(_20366_));
 sky130_fd_sc_hd__nand2_1 _49254_ (.A(_20365_),
    .B(_20366_),
    .Y(_20367_));
 sky130_fd_sc_hd__a31o_1 _49255_ (.A1(_18481_),
    .A2(_19372_),
    .A3(_19375_),
    .B1(_20329_),
    .X(_20368_));
 sky130_fd_sc_hd__or3b_4 _49256_ (.A(_20331_),
    .B(_20367_),
    .C_N(_20368_),
    .X(_20369_));
 sky130_fd_sc_hd__a21bo_1 _49257_ (.A1(_20368_),
    .A2(_20330_),
    .B1_N(_20367_),
    .X(_20370_));
 sky130_fd_sc_hd__and2_2 _49258_ (.A(_20369_),
    .B(_20370_),
    .X(_20371_));
 sky130_fd_sc_hd__nand3_1 _49259_ (.A(_19288_),
    .B(_18501_),
    .C(_19282_),
    .Y(_20372_));
 sky130_fd_sc_hd__clkbuf_2 _49260_ (.A(\delay_line[27][7] ),
    .X(_20373_));
 sky130_fd_sc_hd__nor2_2 _49261_ (.A(_20373_),
    .B(_19277_),
    .Y(_20374_));
 sky130_fd_sc_hd__nor2_1 _49262_ (.A(net333),
    .B(_20373_),
    .Y(_20375_));
 sky130_fd_sc_hd__and2_1 _49263_ (.A(\delay_line[27][5] ),
    .B(\delay_line[27][7] ),
    .X(_20376_));
 sky130_fd_sc_hd__o21ai_1 _49264_ (.A1(_20375_),
    .A2(_20376_),
    .B1(_19276_),
    .Y(_20377_));
 sky130_fd_sc_hd__nand2_2 _49265_ (.A(_18491_),
    .B(_20373_),
    .Y(_20378_));
 sky130_fd_sc_hd__nand3b_1 _49266_ (.A_N(_20375_),
    .B(_20378_),
    .C(_19279_),
    .Y(_20379_));
 sky130_fd_sc_hd__a21oi_1 _49267_ (.A1(_20377_),
    .A2(_20379_),
    .B1(net274),
    .Y(_20380_));
 sky130_fd_sc_hd__nor3_1 _49268_ (.A(_20374_),
    .B(_24336_),
    .C(_20380_),
    .Y(_20381_));
 sky130_fd_sc_hd__clkbuf_2 _49269_ (.A(_20381_),
    .X(_20382_));
 sky130_fd_sc_hd__o21a_1 _49270_ (.A1(_20380_),
    .A2(_20374_),
    .B1(_24336_),
    .X(_20383_));
 sky130_fd_sc_hd__a21oi_1 _49271_ (.A1(_19281_),
    .A2(_22468_),
    .B1(_19284_),
    .Y(_20384_));
 sky130_fd_sc_hd__o21ai_2 _49272_ (.A1(_20382_),
    .A2(_20383_),
    .B1(_20384_),
    .Y(_20385_));
 sky130_fd_sc_hd__o311a_1 _49273_ (.A1(_19273_),
    .A2(_18496_),
    .A3(_19274_),
    .B1(_22457_),
    .C1(_19281_),
    .X(_20386_));
 sky130_fd_sc_hd__nor2_1 _49274_ (.A(_20381_),
    .B(_20383_),
    .Y(_20387_));
 sky130_fd_sc_hd__o21ai_1 _49275_ (.A1(_19284_),
    .A2(_20386_),
    .B1(_20387_),
    .Y(_20388_));
 sky130_fd_sc_hd__clkbuf_2 _49276_ (.A(_20388_),
    .X(_20389_));
 sky130_fd_sc_hd__nand3b_4 _49277_ (.A_N(_20372_),
    .B(_20385_),
    .C(_20389_),
    .Y(_20390_));
 sky130_fd_sc_hd__a32o_1 _49278_ (.A1(_18501_),
    .A2(_19283_),
    .A3(_19289_),
    .B1(_20385_),
    .B2(_20388_),
    .X(_20391_));
 sky130_fd_sc_hd__a32o_1 _49279_ (.A1(_19291_),
    .A2(_19283_),
    .A3(_19289_),
    .B1(_20390_),
    .B2(_20391_),
    .X(_20392_));
 sky130_fd_sc_hd__and3_1 _49280_ (.A(_19291_),
    .B(_19283_),
    .C(_19289_),
    .X(_20393_));
 sky130_fd_sc_hd__nand3_4 _49281_ (.A(_20391_),
    .B(_20393_),
    .C(_20390_),
    .Y(_20394_));
 sky130_fd_sc_hd__or3b_2 _49282_ (.A(_06469_),
    .B(_24314_),
    .C_N(_19266_),
    .X(_20395_));
 sky130_fd_sc_hd__a21o_1 _49283_ (.A1(_24347_),
    .A2(_19266_),
    .B1(_06590_),
    .X(_20396_));
 sky130_fd_sc_hd__clkbuf_2 _49284_ (.A(\delay_line[26][6] ),
    .X(_20397_));
 sky130_fd_sc_hd__a21o_1 _49285_ (.A1(_20395_),
    .A2(_20396_),
    .B1(_20397_),
    .X(_20398_));
 sky130_fd_sc_hd__nand3_4 _49286_ (.A(_20395_),
    .B(_20396_),
    .C(_20397_),
    .Y(_20399_));
 sky130_fd_sc_hd__a2bb2o_1 _49287_ (.A1_N(_19263_),
    .A2_N(_19265_),
    .B1(_18490_),
    .B2(_19268_),
    .X(_20400_));
 sky130_fd_sc_hd__nand3_2 _49288_ (.A(_20398_),
    .B(_20399_),
    .C(_20400_),
    .Y(_20401_));
 sky130_fd_sc_hd__a21o_1 _49289_ (.A1(_20398_),
    .A2(_20399_),
    .B1(_20400_),
    .X(_20402_));
 sky130_fd_sc_hd__and2_1 _49290_ (.A(_20401_),
    .B(_20402_),
    .X(_20403_));
 sky130_fd_sc_hd__nand3_2 _49291_ (.A(_20392_),
    .B(_20394_),
    .C(_20403_),
    .Y(_20404_));
 sky130_fd_sc_hd__inv_2 _49292_ (.A(_20404_),
    .Y(_20405_));
 sky130_fd_sc_hd__a21oi_1 _49293_ (.A1(_20392_),
    .A2(_20394_),
    .B1(_20403_),
    .Y(_20406_));
 sky130_fd_sc_hd__clkbuf_2 _49294_ (.A(\delay_line[28][7] ),
    .X(_20407_));
 sky130_fd_sc_hd__nand2_1 _49295_ (.A(_18510_),
    .B(_19295_),
    .Y(_20408_));
 sky130_fd_sc_hd__or2b_1 _49296_ (.A(\delay_line[28][7] ),
    .B_N(_19295_),
    .X(_20409_));
 sky130_fd_sc_hd__buf_1 _49297_ (.A(\delay_line[28][7] ),
    .X(_20410_));
 sky130_fd_sc_hd__nand2_1 _49298_ (.A(_19300_),
    .B(_20410_),
    .Y(_20411_));
 sky130_fd_sc_hd__nand3_1 _49299_ (.A(_20408_),
    .B(_20409_),
    .C(_20411_),
    .Y(_20412_));
 sky130_fd_sc_hd__o211ai_2 _49300_ (.A1(_20407_),
    .A2(_20408_),
    .B1(_01117_),
    .C1(_20412_),
    .Y(_20413_));
 sky130_fd_sc_hd__o21ai_1 _49301_ (.A1(_20407_),
    .A2(_20408_),
    .B1(_20412_),
    .Y(_20414_));
 sky130_fd_sc_hd__nand2_1 _49302_ (.A(_15921_),
    .B(_20414_),
    .Y(_20415_));
 sky130_fd_sc_hd__a22o_1 _49303_ (.A1(_19301_),
    .A2(_18513_),
    .B1(_19299_),
    .B2(_24369_),
    .X(_20416_));
 sky130_fd_sc_hd__a21o_1 _49304_ (.A1(_20413_),
    .A2(_20415_),
    .B1(_20416_),
    .X(_20417_));
 sky130_fd_sc_hd__nand3_4 _49305_ (.A(_20416_),
    .B(_20413_),
    .C(_20415_),
    .Y(_20418_));
 sky130_fd_sc_hd__nand3_4 _49306_ (.A(_20417_),
    .B(_24380_),
    .C(_20418_),
    .Y(_20419_));
 sky130_fd_sc_hd__a21o_1 _49307_ (.A1(_20418_),
    .A2(_20417_),
    .B1(_24369_),
    .X(_20420_));
 sky130_fd_sc_hd__nand2_1 _49308_ (.A(_20419_),
    .B(_20420_),
    .Y(_20421_));
 sky130_fd_sc_hd__a21boi_1 _49309_ (.A1(_22259_),
    .A2(_19309_),
    .B1_N(_19307_),
    .Y(_20422_));
 sky130_fd_sc_hd__nand2_1 _49310_ (.A(_20421_),
    .B(_20422_),
    .Y(_20423_));
 sky130_fd_sc_hd__o2111a_1 _49311_ (.A1(_18515_),
    .A2(_18516_),
    .B1(_18509_),
    .C1(_19310_),
    .D1(_19311_),
    .X(_20424_));
 sky130_fd_sc_hd__nand3b_4 _49312_ (.A_N(_20422_),
    .B(_20419_),
    .C(_20420_),
    .Y(_20425_));
 sky130_fd_sc_hd__nand3_1 _49313_ (.A(_20423_),
    .B(_20424_),
    .C(_20425_),
    .Y(_20426_));
 sky130_fd_sc_hd__a2bb2o_1 _49314_ (.A1_N(_18519_),
    .A2_N(_19312_),
    .B1(_20425_),
    .B2(_20423_),
    .X(_20427_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49315_ (.A(_18508_),
    .X(_20428_));
 sky130_fd_sc_hd__and4b_1 _49316_ (.A_N(_15954_),
    .B(_18521_),
    .C(_18518_),
    .D(_20428_),
    .X(_20429_));
 sky130_fd_sc_hd__nor2_1 _49317_ (.A(_18522_),
    .B(_19312_),
    .Y(_20430_));
 sky130_fd_sc_hd__a221o_1 _49318_ (.A1(_20426_),
    .A2(_20427_),
    .B1(_20429_),
    .B2(_19315_),
    .C1(_20430_),
    .X(_20431_));
 sky130_fd_sc_hd__nand3_1 _49319_ (.A(_20423_),
    .B(_20430_),
    .C(_20425_),
    .Y(_20432_));
 sky130_fd_sc_hd__inv_2 _49320_ (.A(_20418_),
    .Y(_20433_));
 sky130_fd_sc_hd__nand2_1 _49321_ (.A(_20429_),
    .B(_20433_),
    .Y(_20434_));
 sky130_fd_sc_hd__and3_1 _49322_ (.A(_20431_),
    .B(_20432_),
    .C(_20434_),
    .X(_20435_));
 sky130_fd_sc_hd__or3b_2 _49323_ (.A(_20405_),
    .B(_20406_),
    .C_N(_20435_),
    .X(_20436_));
 sky130_fd_sc_hd__o21bai_1 _49324_ (.A1(_20405_),
    .A2(_20406_),
    .B1_N(_20435_),
    .Y(_20437_));
 sky130_fd_sc_hd__nand2_1 _49325_ (.A(_20436_),
    .B(_20437_),
    .Y(_20438_));
 sky130_fd_sc_hd__o21ba_1 _49326_ (.A1(_19293_),
    .A2(_19316_),
    .B1_N(_19294_),
    .X(_20439_));
 sky130_fd_sc_hd__and2_1 _49327_ (.A(_20438_),
    .B(_20439_),
    .X(_20440_));
 sky130_fd_sc_hd__nor2_1 _49328_ (.A(_20439_),
    .B(_20438_),
    .Y(_20441_));
 sky130_fd_sc_hd__nor2_2 _49329_ (.A(_20440_),
    .B(_20441_),
    .Y(_20442_));
 sky130_fd_sc_hd__xnor2_4 _49330_ (.A(_20371_),
    .B(_20442_),
    .Y(_20443_));
 sky130_fd_sc_hd__or2_1 _49331_ (.A(_20301_),
    .B(_20443_),
    .X(_20444_));
 sky130_fd_sc_hd__nand2_1 _49332_ (.A(_20443_),
    .B(_20301_),
    .Y(_20445_));
 sky130_fd_sc_hd__a211oi_1 _49333_ (.A1(_20444_),
    .A2(_20445_),
    .B1(_19321_),
    .C1(net114),
    .Y(_20446_));
 sky130_fd_sc_hd__inv_2 _49334_ (.A(_20446_),
    .Y(_20447_));
 sky130_fd_sc_hd__o211ai_2 _49335_ (.A1(_19321_),
    .A2(net114),
    .B1(_20444_),
    .C1(_20445_),
    .Y(_20448_));
 sky130_fd_sc_hd__buf_1 _49336_ (.A(\delay_line[22][6] ),
    .X(_20449_));
 sky130_fd_sc_hd__clkbuf_2 _49337_ (.A(_20449_),
    .X(_20450_));
 sky130_fd_sc_hd__xor2_2 _49338_ (.A(_06865_),
    .B(_20450_),
    .X(_20451_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49339_ (.A(_20451_),
    .X(_20452_));
 sky130_fd_sc_hd__o21a_1 _49340_ (.A1(_19504_),
    .A2(_19506_),
    .B1(_20452_),
    .X(_20453_));
 sky130_fd_sc_hd__clkbuf_2 _49341_ (.A(_19502_),
    .X(_20454_));
 sky130_fd_sc_hd__a211oi_1 _49342_ (.A1(_01424_),
    .A2(_20454_),
    .B1(_19507_),
    .C1(_20452_),
    .Y(_20455_));
 sky130_fd_sc_hd__a211oi_4 _49343_ (.A1(_18308_),
    .A2(_18313_),
    .B1(_19517_),
    .C1(_19520_),
    .Y(_20456_));
 sky130_fd_sc_hd__o21ai_4 _49344_ (.A1(net346),
    .A2(_19510_),
    .B1(_19511_),
    .Y(_20457_));
 sky130_fd_sc_hd__buf_1 _49345_ (.A(\delay_line[24][3] ),
    .X(_20458_));
 sky130_fd_sc_hd__o21bai_1 _49346_ (.A1(_19510_),
    .A2(_19514_),
    .B1_N(_20458_),
    .Y(_20459_));
 sky130_fd_sc_hd__or2_1 _49347_ (.A(\delay_line[24][1] ),
    .B(net344),
    .X(_20460_));
 sky130_fd_sc_hd__nand2_1 _49348_ (.A(_01435_),
    .B(_06898_),
    .Y(_20461_));
 sky130_fd_sc_hd__nand3_1 _49349_ (.A(_20460_),
    .B(_20458_),
    .C(_20461_),
    .Y(_20462_));
 sky130_fd_sc_hd__clkbuf_2 _49350_ (.A(\delay_line[24][6] ),
    .X(_20463_));
 sky130_fd_sc_hd__clkbuf_2 _49351_ (.A(_20463_),
    .X(_20464_));
 sky130_fd_sc_hd__nand3_1 _49352_ (.A(_20459_),
    .B(_20462_),
    .C(_20464_),
    .Y(_20465_));
 sky130_fd_sc_hd__buf_1 _49353_ (.A(_20465_),
    .X(_20466_));
 sky130_fd_sc_hd__inv_2 _49354_ (.A(_20463_),
    .Y(_20467_));
 sky130_fd_sc_hd__o21ai_1 _49355_ (.A1(_19510_),
    .A2(_19514_),
    .B1(_17007_),
    .Y(_20468_));
 sky130_fd_sc_hd__nand3b_1 _49356_ (.A_N(_17007_),
    .B(_20461_),
    .C(_20460_),
    .Y(_20469_));
 sky130_fd_sc_hd__nand3_1 _49357_ (.A(_20467_),
    .B(_20468_),
    .C(_20469_),
    .Y(_20470_));
 sky130_fd_sc_hd__and3_1 _49358_ (.A(_19516_),
    .B(_20466_),
    .C(_20470_),
    .X(_20471_));
 sky130_fd_sc_hd__a21oi_1 _49359_ (.A1(_20466_),
    .A2(_20470_),
    .B1(_19517_),
    .Y(_20472_));
 sky130_fd_sc_hd__nor2_1 _49360_ (.A(_20471_),
    .B(_20472_),
    .Y(_20473_));
 sky130_fd_sc_hd__xnor2_2 _49361_ (.A(_20457_),
    .B(_20473_),
    .Y(_20474_));
 sky130_fd_sc_hd__buf_1 _49362_ (.A(_20474_),
    .X(_20475_));
 sky130_fd_sc_hd__o21a_1 _49363_ (.A1(_20456_),
    .A2(_19524_),
    .B1(_20475_),
    .X(_20476_));
 sky130_fd_sc_hd__or3_1 _49364_ (.A(_20456_),
    .B(_19524_),
    .C(_20475_),
    .X(_20477_));
 sky130_fd_sc_hd__or4b_1 _49365_ (.A(_20453_),
    .B(_20455_),
    .C(_20476_),
    .D_N(_20477_),
    .X(_20478_));
 sky130_fd_sc_hd__inv_2 _49366_ (.A(_20476_),
    .Y(_20479_));
 sky130_fd_sc_hd__a2bb2o_1 _49367_ (.A1_N(_20453_),
    .A2_N(_20455_),
    .B1(_20479_),
    .B2(_20477_),
    .X(_20480_));
 sky130_fd_sc_hd__a211oi_2 _49368_ (.A1(_18327_),
    .A2(_18331_),
    .B1(_19493_),
    .C1(_19494_),
    .Y(_20481_));
 sky130_fd_sc_hd__nor2_1 _49369_ (.A(_18333_),
    .B(_19497_),
    .Y(_20482_));
 sky130_fd_sc_hd__clkbuf_2 _49370_ (.A(\delay_line[25][7] ),
    .X(_20483_));
 sky130_fd_sc_hd__nand2b_2 _49371_ (.A_N(_20483_),
    .B(_18323_),
    .Y(_20484_));
 sky130_fd_sc_hd__or2b_1 _49372_ (.A(_18323_),
    .B_N(\delay_line[25][7] ),
    .X(_20485_));
 sky130_fd_sc_hd__nand3_1 _49373_ (.A(_19491_),
    .B(_20484_),
    .C(_20485_),
    .Y(_20486_));
 sky130_fd_sc_hd__a21o_1 _49374_ (.A1(_20484_),
    .A2(_20485_),
    .B1(_19491_),
    .X(_20487_));
 sky130_fd_sc_hd__a21oi_1 _49375_ (.A1(_20486_),
    .A2(_20487_),
    .B1(_17226_),
    .Y(_20488_));
 sky130_fd_sc_hd__nand3_1 _49376_ (.A(_20487_),
    .B(_17226_),
    .C(_20486_),
    .Y(_20489_));
 sky130_fd_sc_hd__a21bo_1 _49377_ (.A1(_19490_),
    .A2(_23731_),
    .B1_N(_19492_),
    .X(_20490_));
 sky130_fd_sc_hd__nand3b_2 _49378_ (.A_N(_20488_),
    .B(_20489_),
    .C(_20490_),
    .Y(_20491_));
 sky130_fd_sc_hd__and3_1 _49379_ (.A(_20487_),
    .B(_17139_),
    .C(_20486_),
    .X(_20492_));
 sky130_fd_sc_hd__o21bai_2 _49380_ (.A1(_20488_),
    .A2(_20492_),
    .B1_N(_20490_),
    .Y(_20493_));
 sky130_fd_sc_hd__nand3_2 _49381_ (.A(_20491_),
    .B(_20493_),
    .C(_22358_),
    .Y(_20494_));
 sky130_fd_sc_hd__a21o_1 _49382_ (.A1(_20491_),
    .A2(_20493_),
    .B1(_22369_),
    .X(_20495_));
 sky130_fd_sc_hd__and2_1 _49383_ (.A(_20494_),
    .B(_20495_),
    .X(_20496_));
 sky130_fd_sc_hd__o21ai_1 _49384_ (.A1(_20481_),
    .A2(_20482_),
    .B1(_20496_),
    .Y(_20497_));
 sky130_fd_sc_hd__nand2_1 _49385_ (.A(_20494_),
    .B(_20495_),
    .Y(_20498_));
 sky130_fd_sc_hd__o211ai_1 _49386_ (.A1(_18333_),
    .A2(_19497_),
    .B1(_20498_),
    .C1(_19496_),
    .Y(_20499_));
 sky130_fd_sc_hd__inv_2 _49387_ (.A(_19497_),
    .Y(_20500_));
 sky130_fd_sc_hd__nand4_1 _49388_ (.A(_20497_),
    .B(_20499_),
    .C(_19498_),
    .D(_20500_),
    .Y(_20501_));
 sky130_fd_sc_hd__clkbuf_2 _49389_ (.A(_20501_),
    .X(_20502_));
 sky130_fd_sc_hd__a32o_1 _49390_ (.A1(_19498_),
    .A2(_19495_),
    .A3(_19496_),
    .B1(_20497_),
    .B2(_20499_),
    .X(_20503_));
 sky130_fd_sc_hd__and4_1 _49391_ (.A(_20478_),
    .B(_20480_),
    .C(_20502_),
    .D(_20503_),
    .X(_20504_));
 sky130_fd_sc_hd__a22oi_2 _49392_ (.A1(_20478_),
    .A2(_20480_),
    .B1(_20502_),
    .B2(_20503_),
    .Y(_20505_));
 sky130_fd_sc_hd__o211a_1 _49393_ (.A1(_20504_),
    .A2(_20505_),
    .B1(_19415_),
    .C1(_19430_),
    .X(_20506_));
 sky130_fd_sc_hd__a211oi_2 _49394_ (.A1(_19415_),
    .A2(_19430_),
    .B1(_20504_),
    .C1(_20505_),
    .Y(_20507_));
 sky130_fd_sc_hd__nor2_1 _49395_ (.A(_20506_),
    .B(_20507_),
    .Y(_20508_));
 sky130_fd_sc_hd__o21ai_1 _49396_ (.A1(_19529_),
    .A2(_19500_),
    .B1(_19526_),
    .Y(_20509_));
 sky130_fd_sc_hd__and2_1 _49397_ (.A(_20508_),
    .B(_20509_),
    .X(_20510_));
 sky130_fd_sc_hd__o221a_1 _49398_ (.A1(_19529_),
    .A2(_19500_),
    .B1(_20507_),
    .B2(_20506_),
    .C1(_19526_),
    .X(_20511_));
 sky130_fd_sc_hd__or2_1 _49399_ (.A(_20510_),
    .B(_20511_),
    .X(_20512_));
 sky130_fd_sc_hd__and2_2 _49400_ (.A(_19417_),
    .B(\delay_line[21][6] ),
    .X(_20513_));
 sky130_fd_sc_hd__buf_1 _49401_ (.A(\delay_line[21][6] ),
    .X(_20514_));
 sky130_fd_sc_hd__nor2_1 _49402_ (.A(_19417_),
    .B(_20514_),
    .Y(_20515_));
 sky130_fd_sc_hd__nand2_1 _49403_ (.A(net360),
    .B(\delay_line[21][5] ),
    .Y(_20516_));
 sky130_fd_sc_hd__clkbuf_4 _49404_ (.A(_20516_),
    .X(_20517_));
 sky130_fd_sc_hd__o21ai_4 _49405_ (.A1(_20513_),
    .A2(_20515_),
    .B1(_20517_),
    .Y(_20518_));
 sky130_fd_sc_hd__or2_1 _49406_ (.A(_20514_),
    .B(_20516_),
    .X(_20519_));
 sky130_fd_sc_hd__a21o_1 _49407_ (.A1(_20518_),
    .A2(_20519_),
    .B1(_01600_),
    .X(_20520_));
 sky130_fd_sc_hd__clkbuf_2 _49408_ (.A(\delay_line[21][6] ),
    .X(_20521_));
 sky130_fd_sc_hd__o211ai_4 _49409_ (.A1(_20521_),
    .A2(_20517_),
    .B1(_01600_),
    .C1(_20518_),
    .Y(_20522_));
 sky130_fd_sc_hd__nand2_1 _49410_ (.A(_19421_),
    .B(_19423_),
    .Y(_20523_));
 sky130_fd_sc_hd__a21o_1 _49411_ (.A1(_20520_),
    .A2(_20522_),
    .B1(_20523_),
    .X(_20524_));
 sky130_fd_sc_hd__nand3_2 _49412_ (.A(_20523_),
    .B(_20520_),
    .C(_20522_),
    .Y(_20525_));
 sky130_fd_sc_hd__nand3_2 _49413_ (.A(_20524_),
    .B(_23995_),
    .C(_20525_),
    .Y(_20526_));
 sky130_fd_sc_hd__a21o_1 _49414_ (.A1(_20525_),
    .A2(_20524_),
    .B1(_24006_),
    .X(_20527_));
 sky130_fd_sc_hd__and2_1 _49415_ (.A(_16503_),
    .B(_07305_),
    .X(_20528_));
 sky130_fd_sc_hd__and4b_2 _49416_ (.A_N(_18349_),
    .B(_19422_),
    .C(_19423_),
    .D(_20528_),
    .X(_20529_));
 sky130_fd_sc_hd__and4_1 _49417_ (.A(_19422_),
    .B(_19423_),
    .C(_18349_),
    .D(_18354_),
    .X(_20530_));
 sky130_fd_sc_hd__a211o_1 _49418_ (.A1(_20526_),
    .A2(_20527_),
    .B1(_20529_),
    .C1(_20530_),
    .X(_20531_));
 sky130_fd_sc_hd__inv_2 _49419_ (.A(_20526_),
    .Y(_20532_));
 sky130_fd_sc_hd__a21oi_1 _49420_ (.A1(_20525_),
    .A2(_20524_),
    .B1(_07338_),
    .Y(_20533_));
 sky130_fd_sc_hd__nor2_1 _49421_ (.A(_20532_),
    .B(_20533_),
    .Y(_20534_));
 sky130_fd_sc_hd__o21ai_1 _49422_ (.A1(_20529_),
    .A2(_20530_),
    .B1(_20534_),
    .Y(_20535_));
 sky130_fd_sc_hd__nand2_1 _49423_ (.A(_19424_),
    .B(_19425_),
    .Y(_20536_));
 sky130_fd_sc_hd__nor2_1 _49424_ (.A(_18365_),
    .B(_20536_),
    .Y(_20537_));
 sky130_fd_sc_hd__and3_2 _49425_ (.A(_20531_),
    .B(_20535_),
    .C(_20537_),
    .X(_20538_));
 sky130_fd_sc_hd__o2bb2a_1 _49426_ (.A1_N(_20531_),
    .A2_N(_20535_),
    .B1(_18366_),
    .B2(_20536_),
    .X(_20539_));
 sky130_fd_sc_hd__nor2_1 _49427_ (.A(_20538_),
    .B(_20539_),
    .Y(_20540_));
 sky130_fd_sc_hd__nor4_1 _49428_ (.A(_23940_),
    .B(_18388_),
    .C(_19392_),
    .D(_19396_),
    .Y(_20541_));
 sky130_fd_sc_hd__clkbuf_2 _49429_ (.A(\delay_line[18][6] ),
    .X(_20542_));
 sky130_fd_sc_hd__xor2_2 _49430_ (.A(_07514_),
    .B(_20542_),
    .X(_20543_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49431_ (.A(_20543_),
    .X(_20544_));
 sky130_fd_sc_hd__or3_2 _49432_ (.A(_19397_),
    .B(net260),
    .C(_20544_),
    .X(_20545_));
 sky130_fd_sc_hd__o21ai_2 _49433_ (.A1(_19397_),
    .A2(net260),
    .B1(_20544_),
    .Y(_20546_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49434_ (.A(\delay_line[19][6] ),
    .X(_20547_));
 sky130_fd_sc_hd__and2_2 _49435_ (.A(\delay_line[19][5] ),
    .B(_20547_),
    .X(_20548_));
 sky130_fd_sc_hd__nor2_1 _49436_ (.A(_19402_),
    .B(_20547_),
    .Y(_20549_));
 sky130_fd_sc_hd__nand2_1 _49437_ (.A(net371),
    .B(_19402_),
    .Y(_20550_));
 sky130_fd_sc_hd__o21ai_2 _49438_ (.A1(_20548_),
    .A2(_20549_),
    .B1(_20550_),
    .Y(_20551_));
 sky130_fd_sc_hd__clkbuf_2 _49439_ (.A(_20551_),
    .X(_20552_));
 sky130_fd_sc_hd__inv_2 _49440_ (.A(_20547_),
    .Y(_20553_));
 sky130_fd_sc_hd__nand2_2 _49441_ (.A(_19401_),
    .B(_20553_),
    .Y(_20554_));
 sky130_fd_sc_hd__a21oi_1 _49442_ (.A1(_20552_),
    .A2(_20554_),
    .B1(_07371_),
    .Y(_20555_));
 sky130_fd_sc_hd__and3_1 _49443_ (.A(_20551_),
    .B(_20554_),
    .C(_07360_),
    .X(_20556_));
 sky130_fd_sc_hd__a21boi_1 _49444_ (.A1(_19404_),
    .A2(_23874_),
    .B1_N(_19406_),
    .Y(_20557_));
 sky130_fd_sc_hd__o21ai_2 _49445_ (.A1(_20555_),
    .A2(_20556_),
    .B1(_20557_),
    .Y(_20558_));
 sky130_fd_sc_hd__a21o_1 _49446_ (.A1(_20551_),
    .A2(_20554_),
    .B1(_07360_),
    .X(_20559_));
 sky130_fd_sc_hd__buf_2 _49447_ (.A(_20547_),
    .X(_20560_));
 sky130_fd_sc_hd__clkbuf_2 _49448_ (.A(_20560_),
    .X(_20561_));
 sky130_fd_sc_hd__o211ai_1 _49449_ (.A1(_20561_),
    .A2(_20550_),
    .B1(_07360_),
    .C1(_20552_),
    .Y(_20562_));
 sky130_fd_sc_hd__nand3b_2 _49450_ (.A_N(_20557_),
    .B(_20559_),
    .C(_20562_),
    .Y(_20563_));
 sky130_fd_sc_hd__nand3_1 _49451_ (.A(_20558_),
    .B(_23885_),
    .C(_20563_),
    .Y(_20564_));
 sky130_fd_sc_hd__buf_1 _49452_ (.A(_20564_),
    .X(_20565_));
 sky130_fd_sc_hd__a21o_1 _49453_ (.A1(_20563_),
    .A2(_20558_),
    .B1(_23896_),
    .X(_20566_));
 sky130_fd_sc_hd__clkbuf_2 _49454_ (.A(_19409_),
    .X(_20567_));
 sky130_fd_sc_hd__a221o_1 _49455_ (.A1(_20565_),
    .A2(_20566_),
    .B1(_18381_),
    .B2(_19412_),
    .C1(_20567_),
    .X(_20568_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49456_ (.A(_18376_),
    .X(_20569_));
 sky130_fd_sc_hd__and4_2 _49457_ (.A(_19407_),
    .B(_19408_),
    .C(_20569_),
    .D(_18369_),
    .X(_20570_));
 sky130_fd_sc_hd__and2_1 _49458_ (.A(_20565_),
    .B(_20566_),
    .X(_20571_));
 sky130_fd_sc_hd__o21ai_2 _49459_ (.A1(_20567_),
    .A2(_20570_),
    .B1(_20571_),
    .Y(_20572_));
 sky130_fd_sc_hd__nand4_4 _49460_ (.A(_20568_),
    .B(_18379_),
    .C(_20572_),
    .D(_19412_),
    .Y(_20573_));
 sky130_fd_sc_hd__clkbuf_2 _49461_ (.A(_20569_),
    .X(_20574_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49462_ (.A(_18380_),
    .X(_20575_));
 sky130_fd_sc_hd__or4b_1 _49463_ (.A(_07470_),
    .B(_20574_),
    .C(_07437_),
    .D_N(_20575_),
    .X(_20576_));
 sky130_fd_sc_hd__or2_1 _49464_ (.A(_20567_),
    .B(_19411_),
    .X(_20577_));
 sky130_fd_sc_hd__a2bb2o_1 _49465_ (.A1_N(_20576_),
    .A2_N(_20577_),
    .B1(_20572_),
    .B2(_20568_),
    .X(_20578_));
 sky130_fd_sc_hd__nand4_4 _49466_ (.A(_20545_),
    .B(_20546_),
    .C(_20573_),
    .D(_20578_),
    .Y(_20579_));
 sky130_fd_sc_hd__a22o_1 _49467_ (.A1(_20545_),
    .A2(_20546_),
    .B1(_20573_),
    .B2(_20578_),
    .X(_20580_));
 sky130_fd_sc_hd__nand2_1 _49468_ (.A(_20579_),
    .B(_20580_),
    .Y(_20581_));
 sky130_fd_sc_hd__xnor2_1 _49469_ (.A(_20540_),
    .B(_20581_),
    .Y(_20582_));
 sky130_fd_sc_hd__nor3b_4 _49470_ (.A(_19448_),
    .B(_19449_),
    .C_N(_19451_),
    .Y(_20583_));
 sky130_fd_sc_hd__buf_1 _49471_ (.A(\delay_line[14][2] ),
    .X(_20584_));
 sky130_fd_sc_hd__nor2_1 _49472_ (.A(net393),
    .B(_20584_),
    .Y(_20585_));
 sky130_fd_sc_hd__and2_1 _49473_ (.A(\delay_line[14][1] ),
    .B(\delay_line[14][2] ),
    .X(_20586_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49474_ (.A(\delay_line[14][6] ),
    .X(_20587_));
 sky130_fd_sc_hd__or3b_4 _49475_ (.A(_20585_),
    .B(_20586_),
    .C_N(_20587_),
    .X(_20588_));
 sky130_fd_sc_hd__buf_1 _49476_ (.A(_20587_),
    .X(_20589_));
 sky130_fd_sc_hd__o21bai_4 _49477_ (.A1(_20585_),
    .A2(_20586_),
    .B1_N(_20589_),
    .Y(_20590_));
 sky130_fd_sc_hd__o211a_1 _49478_ (.A1(_19449_),
    .A2(_20583_),
    .B1(_20588_),
    .C1(_20590_),
    .X(_20591_));
 sky130_fd_sc_hd__a221oi_4 _49479_ (.A1(_24061_),
    .A2(_01765_),
    .B1(_20588_),
    .B2(_20590_),
    .C1(_20583_),
    .Y(_20592_));
 sky130_fd_sc_hd__nor3_2 _49480_ (.A(_19455_),
    .B(_20591_),
    .C(_20592_),
    .Y(_20593_));
 sky130_fd_sc_hd__o21a_1 _49481_ (.A1(_20591_),
    .A2(_20592_),
    .B1(_19455_),
    .X(_20594_));
 sky130_fd_sc_hd__nand3_1 _49482_ (.A(net183),
    .B(_19469_),
    .C(_19470_),
    .Y(_20595_));
 sky130_fd_sc_hd__inv_2 _49483_ (.A(\delay_line[15][7] ),
    .Y(_20596_));
 sky130_fd_sc_hd__nand2_1 _49484_ (.A(_20596_),
    .B(_18416_),
    .Y(_20597_));
 sky130_fd_sc_hd__inv_2 _49485_ (.A(\delay_line[15][5] ),
    .Y(_20598_));
 sky130_fd_sc_hd__buf_1 _49486_ (.A(\delay_line[15][7] ),
    .X(_20599_));
 sky130_fd_sc_hd__buf_2 _49487_ (.A(_20599_),
    .X(_20600_));
 sky130_fd_sc_hd__nand2_1 _49488_ (.A(_20598_),
    .B(_20600_),
    .Y(_20601_));
 sky130_fd_sc_hd__nand3_1 _49489_ (.A(_19462_),
    .B(_20597_),
    .C(_20601_),
    .Y(_20602_));
 sky130_fd_sc_hd__and2b_1 _49490_ (.A_N(_20599_),
    .B(_18414_),
    .X(_20603_));
 sky130_fd_sc_hd__nor2_1 _49491_ (.A(_18414_),
    .B(_20596_),
    .Y(_20604_));
 sky130_fd_sc_hd__o21ai_2 _49492_ (.A1(_20603_),
    .A2(_20604_),
    .B1(_19458_),
    .Y(_20605_));
 sky130_fd_sc_hd__buf_1 _49493_ (.A(_01787_),
    .X(_20606_));
 sky130_fd_sc_hd__a21oi_1 _49494_ (.A1(_20602_),
    .A2(_20605_),
    .B1(_20606_),
    .Y(_20607_));
 sky130_fd_sc_hd__and3_1 _49495_ (.A(_20605_),
    .B(_20606_),
    .C(_20602_),
    .X(_20608_));
 sky130_fd_sc_hd__a21bo_1 _49496_ (.A1(_19460_),
    .A2(\delay_line[15][1] ),
    .B1_N(_19463_),
    .X(_20609_));
 sky130_fd_sc_hd__o21bai_1 _49497_ (.A1(_20607_),
    .A2(_20608_),
    .B1_N(_20609_),
    .Y(_20610_));
 sky130_fd_sc_hd__nand3_1 _49498_ (.A(_20605_),
    .B(_20606_),
    .C(_20602_),
    .Y(_20611_));
 sky130_fd_sc_hd__nand3b_2 _49499_ (.A_N(_20607_),
    .B(_20611_),
    .C(_20609_),
    .Y(_20612_));
 sky130_fd_sc_hd__nand3_2 _49500_ (.A(_20610_),
    .B(_22402_),
    .C(_20612_),
    .Y(_20613_));
 sky130_fd_sc_hd__a21o_1 _49501_ (.A1(_20612_),
    .A2(_20610_),
    .B1(_22413_),
    .X(_20614_));
 sky130_fd_sc_hd__nand2_1 _49502_ (.A(_20613_),
    .B(_20614_),
    .Y(_20615_));
 sky130_fd_sc_hd__a21o_1 _49503_ (.A1(_19470_),
    .A2(_20595_),
    .B1(_20615_),
    .X(_20616_));
 sky130_fd_sc_hd__nor2_2 _49504_ (.A(_18432_),
    .B(_19472_),
    .Y(_20617_));
 sky130_fd_sc_hd__o211ai_2 _49505_ (.A1(_18431_),
    .A2(_19471_),
    .B1(_20615_),
    .C1(_19470_),
    .Y(_20618_));
 sky130_fd_sc_hd__and3_1 _49506_ (.A(_20616_),
    .B(_20617_),
    .C(_20618_),
    .X(_20619_));
 sky130_fd_sc_hd__a2bb2o_1 _49507_ (.A1_N(_18432_),
    .A2_N(_19472_),
    .B1(_20618_),
    .B2(_20616_),
    .X(_20620_));
 sky130_fd_sc_hd__or4b_2 _49508_ (.A(_20593_),
    .B(_20594_),
    .C(_20619_),
    .D_N(_20620_),
    .X(_20621_));
 sky130_fd_sc_hd__nand3_1 _49509_ (.A(_20616_),
    .B(_20617_),
    .C(_20618_),
    .Y(_20622_));
 sky130_fd_sc_hd__a2bb2oi_1 _49510_ (.A1_N(_20593_),
    .A2_N(_20594_),
    .B1(_20622_),
    .B2(_20620_),
    .Y(_20623_));
 sky130_fd_sc_hd__inv_2 _49511_ (.A(_20623_),
    .Y(_20624_));
 sky130_fd_sc_hd__o21ai_2 _49512_ (.A1(_24127_),
    .A2(_19433_),
    .B1(_19434_),
    .Y(_20625_));
 sky130_fd_sc_hd__o21ai_1 _49513_ (.A1(_19432_),
    .A2(_19436_),
    .B1(_16667_),
    .Y(_20626_));
 sky130_fd_sc_hd__or2_1 _49514_ (.A(\delay_line[16][1] ),
    .B(\delay_line[16][2] ),
    .X(_20627_));
 sky130_fd_sc_hd__nand2_1 _49515_ (.A(_01864_),
    .B(_07206_),
    .Y(_20628_));
 sky130_fd_sc_hd__nand3_1 _49516_ (.A(_20627_),
    .B(_16656_),
    .C(_20628_),
    .Y(_20629_));
 sky130_fd_sc_hd__clkbuf_2 _49517_ (.A(net385),
    .X(_20630_));
 sky130_fd_sc_hd__nand3_1 _49518_ (.A(_20626_),
    .B(_20629_),
    .C(_20630_),
    .Y(_20631_));
 sky130_fd_sc_hd__buf_1 _49519_ (.A(_20631_),
    .X(_20632_));
 sky130_fd_sc_hd__o21ai_1 _49520_ (.A1(_19433_),
    .A2(_19437_),
    .B1(_16590_),
    .Y(_20633_));
 sky130_fd_sc_hd__nand3_1 _49521_ (.A(_16667_),
    .B(_20628_),
    .C(_20627_),
    .Y(_20634_));
 sky130_fd_sc_hd__nand3b_1 _49522_ (.A_N(_20630_),
    .B(_20633_),
    .C(_20634_),
    .Y(_20635_));
 sky130_fd_sc_hd__and3_1 _49523_ (.A(_19439_),
    .B(_20632_),
    .C(_20635_),
    .X(_20636_));
 sky130_fd_sc_hd__a21oi_1 _49524_ (.A1(_20632_),
    .A2(_20635_),
    .B1(_19439_),
    .Y(_20637_));
 sky130_fd_sc_hd__nor2_1 _49525_ (.A(_20636_),
    .B(_20637_),
    .Y(_20638_));
 sky130_fd_sc_hd__xnor2_2 _49526_ (.A(_20625_),
    .B(_20638_),
    .Y(_20639_));
 sky130_fd_sc_hd__o21ai_1 _49527_ (.A1(_19446_),
    .A2(_19445_),
    .B1(_20639_),
    .Y(_20640_));
 sky130_fd_sc_hd__or3_1 _49528_ (.A(_19446_),
    .B(_19445_),
    .C(_20639_),
    .X(_20641_));
 sky130_fd_sc_hd__and2_1 _49529_ (.A(_20640_),
    .B(_20641_),
    .X(_20642_));
 sky130_fd_sc_hd__nand3_1 _49530_ (.A(_20621_),
    .B(_20624_),
    .C(_20642_),
    .Y(_20643_));
 sky130_fd_sc_hd__a21o_1 _49531_ (.A1(_20621_),
    .A2(_20624_),
    .B1(_20642_),
    .X(_20644_));
 sky130_fd_sc_hd__and2_1 _49532_ (.A(_20643_),
    .B(_20644_),
    .X(_20645_));
 sky130_fd_sc_hd__nor3_4 _49533_ (.A(_19475_),
    .B(_19478_),
    .C(_20645_),
    .Y(_20646_));
 sky130_fd_sc_hd__o21a_2 _49534_ (.A1(_19475_),
    .A2(_19478_),
    .B1(_20645_),
    .X(_20647_));
 sky130_fd_sc_hd__nor2_1 _49535_ (.A(_20646_),
    .B(_20647_),
    .Y(_20648_));
 sky130_fd_sc_hd__and2_1 _49536_ (.A(_20582_),
    .B(_20648_),
    .X(_20649_));
 sky130_fd_sc_hd__nor2_1 _49537_ (.A(_20582_),
    .B(_20648_),
    .Y(_20650_));
 sky130_fd_sc_hd__or2_1 _49538_ (.A(_20649_),
    .B(_20650_),
    .X(_20651_));
 sky130_fd_sc_hd__or3b_1 _49539_ (.A(_19483_),
    .B(net105),
    .C_N(_20651_),
    .X(_20652_));
 sky130_fd_sc_hd__o21bai_4 _49540_ (.A1(_19483_),
    .A2(net105),
    .B1_N(_20651_),
    .Y(_20653_));
 sky130_fd_sc_hd__nand2_2 _49541_ (.A(_20652_),
    .B(_20653_),
    .Y(_20654_));
 sky130_fd_sc_hd__or2_1 _49542_ (.A(_20512_),
    .B(_20654_),
    .X(_20655_));
 sky130_fd_sc_hd__nand2_1 _49543_ (.A(_20512_),
    .B(_20654_),
    .Y(_20656_));
 sky130_fd_sc_hd__a211o_1 _49544_ (.A1(_20655_),
    .A2(_20656_),
    .B1(_19486_),
    .C1(net96),
    .X(_20657_));
 sky130_fd_sc_hd__o211ai_2 _49545_ (.A1(_19486_),
    .A2(net96),
    .B1(_20655_),
    .C1(_20656_),
    .Y(_20658_));
 sky130_fd_sc_hd__nand4_1 _49546_ (.A(_20447_),
    .B(_20448_),
    .C(_20657_),
    .D(_20658_),
    .Y(_20659_));
 sky130_fd_sc_hd__a22o_1 _49547_ (.A1(_20447_),
    .A2(_20448_),
    .B1(_20657_),
    .B2(_20658_),
    .X(_20660_));
 sky130_fd_sc_hd__nand2_1 _49548_ (.A(_20659_),
    .B(_20660_),
    .Y(_20661_));
 sky130_fd_sc_hd__a21oi_1 _49549_ (.A1(_19388_),
    .A2(_19542_),
    .B1(_19541_),
    .Y(_20662_));
 sky130_fd_sc_hd__xnor2_1 _49550_ (.A(_20661_),
    .B(_20662_),
    .Y(_20663_));
 sky130_fd_sc_hd__a21oi_2 _49551_ (.A1(_19546_),
    .A2(_19631_),
    .B1(_19728_),
    .Y(_20664_));
 sky130_fd_sc_hd__a21bo_1 _49552_ (.A1(_19585_),
    .A2(_19621_),
    .B1_N(_19623_),
    .X(_20665_));
 sky130_fd_sc_hd__clkbuf_2 _49553_ (.A(\delay_line[33][7] ),
    .X(_20666_));
 sky130_fd_sc_hd__o21ai_1 _49554_ (.A1(net314),
    .A2(net313),
    .B1(_20666_),
    .Y(_20667_));
 sky130_fd_sc_hd__a21o_1 _49555_ (.A1(_19570_),
    .A2(_05337_),
    .B1(_20667_),
    .X(_20668_));
 sky130_fd_sc_hd__and2_1 _49556_ (.A(\delay_line[33][2] ),
    .B(net313),
    .X(_20669_));
 sky130_fd_sc_hd__nor2_2 _49557_ (.A(_02150_),
    .B(\delay_line[33][3] ),
    .Y(_20670_));
 sky130_fd_sc_hd__inv_2 _49558_ (.A(\delay_line[33][7] ),
    .Y(_20671_));
 sky130_fd_sc_hd__o21ai_1 _49559_ (.A1(_20669_),
    .A2(_20670_),
    .B1(_20671_),
    .Y(_20672_));
 sky130_fd_sc_hd__nand3b_2 _49560_ (.A_N(_19578_),
    .B(_20668_),
    .C(_20672_),
    .Y(_20673_));
 sky130_fd_sc_hd__o2bb2ai_1 _49561_ (.A1_N(_20668_),
    .A2_N(_20672_),
    .B1(_19572_),
    .B2(_19577_),
    .Y(_20674_));
 sky130_fd_sc_hd__or2b_1 _49562_ (.A(_02161_),
    .B_N(_00557_),
    .X(_20675_));
 sky130_fd_sc_hd__a21o_1 _49563_ (.A1(_20673_),
    .A2(_20674_),
    .B1(_20675_),
    .X(_20676_));
 sky130_fd_sc_hd__and2b_1 _49564_ (.A_N(_00557_),
    .B(\delay_line[33][0] ),
    .X(_20677_));
 sky130_fd_sc_hd__a21oi_1 _49565_ (.A1(_19580_),
    .A2(_20677_),
    .B1(_19579_),
    .Y(_20678_));
 sky130_fd_sc_hd__nand3_1 _49566_ (.A(_20675_),
    .B(_20673_),
    .C(_20674_),
    .Y(_20679_));
 sky130_fd_sc_hd__nand3_1 _49567_ (.A(_20676_),
    .B(_20678_),
    .C(_20679_),
    .Y(_20680_));
 sky130_fd_sc_hd__nand3_2 _49568_ (.A(_20680_),
    .B(_00579_),
    .C(_22523_),
    .Y(_20681_));
 sky130_fd_sc_hd__a21o_1 _49569_ (.A1(_20679_),
    .A2(_20676_),
    .B1(_20678_),
    .X(_20682_));
 sky130_fd_sc_hd__a22o_1 _49570_ (.A1(_22523_),
    .A2(_00590_),
    .B1(_20680_),
    .B2(_20682_),
    .X(_20683_));
 sky130_fd_sc_hd__nand3_4 _49571_ (.A(_19583_),
    .B(_20681_),
    .C(_20683_),
    .Y(_20684_));
 sky130_fd_sc_hd__a2bb2o_1 _49572_ (.A1_N(_19569_),
    .A2_N(_19582_),
    .B1(_20681_),
    .B2(_20683_),
    .X(_20685_));
 sky130_fd_sc_hd__buf_1 _49573_ (.A(\delay_line[32][7] ),
    .X(_20686_));
 sky130_fd_sc_hd__nand2_1 _49574_ (.A(_19589_),
    .B(_20686_),
    .Y(_20687_));
 sky130_fd_sc_hd__inv_2 _49575_ (.A(\delay_line[32][6] ),
    .Y(_20688_));
 sky130_fd_sc_hd__inv_2 _49576_ (.A(\delay_line[32][7] ),
    .Y(_20689_));
 sky130_fd_sc_hd__clkbuf_2 _49577_ (.A(_20689_),
    .X(_20690_));
 sky130_fd_sc_hd__nand2_1 _49578_ (.A(_20688_),
    .B(_20690_),
    .Y(_20691_));
 sky130_fd_sc_hd__a21oi_1 _49579_ (.A1(_20687_),
    .A2(_20691_),
    .B1(_18667_),
    .Y(_20692_));
 sky130_fd_sc_hd__clkbuf_2 _49580_ (.A(_20692_),
    .X(_20693_));
 sky130_fd_sc_hd__and2_2 _49581_ (.A(_19589_),
    .B(_20686_),
    .X(_20694_));
 sky130_fd_sc_hd__o21ai_1 _49582_ (.A1(_19589_),
    .A2(_20686_),
    .B1(_18663_),
    .Y(_20695_));
 sky130_fd_sc_hd__buf_2 _49583_ (.A(_20695_),
    .X(_20696_));
 sky130_fd_sc_hd__o21ai_4 _49584_ (.A1(_18671_),
    .A2(_19586_),
    .B1(_19590_),
    .Y(_20697_));
 sky130_fd_sc_hd__o21ai_4 _49585_ (.A1(_20694_),
    .A2(_20696_),
    .B1(_20697_),
    .Y(_20698_));
 sky130_fd_sc_hd__buf_1 _49586_ (.A(_19589_),
    .X(_20699_));
 sky130_fd_sc_hd__buf_1 _49587_ (.A(\delay_line[32][7] ),
    .X(_20700_));
 sky130_fd_sc_hd__a21oi_1 _49588_ (.A1(_20699_),
    .A2(_20700_),
    .B1(_20695_),
    .Y(_20701_));
 sky130_fd_sc_hd__o21bai_2 _49589_ (.A1(_20701_),
    .A2(_20692_),
    .B1_N(_20697_),
    .Y(_20702_));
 sky130_fd_sc_hd__o211a_1 _49590_ (.A1(_20693_),
    .A2(_20698_),
    .B1(_18660_),
    .C1(_20702_),
    .X(_20703_));
 sky130_fd_sc_hd__nor2_1 _49591_ (.A(_20699_),
    .B(_20700_),
    .Y(_20704_));
 sky130_fd_sc_hd__o21bai_2 _49592_ (.A1(_20694_),
    .A2(_20704_),
    .B1_N(_18667_),
    .Y(_20705_));
 sky130_fd_sc_hd__o211ai_2 _49593_ (.A1(_20696_),
    .A2(_20694_),
    .B1(_20697_),
    .C1(_20705_),
    .Y(_20706_));
 sky130_fd_sc_hd__a21oi_1 _49594_ (.A1(_20702_),
    .A2(_20706_),
    .B1(_18660_),
    .Y(_20707_));
 sky130_fd_sc_hd__o21ai_1 _49595_ (.A1(_05260_),
    .A2(_19593_),
    .B1(_19595_),
    .Y(_20708_));
 sky130_fd_sc_hd__o21bai_2 _49596_ (.A1(_20703_),
    .A2(_20707_),
    .B1_N(_20708_),
    .Y(_20709_));
 sky130_fd_sc_hd__o211ai_2 _49597_ (.A1(_20693_),
    .A2(_20698_),
    .B1(_18659_),
    .C1(_20702_),
    .Y(_20710_));
 sky130_fd_sc_hd__a21o_1 _49598_ (.A1(_20702_),
    .A2(_20706_),
    .B1(_18659_),
    .X(_20711_));
 sky130_fd_sc_hd__nand3_1 _49599_ (.A(_20710_),
    .B(_20711_),
    .C(_20708_),
    .Y(_20712_));
 sky130_fd_sc_hd__a21o_1 _49600_ (.A1(_20709_),
    .A2(_20712_),
    .B1(_24457_),
    .X(_20713_));
 sky130_fd_sc_hd__clkbuf_2 _49601_ (.A(_20712_),
    .X(_20714_));
 sky130_fd_sc_hd__nand3_2 _49602_ (.A(_20709_),
    .B(_20714_),
    .C(_24468_),
    .Y(_20715_));
 sky130_fd_sc_hd__nand2_2 _49603_ (.A(_19606_),
    .B(_19605_),
    .Y(_20716_));
 sky130_fd_sc_hd__nand3_2 _49604_ (.A(_20713_),
    .B(_20715_),
    .C(_20716_),
    .Y(_20717_));
 sky130_fd_sc_hd__a21oi_1 _49605_ (.A1(_20709_),
    .A2(_20714_),
    .B1(_24468_),
    .Y(_20718_));
 sky130_fd_sc_hd__and3_1 _49606_ (.A(_20709_),
    .B(_20714_),
    .C(_24468_),
    .X(_20719_));
 sky130_fd_sc_hd__and2_1 _49607_ (.A(_19606_),
    .B(_19605_),
    .X(_20720_));
 sky130_fd_sc_hd__o21ai_2 _49608_ (.A1(_20718_),
    .A2(_20719_),
    .B1(_20720_),
    .Y(_20721_));
 sky130_fd_sc_hd__nand2_1 _49609_ (.A(_19605_),
    .B(_19607_),
    .Y(_20722_));
 sky130_fd_sc_hd__o2bb2ai_1 _49610_ (.A1_N(_20717_),
    .A2_N(_20721_),
    .B1(_18681_),
    .B2(_20722_),
    .Y(_20723_));
 sky130_fd_sc_hd__nand4_2 _49611_ (.A(_20721_),
    .B(_19616_),
    .C(_19613_),
    .D(_20717_),
    .Y(_20724_));
 sky130_fd_sc_hd__a22oi_4 _49612_ (.A1(_19616_),
    .A2(_19610_),
    .B1(_20723_),
    .B2(_20724_),
    .Y(_20725_));
 sky130_fd_sc_hd__a2bb2oi_2 _49613_ (.A1_N(_18681_),
    .A2_N(_20722_),
    .B1(_20717_),
    .B2(_20721_),
    .Y(_20726_));
 sky130_fd_sc_hd__or4_1 _49614_ (.A(_19615_),
    .B(_18685_),
    .C(_19614_),
    .D(_18683_),
    .X(_20727_));
 sky130_fd_sc_hd__nor2_1 _49615_ (.A(_20726_),
    .B(_20727_),
    .Y(_20728_));
 sky130_fd_sc_hd__o211ai_4 _49616_ (.A1(_19608_),
    .A2(_19610_),
    .B1(_19612_),
    .C1(_19617_),
    .Y(_20729_));
 sky130_fd_sc_hd__o21ai_2 _49617_ (.A1(_20725_),
    .A2(_20728_),
    .B1(_20729_),
    .Y(_20730_));
 sky130_fd_sc_hd__or4_1 _49618_ (.A(_18686_),
    .B(_18683_),
    .C(_19619_),
    .D(_20725_),
    .X(_20731_));
 sky130_fd_sc_hd__a22oi_1 _49619_ (.A1(_20684_),
    .A2(_20685_),
    .B1(_20730_),
    .B2(_20731_),
    .Y(_20732_));
 sky130_fd_sc_hd__inv_2 _49620_ (.A(_20732_),
    .Y(_20733_));
 sky130_fd_sc_hd__nand2_1 _49621_ (.A(_19561_),
    .B(_18637_),
    .Y(_20734_));
 sky130_fd_sc_hd__nand3_1 _49622_ (.A(_19552_),
    .B(_19555_),
    .C(_19558_),
    .Y(_20735_));
 sky130_fd_sc_hd__nor2_1 _49623_ (.A(\delay_line[34][4] ),
    .B(_18631_),
    .Y(_20736_));
 sky130_fd_sc_hd__and2_1 _49624_ (.A(_19548_),
    .B(_18631_),
    .X(_20737_));
 sky130_fd_sc_hd__o21bai_1 _49625_ (.A1(_20736_),
    .A2(_20737_),
    .B1_N(_18630_),
    .Y(_20738_));
 sky130_fd_sc_hd__nand2_1 _49626_ (.A(_19548_),
    .B(_18631_),
    .Y(_20739_));
 sky130_fd_sc_hd__nand3b_2 _49627_ (.A_N(_20736_),
    .B(_20739_),
    .C(_05392_),
    .Y(_20740_));
 sky130_fd_sc_hd__clkbuf_2 _49628_ (.A(\delay_line[34][7] ),
    .X(_20741_));
 sky130_fd_sc_hd__nand3_1 _49629_ (.A(_17810_),
    .B(_19553_),
    .C(_20741_),
    .Y(_20742_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49630_ (.A(\delay_line[34][7] ),
    .X(_20743_));
 sky130_fd_sc_hd__a21o_1 _49631_ (.A1(_19548_),
    .A2(_19549_),
    .B1(_20743_),
    .X(_20744_));
 sky130_fd_sc_hd__nand2_1 _49632_ (.A(_20742_),
    .B(_20744_),
    .Y(_20745_));
 sky130_fd_sc_hd__a21oi_1 _49633_ (.A1(_20738_),
    .A2(_20740_),
    .B1(_20745_),
    .Y(_20746_));
 sky130_fd_sc_hd__and3_1 _49634_ (.A(_20738_),
    .B(_20740_),
    .C(_20745_),
    .X(_20747_));
 sky130_fd_sc_hd__a211o_1 _49635_ (.A1(_19555_),
    .A2(_20735_),
    .B1(_20746_),
    .C1(_20747_),
    .X(_20748_));
 sky130_fd_sc_hd__and3b_1 _49636_ (.A_N(\delay_line[34][0] ),
    .B(_02249_),
    .C(_05403_),
    .X(_20749_));
 sky130_fd_sc_hd__a21oi_1 _49637_ (.A1(\delay_line[34][0] ),
    .A2(_19557_),
    .B1(_20749_),
    .Y(_20750_));
 sky130_fd_sc_hd__o211ai_2 _49638_ (.A1(_20746_),
    .A2(_20747_),
    .B1(_19555_),
    .C1(_20735_),
    .Y(_20751_));
 sky130_fd_sc_hd__and3_1 _49639_ (.A(_20748_),
    .B(_20750_),
    .C(_20751_),
    .X(_20752_));
 sky130_fd_sc_hd__a21oi_1 _49640_ (.A1(_20751_),
    .A2(_20748_),
    .B1(_20750_),
    .Y(_20753_));
 sky130_fd_sc_hd__or2_1 _49641_ (.A(_20752_),
    .B(_20753_),
    .X(_20754_));
 sky130_fd_sc_hd__and3_1 _49642_ (.A(_19562_),
    .B(_20734_),
    .C(_20754_),
    .X(_20755_));
 sky130_fd_sc_hd__a21oi_1 _49643_ (.A1(_19562_),
    .A2(_20734_),
    .B1(_20754_),
    .Y(_20756_));
 sky130_fd_sc_hd__a21boi_2 _49644_ (.A1(_18648_),
    .A2(_19565_),
    .B1_N(_19566_),
    .Y(_20757_));
 sky130_fd_sc_hd__o21a_1 _49645_ (.A1(_20755_),
    .A2(_20756_),
    .B1(_20757_),
    .X(_20758_));
 sky130_fd_sc_hd__nor3_1 _49646_ (.A(_20755_),
    .B(_20756_),
    .C(_20757_),
    .Y(_20759_));
 sky130_fd_sc_hd__nor2_1 _49647_ (.A(_20758_),
    .B(_20759_),
    .Y(_20760_));
 sky130_fd_sc_hd__o2111ai_4 _49648_ (.A1(_20725_),
    .A2(_20729_),
    .B1(_20684_),
    .C1(_20730_),
    .D1(_20685_),
    .Y(_20761_));
 sky130_fd_sc_hd__nand3_1 _49649_ (.A(_20733_),
    .B(_20760_),
    .C(_20761_),
    .Y(_20762_));
 sky130_fd_sc_hd__a21o_1 _49650_ (.A1(_20761_),
    .A2(_20733_),
    .B1(_20760_),
    .X(_20763_));
 sky130_fd_sc_hd__a211oi_1 _49651_ (.A1(_20762_),
    .A2(_20763_),
    .B1(_19349_),
    .C1(net141),
    .Y(_20764_));
 sky130_fd_sc_hd__o211a_1 _49652_ (.A1(_19349_),
    .A2(net141),
    .B1(_20762_),
    .C1(_20763_),
    .X(_20765_));
 sky130_fd_sc_hd__nor2_1 _49653_ (.A(_20764_),
    .B(_20765_),
    .Y(_20766_));
 sky130_fd_sc_hd__xnor2_1 _49654_ (.A(_20665_),
    .B(_20766_),
    .Y(_20767_));
 sky130_fd_sc_hd__o211ai_1 _49655_ (.A1(_19628_),
    .A2(_19547_),
    .B1(_19627_),
    .C1(_20767_),
    .Y(_20768_));
 sky130_fd_sc_hd__a21o_1 _49656_ (.A1(_19627_),
    .A2(_19629_),
    .B1(_20767_),
    .X(_20769_));
 sky130_fd_sc_hd__and2_1 _49657_ (.A(_20768_),
    .B(_20769_),
    .X(_20770_));
 sky130_fd_sc_hd__buf_1 _49658_ (.A(_19636_),
    .X(_20771_));
 sky130_fd_sc_hd__a21oi_1 _49659_ (.A1(_19633_),
    .A2(_20771_),
    .B1(\delay_line[40][7] ),
    .Y(_20772_));
 sky130_fd_sc_hd__and3_1 _49660_ (.A(_19633_),
    .B(_20771_),
    .C(\delay_line[40][7] ),
    .X(_20773_));
 sky130_fd_sc_hd__nor3b_2 _49661_ (.A(_20772_),
    .B(_20773_),
    .C_N(_05689_),
    .Y(_20774_));
 sky130_fd_sc_hd__o21ba_1 _49662_ (.A1(_20772_),
    .A2(_20773_),
    .B1_N(_05689_),
    .X(_20775_));
 sky130_fd_sc_hd__o211ai_2 _49663_ (.A1(_20774_),
    .A2(_20775_),
    .B1(_19637_),
    .C1(_19640_),
    .Y(_20776_));
 sky130_fd_sc_hd__inv_2 _49664_ (.A(_20776_),
    .Y(_20777_));
 sky130_fd_sc_hd__a211oi_2 _49665_ (.A1(_19637_),
    .A2(_19640_),
    .B1(_20774_),
    .C1(_20775_),
    .Y(_20778_));
 sky130_fd_sc_hd__nand2_1 _49666_ (.A(_19642_),
    .B(_19635_),
    .Y(_20779_));
 sky130_fd_sc_hd__o21ai_1 _49667_ (.A1(_19644_),
    .A2(_19643_),
    .B1(_20779_),
    .Y(_20780_));
 sky130_fd_sc_hd__or3b_2 _49668_ (.A(_20777_),
    .B(_20778_),
    .C_N(_20780_),
    .X(_20781_));
 sky130_fd_sc_hd__o221ai_4 _49669_ (.A1(_20777_),
    .A2(_20778_),
    .B1(_19644_),
    .B2(_19643_),
    .C1(_20779_),
    .Y(_20782_));
 sky130_fd_sc_hd__and3_1 _49670_ (.A(_17780_),
    .B(_18599_),
    .C(_19647_),
    .X(_20783_));
 sky130_fd_sc_hd__nor2_1 _49671_ (.A(_19649_),
    .B(\delay_line[38][7] ),
    .Y(_20784_));
 sky130_fd_sc_hd__nand2_1 _49672_ (.A(\delay_line[38][4] ),
    .B(\delay_line[38][7] ),
    .Y(_20785_));
 sky130_fd_sc_hd__nor2b_1 _49673_ (.A(_20784_),
    .B_N(_20785_),
    .Y(_20786_));
 sky130_fd_sc_hd__buf_1 _49674_ (.A(\delay_line[38][6] ),
    .X(_20787_));
 sky130_fd_sc_hd__o211a_1 _49675_ (.A1(net289),
    .A2(\delay_line[38][6] ),
    .B1(\delay_line[38][5] ),
    .C1(net290),
    .X(_20788_));
 sky130_fd_sc_hd__a21oi_1 _49676_ (.A1(\delay_line[38][3] ),
    .A2(_20787_),
    .B1(_20788_),
    .Y(_20789_));
 sky130_fd_sc_hd__xor2_1 _49677_ (.A(_20786_),
    .B(_20789_),
    .X(_20790_));
 sky130_fd_sc_hd__o21ba_1 _49678_ (.A1(_19652_),
    .A2(_20783_),
    .B1_N(_20790_),
    .X(_20791_));
 sky130_fd_sc_hd__nand2_1 _49679_ (.A(_19647_),
    .B(_19646_),
    .Y(_20792_));
 sky130_fd_sc_hd__and3b_1 _49680_ (.A_N(_19652_),
    .B(_20790_),
    .C(_20792_),
    .X(_20793_));
 sky130_fd_sc_hd__nor2_1 _49681_ (.A(net283),
    .B(net282),
    .Y(_20794_));
 sky130_fd_sc_hd__nand2_1 _49682_ (.A(\delay_line[39][6] ),
    .B(net282),
    .Y(_20795_));
 sky130_fd_sc_hd__or3b_1 _49683_ (.A(_19660_),
    .B(_20794_),
    .C_N(_20795_),
    .X(_20796_));
 sky130_fd_sc_hd__inv_2 _49684_ (.A(net282),
    .Y(_20797_));
 sky130_fd_sc_hd__nand2_1 _49685_ (.A(_19661_),
    .B(_20797_),
    .Y(_20798_));
 sky130_fd_sc_hd__a21o_1 _49686_ (.A1(_20798_),
    .A2(_20795_),
    .B1(_18606_),
    .X(_20799_));
 sky130_fd_sc_hd__nand2_1 _49687_ (.A(_20796_),
    .B(_20799_),
    .Y(_20800_));
 sky130_fd_sc_hd__a21oi_2 _49688_ (.A1(_19658_),
    .A2(_19659_),
    .B1(_20800_),
    .Y(_20801_));
 sky130_fd_sc_hd__a311oi_2 _49689_ (.A1(_19657_),
    .A2(_19658_),
    .A3(_20800_),
    .B1(_19656_),
    .C1(_20801_),
    .Y(_20802_));
 sky130_fd_sc_hd__and3_1 _49690_ (.A(_19658_),
    .B(_19659_),
    .C(_20800_),
    .X(_20803_));
 sky130_fd_sc_hd__o21a_1 _49691_ (.A1(_20801_),
    .A2(_20803_),
    .B1(_19656_),
    .X(_20804_));
 sky130_fd_sc_hd__o211ai_1 _49692_ (.A1(_18609_),
    .A2(_19655_),
    .B1(_19659_),
    .C1(_19664_),
    .Y(_20805_));
 sky130_fd_sc_hd__o21a_1 _49693_ (.A1(_20802_),
    .A2(_20804_),
    .B1(_20805_),
    .X(_20806_));
 sky130_fd_sc_hd__buf_1 _49694_ (.A(_20802_),
    .X(_20807_));
 sky130_fd_sc_hd__a211oi_1 _49695_ (.A1(_20805_),
    .A2(_19667_),
    .B1(_20807_),
    .C1(_20804_),
    .Y(_20808_));
 sky130_fd_sc_hd__a21o_1 _49696_ (.A1(_19667_),
    .A2(_20806_),
    .B1(_20808_),
    .X(_20809_));
 sky130_fd_sc_hd__nor3b_1 _49697_ (.A(_19671_),
    .B(_19672_),
    .C_N(_20809_),
    .Y(_20810_));
 sky130_fd_sc_hd__o21ba_1 _49698_ (.A1(_19671_),
    .A2(_19672_),
    .B1_N(_20809_),
    .X(_20811_));
 sky130_fd_sc_hd__o22ai_2 _49699_ (.A1(_20791_),
    .A2(_20793_),
    .B1(_20810_),
    .B2(_20811_),
    .Y(_20812_));
 sky130_fd_sc_hd__or4_2 _49700_ (.A(_20791_),
    .B(_20793_),
    .C(_20810_),
    .D(_20811_),
    .X(_20813_));
 sky130_fd_sc_hd__and4_2 _49701_ (.A(_20781_),
    .B(_20782_),
    .C(_20812_),
    .D(_20813_),
    .X(_20814_));
 sky130_fd_sc_hd__a22oi_4 _49702_ (.A1(_20781_),
    .A2(_20782_),
    .B1(_20812_),
    .B2(_20813_),
    .Y(_20815_));
 sky130_fd_sc_hd__and3b_1 _49703_ (.A_N(_05986_),
    .B(_18570_),
    .C(_19681_),
    .X(_20816_));
 sky130_fd_sc_hd__nor2b_1 _49704_ (.A(_18570_),
    .B_N(net292),
    .Y(_20817_));
 sky130_fd_sc_hd__and2b_1 _49705_ (.A_N(\delay_line[37][7] ),
    .B(_18570_),
    .X(_20818_));
 sky130_fd_sc_hd__nor2_1 _49706_ (.A(_20817_),
    .B(_20818_),
    .Y(_20819_));
 sky130_fd_sc_hd__o21ai_1 _49707_ (.A1(_19678_),
    .A2(_20816_),
    .B1(_20819_),
    .Y(_20820_));
 sky130_fd_sc_hd__or3_1 _49708_ (.A(_19678_),
    .B(_20819_),
    .C(_20816_),
    .X(_20821_));
 sky130_fd_sc_hd__a31o_1 _49709_ (.A1(_19679_),
    .A2(_17521_),
    .A3(_18572_),
    .B1(_19686_),
    .X(_20822_));
 sky130_fd_sc_hd__and3_1 _49710_ (.A(_20820_),
    .B(_20821_),
    .C(_20822_),
    .X(_20823_));
 sky130_fd_sc_hd__a21oi_1 _49711_ (.A1(_20820_),
    .A2(_20821_),
    .B1(_20822_),
    .Y(_20824_));
 sky130_fd_sc_hd__and2b_1 _49712_ (.A_N(\delay_line[36][2] ),
    .B(\delay_line[36][4] ),
    .X(_20825_));
 sky130_fd_sc_hd__and2b_1 _49713_ (.A_N(\delay_line[36][4] ),
    .B(\delay_line[36][2] ),
    .X(_20826_));
 sky130_fd_sc_hd__nor2_1 _49714_ (.A(_20825_),
    .B(_20826_),
    .Y(_20827_));
 sky130_fd_sc_hd__or2b_1 _49715_ (.A(\delay_line[36][1] ),
    .B_N(\delay_line[36][3] ),
    .X(_20828_));
 sky130_fd_sc_hd__a21boi_1 _49716_ (.A1(_18545_),
    .A2(_19716_),
    .B1_N(_20828_),
    .Y(_20829_));
 sky130_fd_sc_hd__xor2_1 _49717_ (.A(_20827_),
    .B(_20829_),
    .X(_20830_));
 sky130_fd_sc_hd__o31a_1 _49718_ (.A1(_05931_),
    .A2(_18546_),
    .A3(_19718_),
    .B1(_20830_),
    .X(_20831_));
 sky130_fd_sc_hd__nor4_1 _49719_ (.A(\delay_line[36][0] ),
    .B(_18545_),
    .C(_19718_),
    .D(_20830_),
    .Y(_20832_));
 sky130_fd_sc_hd__clkbuf_2 _49720_ (.A(_18550_),
    .X(_20833_));
 sky130_fd_sc_hd__buf_1 _49721_ (.A(\delay_line[35][7] ),
    .X(_20834_));
 sky130_fd_sc_hd__buf_1 _49722_ (.A(_19690_),
    .X(_20835_));
 sky130_fd_sc_hd__and2b_1 _49723_ (.A_N(_20834_),
    .B(_20835_),
    .X(_20836_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49724_ (.A(_20835_),
    .X(_20837_));
 sky130_fd_sc_hd__buf_1 _49725_ (.A(_20834_),
    .X(_20838_));
 sky130_fd_sc_hd__o21ai_1 _49726_ (.A1(_20837_),
    .A2(_20838_),
    .B1(_20833_),
    .Y(_20839_));
 sky130_fd_sc_hd__and2_1 _49727_ (.A(_20835_),
    .B(_20834_),
    .X(_20840_));
 sky130_fd_sc_hd__o22a_1 _49728_ (.A1(_20833_),
    .A2(_20836_),
    .B1(_20839_),
    .B2(_20840_),
    .X(_20841_));
 sky130_fd_sc_hd__clkbuf_2 _49729_ (.A(_20838_),
    .X(_20842_));
 sky130_fd_sc_hd__nor2_1 _49730_ (.A(_20842_),
    .B(_19691_),
    .Y(_20843_));
 sky130_fd_sc_hd__o211a_1 _49731_ (.A1(_20841_),
    .A2(_20843_),
    .B1(_19696_),
    .C1(_19704_),
    .X(_20844_));
 sky130_fd_sc_hd__a211oi_2 _49732_ (.A1(_19696_),
    .A2(_19704_),
    .B1(_20841_),
    .C1(_20843_),
    .Y(_20845_));
 sky130_fd_sc_hd__o21a_1 _49733_ (.A1(_20844_),
    .A2(_20845_),
    .B1(_05832_),
    .X(_20846_));
 sky130_fd_sc_hd__nor3_2 _49734_ (.A(_05832_),
    .B(_20844_),
    .C(_20845_),
    .Y(_20847_));
 sky130_fd_sc_hd__a211oi_1 _49735_ (.A1(_19705_),
    .A2(_19707_),
    .B1(_20846_),
    .C1(_20847_),
    .Y(_20848_));
 sky130_fd_sc_hd__o221a_1 _49736_ (.A1(_22677_),
    .A2(_19701_),
    .B1(_20846_),
    .B2(_20847_),
    .C1(_19705_),
    .X(_20849_));
 sky130_fd_sc_hd__nor2_1 _49737_ (.A(_20848_),
    .B(_20849_),
    .Y(_20850_));
 sky130_fd_sc_hd__o211ai_2 _49738_ (.A1(_19710_),
    .A2(_18565_),
    .B1(_19708_),
    .C1(_19711_),
    .Y(_20851_));
 sky130_fd_sc_hd__xor2_1 _49739_ (.A(_20850_),
    .B(_20851_),
    .X(_20852_));
 sky130_fd_sc_hd__o21bai_1 _49740_ (.A1(_20831_),
    .A2(_20832_),
    .B1_N(_20852_),
    .Y(_20853_));
 sky130_fd_sc_hd__or3b_1 _49741_ (.A(_20831_),
    .B(_20832_),
    .C_N(_20852_),
    .X(_20854_));
 sky130_fd_sc_hd__or4bb_2 _49742_ (.A(_20823_),
    .B(_20824_),
    .C_N(_20853_),
    .D_N(_20854_),
    .X(_20855_));
 sky130_fd_sc_hd__a2bb2o_1 _49743_ (.A1_N(_20823_),
    .A2_N(_20824_),
    .B1(_20853_),
    .B2(_20854_),
    .X(_20856_));
 sky130_fd_sc_hd__a221oi_2 _49744_ (.A1(_19687_),
    .A2(_19722_),
    .B1(_20855_),
    .B2(_20856_),
    .C1(_19720_),
    .Y(_20857_));
 sky130_fd_sc_hd__and3b_1 _49745_ (.A_N(_19720_),
    .B(_19721_),
    .C(_19687_),
    .X(_20858_));
 sky130_fd_sc_hd__o211a_1 _49746_ (.A1(_19720_),
    .A2(_20858_),
    .B1(_20855_),
    .C1(_20856_),
    .X(_20859_));
 sky130_fd_sc_hd__nor4_1 _49747_ (.A(_20814_),
    .B(_20815_),
    .C(_20857_),
    .D(_20859_),
    .Y(_20860_));
 sky130_fd_sc_hd__o22a_1 _49748_ (.A1(_20814_),
    .A2(_20815_),
    .B1(_20857_),
    .B2(_20859_),
    .X(_20861_));
 sky130_fd_sc_hd__nor2_2 _49749_ (.A(net104),
    .B(_20861_),
    .Y(_20862_));
 sky130_fd_sc_hd__xor2_1 _49750_ (.A(_20770_),
    .B(_20862_),
    .X(_20863_));
 sky130_fd_sc_hd__and2_1 _49751_ (.A(_19384_),
    .B(_19387_),
    .X(_20864_));
 sky130_fd_sc_hd__or2b_1 _49752_ (.A(_20863_),
    .B_N(_20864_),
    .X(_20865_));
 sky130_fd_sc_hd__a21bo_1 _49753_ (.A1(_19384_),
    .A2(_19387_),
    .B1_N(_20863_),
    .X(_20866_));
 sky130_fd_sc_hd__nand2_1 _49754_ (.A(_20865_),
    .B(_20866_),
    .Y(_20867_));
 sky130_fd_sc_hd__xnor2_1 _49755_ (.A(_20664_),
    .B(_20867_),
    .Y(_20868_));
 sky130_fd_sc_hd__xnor2_2 _49756_ (.A(_20663_),
    .B(_20868_),
    .Y(_20869_));
 sky130_fd_sc_hd__xor2_2 _49757_ (.A(_20300_),
    .B(_20869_),
    .X(_20870_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49758_ (.A(_20289_),
    .X(_20871_));
 sky130_fd_sc_hd__o22ai_1 _49759_ (.A1(_19847_),
    .A2(_19850_),
    .B1(_20288_),
    .B2(_20871_),
    .Y(_20872_));
 sky130_fd_sc_hd__nand3b_1 _49760_ (.A_N(_20293_),
    .B(_20284_),
    .C(_20286_),
    .Y(_20873_));
 sky130_fd_sc_hd__nand3b_2 _49761_ (.A_N(_20295_),
    .B(_20872_),
    .C(_20873_),
    .Y(_20874_));
 sky130_fd_sc_hd__o32a_1 _49762_ (.A1(_19231_),
    .A2(_19229_),
    .A3(_19247_),
    .B1(_19240_),
    .B2(_19239_),
    .X(_20875_));
 sky130_fd_sc_hd__o2bb2ai_2 _49763_ (.A1_N(_20874_),
    .A2_N(_20297_),
    .B1(_20875_),
    .B2(_19235_),
    .Y(_20876_));
 sky130_fd_sc_hd__o211ai_2 _49764_ (.A1(_20296_),
    .A2(_20299_),
    .B1(_20870_),
    .C1(_20876_),
    .Y(_20877_));
 sky130_fd_sc_hd__o2111ai_4 _49765_ (.A1(_19242_),
    .A2(net60),
    .B1(_19248_),
    .C1(_20874_),
    .D1(_20297_),
    .Y(_20878_));
 sky130_fd_sc_hd__a21o_1 _49766_ (.A1(_20878_),
    .A2(_20876_),
    .B1(_20870_),
    .X(_20879_));
 sky130_fd_sc_hd__nand3_2 _49767_ (.A(_19844_),
    .B(_20877_),
    .C(_20879_),
    .Y(_20880_));
 sky130_fd_sc_hd__o211a_1 _49768_ (.A1(_20296_),
    .A2(_20299_),
    .B1(_20870_),
    .C1(_20876_),
    .X(_20881_));
 sky130_fd_sc_hd__a21oi_1 _49769_ (.A1(_20878_),
    .A2(_20876_),
    .B1(_20870_),
    .Y(_20882_));
 sky130_fd_sc_hd__o31a_1 _49770_ (.A1(_19739_),
    .A2(_19256_),
    .A3(_19259_),
    .B1(_19843_),
    .X(_20883_));
 sky130_fd_sc_hd__o21ai_2 _49771_ (.A1(_20881_),
    .A2(_20882_),
    .B1(_20883_),
    .Y(_20884_));
 sky130_fd_sc_hd__o211ai_1 _49772_ (.A1(_19841_),
    .A2(_19842_),
    .B1(_20880_),
    .C1(_20884_),
    .Y(_20885_));
 sky130_fd_sc_hd__nand2_1 _49773_ (.A(_20880_),
    .B(_20884_),
    .Y(_20886_));
 sky130_fd_sc_hd__nor2_1 _49774_ (.A(_19841_),
    .B(_19842_),
    .Y(_20887_));
 sky130_fd_sc_hd__nand2_1 _49775_ (.A(_20886_),
    .B(_20887_),
    .Y(_20888_));
 sky130_fd_sc_hd__nand3b_2 _49776_ (.A_N(_19788_),
    .B(_20885_),
    .C(_20888_),
    .Y(_20889_));
 sky130_fd_sc_hd__o21ai_1 _49777_ (.A1(_19841_),
    .A2(_19842_),
    .B1(_20886_),
    .Y(_20890_));
 sky130_fd_sc_hd__nand3_1 _49778_ (.A(_20887_),
    .B(_20880_),
    .C(_20884_),
    .Y(_20891_));
 sky130_fd_sc_hd__nand3_2 _49779_ (.A(_19788_),
    .B(_20890_),
    .C(_20891_),
    .Y(_20892_));
 sky130_fd_sc_hd__and3_1 _49780_ (.A(_05161_),
    .B(_18765_),
    .C(_19762_),
    .X(_20893_));
 sky130_fd_sc_hd__a21oi_2 _49781_ (.A1(_18752_),
    .A2(_18831_),
    .B1(_18830_),
    .Y(_20894_));
 sky130_fd_sc_hd__nand2_2 _49782_ (.A(_18782_),
    .B(_19761_),
    .Y(_20895_));
 sky130_fd_sc_hd__clkbuf_2 _49783_ (.A(_19825_),
    .X(_20896_));
 sky130_fd_sc_hd__nor2_1 _49784_ (.A(_20896_),
    .B(_18824_),
    .Y(_20897_));
 sky130_fd_sc_hd__clkbuf_2 _49785_ (.A(_10778_),
    .X(_20898_));
 sky130_fd_sc_hd__o32a_1 _49786_ (.A1(_20896_),
    .A2(_10833_),
    .A3(_19757_),
    .B1(_20897_),
    .B2(_20898_),
    .X(_20899_));
 sky130_fd_sc_hd__a311oi_2 _49787_ (.A1(_18733_),
    .A2(_18819_),
    .A3(_18820_),
    .B1(_18826_),
    .C1(_20899_),
    .Y(_20900_));
 sky130_fd_sc_hd__o21a_2 _49788_ (.A1(_18821_),
    .A2(_18826_),
    .B1(_20899_),
    .X(_20901_));
 sky130_fd_sc_hd__a311oi_2 _49789_ (.A1(_19757_),
    .A2(_18780_),
    .A3(_05172_),
    .B1(_20900_),
    .C1(_20901_),
    .Y(_20902_));
 sky130_fd_sc_hd__o2111a_1 _49790_ (.A1(_20900_),
    .A2(_20901_),
    .B1(_19757_),
    .C1(_18780_),
    .D1(_05172_),
    .X(_20903_));
 sky130_fd_sc_hd__nor2_1 _49791_ (.A(_20902_),
    .B(_20903_),
    .Y(_20904_));
 sky130_fd_sc_hd__xor2_2 _49792_ (.A(_20895_),
    .B(_20904_),
    .X(_20905_));
 sky130_fd_sc_hd__xnor2_2 _49793_ (.A(_20894_),
    .B(_20905_),
    .Y(_20906_));
 sky130_fd_sc_hd__xnor2_2 _49794_ (.A(_20893_),
    .B(_20906_),
    .Y(_20907_));
 sky130_fd_sc_hd__inv_2 _49795_ (.A(_20907_),
    .Y(_20908_));
 sky130_fd_sc_hd__nand3_1 _49796_ (.A(_20889_),
    .B(_20892_),
    .C(_20908_),
    .Y(_20909_));
 sky130_fd_sc_hd__nand2_1 _49797_ (.A(_20889_),
    .B(_20892_),
    .Y(_20910_));
 sky130_fd_sc_hd__nand2_1 _49798_ (.A(_20910_),
    .B(_20907_),
    .Y(_20911_));
 sky130_fd_sc_hd__nand3b_2 _49799_ (.A_N(_19787_),
    .B(_20909_),
    .C(_20911_),
    .Y(_20912_));
 sky130_fd_sc_hd__nand2_1 _49800_ (.A(_20910_),
    .B(_20908_),
    .Y(_20913_));
 sky130_fd_sc_hd__nand3_1 _49801_ (.A(_20889_),
    .B(_20892_),
    .C(_20907_),
    .Y(_20914_));
 sky130_fd_sc_hd__nand3_1 _49802_ (.A(_19787_),
    .B(_20913_),
    .C(_20914_),
    .Y(_20915_));
 sky130_fd_sc_hd__and3_1 _49803_ (.A(_20912_),
    .B(_19764_),
    .C(_20915_),
    .X(_20916_));
 sky130_fd_sc_hd__nand2_1 _49804_ (.A(_19779_),
    .B(_19782_),
    .Y(_20917_));
 sky130_fd_sc_hd__a21oi_1 _49805_ (.A1(_18767_),
    .A2(_18757_),
    .B1(_18760_),
    .Y(_20918_));
 sky130_fd_sc_hd__o2bb2ai_1 _49806_ (.A1_N(_20915_),
    .A2_N(_20912_),
    .B1(_19763_),
    .B2(_20918_),
    .Y(_20919_));
 sky130_fd_sc_hd__nand2_1 _49807_ (.A(_20917_),
    .B(_20919_),
    .Y(_20920_));
 sky130_fd_sc_hd__nand3_1 _49808_ (.A(_20912_),
    .B(_19764_),
    .C(_20915_),
    .Y(_20921_));
 sky130_fd_sc_hd__a21oi_2 _49809_ (.A1(_20921_),
    .A2(_20919_),
    .B1(_20917_),
    .Y(_20922_));
 sky130_fd_sc_hd__o21bai_1 _49810_ (.A1(_20916_),
    .A2(_20920_),
    .B1_N(_20922_),
    .Y(_20923_));
 sky130_fd_sc_hd__xor2_1 _49811_ (.A(_19786_),
    .B(_20923_),
    .X(_00038_));
 sky130_fd_sc_hd__o22ai_4 _49812_ (.A1(_20916_),
    .A2(_20920_),
    .B1(_20922_),
    .B2(_19786_),
    .Y(_20924_));
 sky130_fd_sc_hd__a21bo_1 _49813_ (.A1(_20887_),
    .A2(_20884_),
    .B1_N(_20880_),
    .X(_20925_));
 sky130_fd_sc_hd__o31a_1 _49814_ (.A1(_19789_),
    .A2(_19803_),
    .A3(_19804_),
    .B1(_18807_),
    .X(_20926_));
 sky130_fd_sc_hd__a21oi_1 _49815_ (.A1(_19789_),
    .A2(_19805_),
    .B1(_20926_),
    .Y(_20927_));
 sky130_fd_sc_hd__xnor2_2 _49816_ (.A(_11416_),
    .B(_18800_),
    .Y(_20928_));
 sky130_fd_sc_hd__and2_1 _49817_ (.A(\delay_line[20][7] ),
    .B(\delay_line[20][8] ),
    .X(_20929_));
 sky130_fd_sc_hd__buf_1 _49818_ (.A(\delay_line[20][8] ),
    .X(_20930_));
 sky130_fd_sc_hd__nor2_1 _49819_ (.A(\delay_line[20][7] ),
    .B(_20930_),
    .Y(_20931_));
 sky130_fd_sc_hd__or3b_1 _49820_ (.A(_20929_),
    .B(_20931_),
    .C_N(_19791_),
    .X(_20932_));
 sky130_fd_sc_hd__a2bb2o_1 _49821_ (.A1_N(_20929_),
    .A2_N(_20931_),
    .B1(_19790_),
    .B2(_19792_),
    .X(_20933_));
 sky130_fd_sc_hd__and3b_1 _49822_ (.A_N(_20928_),
    .B(_20932_),
    .C(_20933_),
    .X(_20934_));
 sky130_fd_sc_hd__a21boi_1 _49823_ (.A1(_20933_),
    .A2(_20932_),
    .B1_N(_20928_),
    .Y(_20935_));
 sky130_fd_sc_hd__o22a_1 _49824_ (.A1(_19795_),
    .A2(_19796_),
    .B1(_19794_),
    .B2(_19799_),
    .X(_20936_));
 sky130_fd_sc_hd__o21a_1 _49825_ (.A1(_20934_),
    .A2(_20935_),
    .B1(_20936_),
    .X(_20937_));
 sky130_fd_sc_hd__or3_1 _49826_ (.A(_20934_),
    .B(_20935_),
    .C(_20936_),
    .X(_20938_));
 sky130_fd_sc_hd__and3b_1 _49827_ (.A_N(_20937_),
    .B(_19847_),
    .C(_20938_),
    .X(_20939_));
 sky130_fd_sc_hd__inv_2 _49828_ (.A(_20938_),
    .Y(_20940_));
 sky130_fd_sc_hd__o21a_1 _49829_ (.A1(_20940_),
    .A2(_20937_),
    .B1(_20290_),
    .X(_20941_));
 sky130_fd_sc_hd__or3b_1 _49830_ (.A(_20939_),
    .B(_20941_),
    .C_N(_19803_),
    .X(_20942_));
 sky130_fd_sc_hd__o21bai_1 _49831_ (.A1(_20939_),
    .A2(_20941_),
    .B1_N(_19803_),
    .Y(_20943_));
 sky130_fd_sc_hd__and2_1 _49832_ (.A(_20942_),
    .B(_20943_),
    .X(_20944_));
 sky130_fd_sc_hd__xnor2_1 _49833_ (.A(_20927_),
    .B(_20944_),
    .Y(_20945_));
 sky130_fd_sc_hd__clkbuf_2 _49834_ (.A(_11020_),
    .X(_20946_));
 sky130_fd_sc_hd__a21oi_2 _49835_ (.A1(_11042_),
    .A2(_19798_),
    .B1(_18737_),
    .Y(_20947_));
 sky130_fd_sc_hd__nor2_1 _49836_ (.A(_20947_),
    .B(_18743_),
    .Y(_20948_));
 sky130_fd_sc_hd__and2_1 _49837_ (.A(_18743_),
    .B(_20947_),
    .X(_20949_));
 sky130_fd_sc_hd__nor3_2 _49838_ (.A(_10943_),
    .B(_20948_),
    .C(_20949_),
    .Y(_20950_));
 sky130_fd_sc_hd__o21a_1 _49839_ (.A1(_20948_),
    .A2(_20949_),
    .B1(_10954_),
    .X(_20951_));
 sky130_fd_sc_hd__or2_2 _49840_ (.A(_19814_),
    .B(_10756_),
    .X(_20952_));
 sky130_fd_sc_hd__o221ai_4 _49841_ (.A1(_19819_),
    .A2(_19817_),
    .B1(_20950_),
    .B2(_20951_),
    .C1(_20952_),
    .Y(_20953_));
 sky130_fd_sc_hd__a21o_1 _49842_ (.A1(_10756_),
    .A2(_19815_),
    .B1(_10998_),
    .X(_20954_));
 sky130_fd_sc_hd__a211oi_4 _49843_ (.A1(_20952_),
    .A2(_20954_),
    .B1(net208),
    .C1(_20951_),
    .Y(_20955_));
 sky130_fd_sc_hd__inv_2 _49844_ (.A(_20955_),
    .Y(_20956_));
 sky130_fd_sc_hd__or2_1 _49845_ (.A(\delay_line[17][7] ),
    .B(net377),
    .X(_20957_));
 sky130_fd_sc_hd__nand2_2 _49846_ (.A(\delay_line[17][7] ),
    .B(net377),
    .Y(_20958_));
 sky130_fd_sc_hd__and2_1 _49847_ (.A(_20957_),
    .B(_20958_),
    .X(_20959_));
 sky130_fd_sc_hd__xor2_1 _49848_ (.A(_22172_),
    .B(_20959_),
    .X(_20960_));
 sky130_fd_sc_hd__a21o_1 _49849_ (.A1(_20953_),
    .A2(_20956_),
    .B1(_20960_),
    .X(_20961_));
 sky130_fd_sc_hd__nand3_1 _49850_ (.A(_20956_),
    .B(_20960_),
    .C(_20953_),
    .Y(_20962_));
 sky130_fd_sc_hd__a221o_1 _49851_ (.A1(_20946_),
    .A2(net181),
    .B1(_20961_),
    .B2(_20962_),
    .C1(_19821_),
    .X(_20963_));
 sky130_fd_sc_hd__buf_1 _49852_ (.A(_19809_),
    .X(_20964_));
 sky130_fd_sc_hd__buf_1 _49853_ (.A(_20964_),
    .X(_20965_));
 sky130_fd_sc_hd__nand2_1 _49854_ (.A(_20896_),
    .B(_19827_),
    .Y(_20966_));
 sky130_fd_sc_hd__buf_2 _49855_ (.A(_19827_),
    .X(_20967_));
 sky130_fd_sc_hd__or2b_1 _49856_ (.A(_19825_),
    .B_N(_20964_),
    .X(_20968_));
 sky130_fd_sc_hd__o211a_1 _49857_ (.A1(_20965_),
    .A2(_20966_),
    .B1(_20967_),
    .C1(_20968_),
    .X(_20969_));
 sky130_fd_sc_hd__a21o_1 _49858_ (.A1(_20946_),
    .A2(net181),
    .B1(_19821_),
    .X(_20970_));
 sky130_fd_sc_hd__nand3_2 _49859_ (.A(_20970_),
    .B(_20961_),
    .C(_20962_),
    .Y(_20971_));
 sky130_fd_sc_hd__nand3_1 _49860_ (.A(_20963_),
    .B(_20969_),
    .C(_20971_),
    .Y(_20972_));
 sky130_fd_sc_hd__a21o_1 _49861_ (.A1(_20971_),
    .A2(_20963_),
    .B1(_20969_),
    .X(_20973_));
 sky130_fd_sc_hd__and2_1 _49862_ (.A(_20972_),
    .B(_20973_),
    .X(_20974_));
 sky130_fd_sc_hd__xnor2_1 _49863_ (.A(_20945_),
    .B(_20974_),
    .Y(_20975_));
 sky130_fd_sc_hd__a21bo_1 _49864_ (.A1(_20874_),
    .A2(_20299_),
    .B1_N(_20975_),
    .X(_20976_));
 sky130_fd_sc_hd__a211o_1 _49865_ (.A1(_20297_),
    .A2(_20298_),
    .B1(_20975_),
    .C1(_20296_),
    .X(_20977_));
 sky130_fd_sc_hd__nor2_1 _49866_ (.A(_18749_),
    .B(_18808_),
    .Y(_20978_));
 sky130_fd_sc_hd__a32o_1 _49867_ (.A1(_19808_),
    .A2(_19830_),
    .A3(_19831_),
    .B1(_20978_),
    .B2(_19806_),
    .X(_20979_));
 sky130_fd_sc_hd__a21oi_1 _49868_ (.A1(_20976_),
    .A2(_20977_),
    .B1(_20979_),
    .Y(_20980_));
 sky130_fd_sc_hd__and3_1 _49869_ (.A(_20976_),
    .B(_20977_),
    .C(_20979_),
    .X(_20981_));
 sky130_fd_sc_hd__or2_1 _49870_ (.A(_20662_),
    .B(_20661_),
    .X(_20982_));
 sky130_fd_sc_hd__or2_1 _49871_ (.A(_20663_),
    .B(_20868_),
    .X(_20983_));
 sky130_fd_sc_hd__a21bo_1 _49872_ (.A1(_20768_),
    .A2(_20862_),
    .B1_N(_20769_),
    .X(_20984_));
 sky130_fd_sc_hd__nor2_1 _49873_ (.A(net282),
    .B(net281),
    .Y(_20985_));
 sky130_fd_sc_hd__buf_1 _49874_ (.A(_20797_),
    .X(_20986_));
 sky130_fd_sc_hd__inv_2 _49875_ (.A(\delay_line[39][8] ),
    .Y(_20987_));
 sky130_fd_sc_hd__nor2_1 _49876_ (.A(_20986_),
    .B(_20987_),
    .Y(_20988_));
 sky130_fd_sc_hd__or3_1 _49877_ (.A(_19662_),
    .B(_20985_),
    .C(_20988_),
    .X(_20989_));
 sky130_fd_sc_hd__o21ai_1 _49878_ (.A1(_20985_),
    .A2(_20988_),
    .B1(_19662_),
    .Y(_20990_));
 sky130_fd_sc_hd__nand2_1 _49879_ (.A(_20989_),
    .B(_20990_),
    .Y(_20991_));
 sky130_fd_sc_hd__a21oi_2 _49880_ (.A1(_20795_),
    .A2(_20796_),
    .B1(_20991_),
    .Y(_20992_));
 sky130_fd_sc_hd__a311oi_2 _49881_ (.A1(_20794_),
    .A2(_20795_),
    .A3(_20991_),
    .B1(_19660_),
    .C1(_20992_),
    .Y(_20993_));
 sky130_fd_sc_hd__and3_1 _49882_ (.A(_20795_),
    .B(_20796_),
    .C(_20991_),
    .X(_20994_));
 sky130_fd_sc_hd__o21a_1 _49883_ (.A1(_20992_),
    .A2(_20994_),
    .B1(_19660_),
    .X(_20995_));
 sky130_fd_sc_hd__or2_1 _49884_ (.A(_20993_),
    .B(_20995_),
    .X(_20996_));
 sky130_fd_sc_hd__or2b_1 _49885_ (.A(_20801_),
    .B_N(_20996_),
    .X(_20997_));
 sky130_fd_sc_hd__o21bai_1 _49886_ (.A1(_20801_),
    .A2(_20807_),
    .B1_N(_20996_),
    .Y(_20998_));
 sky130_fd_sc_hd__o221a_1 _49887_ (.A1(_20997_),
    .A2(_20807_),
    .B1(_20808_),
    .B2(_20811_),
    .C1(_20998_),
    .X(_20999_));
 sky130_fd_sc_hd__o21a_1 _49888_ (.A1(_20807_),
    .A2(_20997_),
    .B1(_20998_),
    .X(_21000_));
 sky130_fd_sc_hd__or3_1 _49889_ (.A(_20808_),
    .B(_20811_),
    .C(_21000_),
    .X(_21001_));
 sky130_fd_sc_hd__inv_2 _49890_ (.A(_21001_),
    .Y(_21002_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49891_ (.A(\delay_line[38][5] ),
    .X(_21003_));
 sky130_fd_sc_hd__nor2_1 _49892_ (.A(_21003_),
    .B(net287),
    .Y(_21004_));
 sky130_fd_sc_hd__and2_1 _49893_ (.A(_21003_),
    .B(net287),
    .X(_21005_));
 sky130_fd_sc_hd__nor2_1 _49894_ (.A(_21004_),
    .B(_21005_),
    .Y(_21006_));
 sky130_fd_sc_hd__o211ai_1 _49895_ (.A1(_19649_),
    .A2(\delay_line[38][7] ),
    .B1(_20787_),
    .C1(_05568_),
    .Y(_21007_));
 sky130_fd_sc_hd__and3_1 _49896_ (.A(_21006_),
    .B(_21007_),
    .C(_20785_),
    .X(_21008_));
 sky130_fd_sc_hd__a21oi_1 _49897_ (.A1(_20785_),
    .A2(_21007_),
    .B1(_21006_),
    .Y(_21009_));
 sky130_fd_sc_hd__a31o_1 _49898_ (.A1(_18596_),
    .A2(_19647_),
    .A3(_20786_),
    .B1(_20791_),
    .X(_21010_));
 sky130_fd_sc_hd__nor3_1 _49899_ (.A(_21008_),
    .B(_21009_),
    .C(_21010_),
    .Y(_21011_));
 sky130_fd_sc_hd__o21ai_1 _49900_ (.A1(_21008_),
    .A2(_21009_),
    .B1(_21010_),
    .Y(_21012_));
 sky130_fd_sc_hd__or2b_1 _49901_ (.A(_21011_),
    .B_N(_21012_),
    .X(_21013_));
 sky130_fd_sc_hd__o21a_1 _49902_ (.A1(_20999_),
    .A2(_21002_),
    .B1(_21013_),
    .X(_21014_));
 sky130_fd_sc_hd__inv_2 _49903_ (.A(_21014_),
    .Y(_21015_));
 sky130_fd_sc_hd__inv_2 _49904_ (.A(\delay_line[40][7] ),
    .Y(_21016_));
 sky130_fd_sc_hd__clkbuf_2 _49905_ (.A(_21016_),
    .X(_21017_));
 sky130_fd_sc_hd__a31o_1 _49906_ (.A1(\delay_line[40][5] ),
    .A2(_20771_),
    .A3(_21017_),
    .B1(_20774_),
    .X(_21018_));
 sky130_fd_sc_hd__buf_1 _49907_ (.A(\delay_line[40][8] ),
    .X(_21019_));
 sky130_fd_sc_hd__or3b_1 _49908_ (.A(\delay_line[40][8] ),
    .B(_21016_),
    .C_N(_19636_),
    .X(_21020_));
 sky130_fd_sc_hd__or3b_1 _49909_ (.A(_19636_),
    .B(_21016_),
    .C_N(_21019_),
    .X(_21021_));
 sky130_fd_sc_hd__o211a_1 _49910_ (.A1(\delay_line[40][7] ),
    .A2(_21019_),
    .B1(_21020_),
    .C1(_21021_),
    .X(_21022_));
 sky130_fd_sc_hd__nand2_1 _49911_ (.A(_17769_),
    .B(_21022_),
    .Y(_21023_));
 sky130_fd_sc_hd__or2_1 _49912_ (.A(_17769_),
    .B(_21022_),
    .X(_21024_));
 sky130_fd_sc_hd__and3_1 _49913_ (.A(_21018_),
    .B(_21023_),
    .C(_21024_),
    .X(_21025_));
 sky130_fd_sc_hd__a21oi_1 _49914_ (.A1(_21023_),
    .A2(_21024_),
    .B1(_21018_),
    .Y(_21026_));
 sky130_fd_sc_hd__a21oi_1 _49915_ (.A1(_20776_),
    .A2(_20780_),
    .B1(_20778_),
    .Y(_21027_));
 sky130_fd_sc_hd__or3_1 _49916_ (.A(_21025_),
    .B(_21026_),
    .C(_21027_),
    .X(_21028_));
 sky130_fd_sc_hd__o21ai_1 _49917_ (.A1(_21025_),
    .A2(_21026_),
    .B1(_21027_),
    .Y(_21029_));
 sky130_fd_sc_hd__and2_1 _49918_ (.A(_21028_),
    .B(_21029_),
    .X(_21030_));
 sky130_fd_sc_hd__or3_1 _49919_ (.A(_21013_),
    .B(_20999_),
    .C(_21002_),
    .X(_21031_));
 sky130_fd_sc_hd__nand3_1 _49920_ (.A(_21015_),
    .B(_21030_),
    .C(_21031_),
    .Y(_21032_));
 sky130_fd_sc_hd__a21o_1 _49921_ (.A1(_21031_),
    .A2(_21015_),
    .B1(_21030_),
    .X(_21033_));
 sky130_fd_sc_hd__and2_2 _49922_ (.A(_21032_),
    .B(_21033_),
    .X(_21034_));
 sky130_fd_sc_hd__or2b_1 _49923_ (.A(_19679_),
    .B_N(\delay_line[37][8] ),
    .X(_21035_));
 sky130_fd_sc_hd__buf_1 _49924_ (.A(\delay_line[37][8] ),
    .X(_21036_));
 sky130_fd_sc_hd__or2b_1 _49925_ (.A(_21036_),
    .B_N(_19679_),
    .X(_21037_));
 sky130_fd_sc_hd__and3b_1 _49926_ (.A_N(_18576_),
    .B(_19679_),
    .C(_20819_),
    .X(_21038_));
 sky130_fd_sc_hd__o2bb2a_1 _49927_ (.A1_N(_21035_),
    .A2_N(_21037_),
    .B1(_21038_),
    .B2(_20817_),
    .X(_21039_));
 sky130_fd_sc_hd__a21oi_1 _49928_ (.A1(_19678_),
    .A2(_20819_),
    .B1(_20817_),
    .Y(_21040_));
 sky130_fd_sc_hd__and3_1 _49929_ (.A(_21040_),
    .B(_21037_),
    .C(_21035_),
    .X(_21041_));
 sky130_fd_sc_hd__a31o_1 _49930_ (.A1(net292),
    .A2(_18569_),
    .A3(_19681_),
    .B1(_20823_),
    .X(_21042_));
 sky130_fd_sc_hd__or3_1 _49931_ (.A(_21039_),
    .B(_21041_),
    .C(_21042_),
    .X(_21043_));
 sky130_fd_sc_hd__o21ai_1 _49932_ (.A1(_21039_),
    .A2(_21041_),
    .B1(_21042_),
    .Y(_21044_));
 sky130_fd_sc_hd__nand2_1 _49933_ (.A(_21043_),
    .B(_21044_),
    .Y(_21045_));
 sky130_fd_sc_hd__buf_1 _49934_ (.A(\delay_line[36][4] ),
    .X(_21046_));
 sky130_fd_sc_hd__and3_1 _49935_ (.A(_18545_),
    .B(_21046_),
    .C(_19716_),
    .X(_21047_));
 sky130_fd_sc_hd__and2b_1 _49936_ (.A_N(_19715_),
    .B(\delay_line[36][5] ),
    .X(_21048_));
 sky130_fd_sc_hd__buf_1 _49937_ (.A(\delay_line[36][5] ),
    .X(_21049_));
 sky130_fd_sc_hd__and2b_1 _49938_ (.A_N(_21049_),
    .B(_19715_),
    .X(_21050_));
 sky130_fd_sc_hd__nor2_1 _49939_ (.A(_21048_),
    .B(_21050_),
    .Y(_21051_));
 sky130_fd_sc_hd__o21ba_1 _49940_ (.A1(_20828_),
    .A2(_20826_),
    .B1_N(_20825_),
    .X(_21052_));
 sky130_fd_sc_hd__xnor2_1 _49941_ (.A(_21051_),
    .B(_21052_),
    .Y(_21053_));
 sky130_fd_sc_hd__o21ai_2 _49942_ (.A1(net236),
    .A2(_21047_),
    .B1(_21053_),
    .Y(_21054_));
 sky130_fd_sc_hd__a311o_1 _49943_ (.A1(_18546_),
    .A2(_21046_),
    .A3(_19716_),
    .B1(net236),
    .C1(_21053_),
    .X(_21055_));
 sky130_fd_sc_hd__nand2_2 _49944_ (.A(_21054_),
    .B(_21055_),
    .Y(_21056_));
 sky130_fd_sc_hd__nor2_1 _49945_ (.A(\delay_line[35][7] ),
    .B(\delay_line[35][8] ),
    .Y(_21057_));
 sky130_fd_sc_hd__nand2_1 _49946_ (.A(\delay_line[35][7] ),
    .B(\delay_line[35][8] ),
    .Y(_21058_));
 sky130_fd_sc_hd__nand3b_1 _49947_ (.A_N(_21057_),
    .B(_21058_),
    .C(_20835_),
    .Y(_21059_));
 sky130_fd_sc_hd__and2_1 _49948_ (.A(\delay_line[35][7] ),
    .B(\delay_line[35][8] ),
    .X(_21060_));
 sky130_fd_sc_hd__o21bai_2 _49949_ (.A1(_21057_),
    .A2(_21060_),
    .B1_N(_19690_),
    .Y(_21061_));
 sky130_fd_sc_hd__o21a_1 _49950_ (.A1(_20835_),
    .A2(_20834_),
    .B1(_20833_),
    .X(_21062_));
 sky130_fd_sc_hd__a221oi_2 _49951_ (.A1(_20837_),
    .A2(_20834_),
    .B1(_21059_),
    .B2(_21061_),
    .C1(_21062_),
    .Y(_21063_));
 sky130_fd_sc_hd__inv_2 _49952_ (.A(_21063_),
    .Y(_21064_));
 sky130_fd_sc_hd__o211ai_2 _49953_ (.A1(_20840_),
    .A2(_21062_),
    .B1(_21059_),
    .C1(_21061_),
    .Y(_21065_));
 sky130_fd_sc_hd__and3_1 _49954_ (.A(_21064_),
    .B(_20841_),
    .C(_21065_),
    .X(_21066_));
 sky130_fd_sc_hd__a21o_1 _49955_ (.A1(_21065_),
    .A2(_21064_),
    .B1(_20841_),
    .X(_21067_));
 sky130_fd_sc_hd__inv_2 _49956_ (.A(_21067_),
    .Y(_21068_));
 sky130_fd_sc_hd__or3_1 _49957_ (.A(_04327_),
    .B(_21066_),
    .C(_21068_),
    .X(_21069_));
 sky130_fd_sc_hd__o21ai_1 _49958_ (.A1(_21066_),
    .A2(_21068_),
    .B1(_04338_),
    .Y(_21070_));
 sky130_fd_sc_hd__o211a_1 _49959_ (.A1(_20845_),
    .A2(_20847_),
    .B1(_21069_),
    .C1(_21070_),
    .X(_21071_));
 sky130_fd_sc_hd__a211oi_1 _49960_ (.A1(_21069_),
    .A2(_21070_),
    .B1(_20845_),
    .C1(_20847_),
    .Y(_21072_));
 sky130_fd_sc_hd__nor2_1 _49961_ (.A(_21071_),
    .B(_21072_),
    .Y(_21073_));
 sky130_fd_sc_hd__a21o_1 _49962_ (.A1(_20851_),
    .A2(_20850_),
    .B1(_20848_),
    .X(_21074_));
 sky130_fd_sc_hd__xnor2_2 _49963_ (.A(_21073_),
    .B(_21074_),
    .Y(_21075_));
 sky130_fd_sc_hd__xnor2_1 _49964_ (.A(_21056_),
    .B(_21075_),
    .Y(_21076_));
 sky130_fd_sc_hd__or2_2 _49965_ (.A(_21045_),
    .B(_21076_),
    .X(_21077_));
 sky130_fd_sc_hd__nand2_1 _49966_ (.A(_21045_),
    .B(_21076_),
    .Y(_21078_));
 sky130_fd_sc_hd__nand2_1 _49967_ (.A(_21077_),
    .B(_21078_),
    .Y(_21079_));
 sky130_fd_sc_hd__and3_1 _49968_ (.A(_20854_),
    .B(_20855_),
    .C(_21079_),
    .X(_21080_));
 sky130_fd_sc_hd__a21oi_1 _49969_ (.A1(_20854_),
    .A2(_20855_),
    .B1(_21079_),
    .Y(_21081_));
 sky130_fd_sc_hd__nor2_2 _49970_ (.A(_21080_),
    .B(_21081_),
    .Y(_21082_));
 sky130_fd_sc_hd__xnor2_4 _49971_ (.A(_21034_),
    .B(_21082_),
    .Y(_21083_));
 sky130_fd_sc_hd__and2_1 _49972_ (.A(\delay_line[34][6] ),
    .B(\delay_line[34][8] ),
    .X(_21084_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _49973_ (.A(\delay_line[34][8] ),
    .X(_21085_));
 sky130_fd_sc_hd__nor2_1 _49974_ (.A(_19549_),
    .B(_21085_),
    .Y(_21086_));
 sky130_fd_sc_hd__inv_2 _49975_ (.A(_20743_),
    .Y(_21087_));
 sky130_fd_sc_hd__o21ai_1 _49976_ (.A1(_21084_),
    .A2(_21086_),
    .B1(_21087_),
    .Y(_21088_));
 sky130_fd_sc_hd__nor2_1 _49977_ (.A(_20736_),
    .B(_20737_),
    .Y(_21089_));
 sky130_fd_sc_hd__nand2_1 _49978_ (.A(_19553_),
    .B(_21085_),
    .Y(_21090_));
 sky130_fd_sc_hd__nand3b_1 _49979_ (.A_N(_21086_),
    .B(_20741_),
    .C(_21090_),
    .Y(_21091_));
 sky130_fd_sc_hd__nand3_1 _49980_ (.A(_21088_),
    .B(_21089_),
    .C(_21091_),
    .Y(_21092_));
 sky130_fd_sc_hd__a2bb2o_1 _49981_ (.A1_N(_20736_),
    .A2_N(_20737_),
    .B1(_21091_),
    .B2(_21088_),
    .X(_21093_));
 sky130_fd_sc_hd__a32o_1 _49982_ (.A1(_20738_),
    .A2(_20740_),
    .A3(_20745_),
    .B1(_19551_),
    .B2(_21087_),
    .X(_21094_));
 sky130_fd_sc_hd__a21o_1 _49983_ (.A1(_21092_),
    .A2(_21093_),
    .B1(_21094_),
    .X(_21095_));
 sky130_fd_sc_hd__nand3_1 _49984_ (.A(_21094_),
    .B(_21092_),
    .C(_21093_),
    .Y(_21096_));
 sky130_fd_sc_hd__clkbuf_2 _49985_ (.A(_20739_),
    .X(_21097_));
 sky130_fd_sc_hd__a21oi_2 _49986_ (.A1(_21097_),
    .A2(_20740_),
    .B1(_00601_),
    .Y(_21098_));
 sky130_fd_sc_hd__and3_1 _49987_ (.A(_20740_),
    .B(_00601_),
    .C(_21097_),
    .X(_21099_));
 sky130_fd_sc_hd__or2_1 _49988_ (.A(_21098_),
    .B(_21099_),
    .X(_21100_));
 sky130_fd_sc_hd__a21o_1 _49989_ (.A1(_21095_),
    .A2(_21096_),
    .B1(_21100_),
    .X(_21101_));
 sky130_fd_sc_hd__o211ai_1 _49990_ (.A1(_21098_),
    .A2(_21099_),
    .B1(_21095_),
    .C1(_21096_),
    .Y(_21102_));
 sky130_fd_sc_hd__a21boi_1 _49991_ (.A1(_20750_),
    .A2(_20751_),
    .B1_N(_20748_),
    .Y(_21103_));
 sky130_fd_sc_hd__nand3_1 _49992_ (.A(_21101_),
    .B(_21102_),
    .C(_21103_),
    .Y(_21104_));
 sky130_fd_sc_hd__a21o_1 _49993_ (.A1(_21101_),
    .A2(_21102_),
    .B1(_21103_),
    .X(_21105_));
 sky130_fd_sc_hd__a21o_1 _49994_ (.A1(_21104_),
    .A2(_21105_),
    .B1(_20749_),
    .X(_21106_));
 sky130_fd_sc_hd__nand3_1 _49995_ (.A(_21105_),
    .B(_20749_),
    .C(_21104_),
    .Y(_21107_));
 sky130_fd_sc_hd__and2_1 _49996_ (.A(_21106_),
    .B(_21107_),
    .X(_21108_));
 sky130_fd_sc_hd__o21bai_2 _49997_ (.A1(_20755_),
    .A2(_20757_),
    .B1_N(_20756_),
    .Y(_21109_));
 sky130_fd_sc_hd__xor2_1 _49998_ (.A(_21108_),
    .B(_21109_),
    .X(_21110_));
 sky130_fd_sc_hd__nor2_1 _49999_ (.A(_20718_),
    .B(_20719_),
    .Y(_21111_));
 sky130_fd_sc_hd__clkbuf_2 _50000_ (.A(_20688_),
    .X(_21112_));
 sky130_fd_sc_hd__inv_2 _50001_ (.A(\delay_line[32][8] ),
    .Y(_21113_));
 sky130_fd_sc_hd__nand2_1 _50002_ (.A(_20690_),
    .B(_21113_),
    .Y(_21114_));
 sky130_fd_sc_hd__buf_1 _50003_ (.A(\delay_line[32][8] ),
    .X(_21115_));
 sky130_fd_sc_hd__buf_2 _50004_ (.A(_21115_),
    .X(_21116_));
 sky130_fd_sc_hd__nand2_1 _50005_ (.A(_20700_),
    .B(_21116_),
    .Y(_21117_));
 sky130_fd_sc_hd__o2111ai_4 _50006_ (.A1(_21112_),
    .A2(_20690_),
    .B1(_20696_),
    .C1(_21114_),
    .D1(_21117_),
    .Y(_21118_));
 sky130_fd_sc_hd__nor2_1 _50007_ (.A(_20700_),
    .B(_21116_),
    .Y(_21119_));
 sky130_fd_sc_hd__and2_1 _50008_ (.A(_20686_),
    .B(_21115_),
    .X(_21120_));
 sky130_fd_sc_hd__o2bb2ai_1 _50009_ (.A1_N(_20687_),
    .A2_N(_20696_),
    .B1(_21119_),
    .B2(_21120_),
    .Y(_21121_));
 sky130_fd_sc_hd__nor2_1 _50010_ (.A(_19586_),
    .B(_19587_),
    .Y(_21122_));
 sky130_fd_sc_hd__nand3_2 _50011_ (.A(_21118_),
    .B(_21121_),
    .C(_21122_),
    .Y(_21123_));
 sky130_fd_sc_hd__a21o_1 _50012_ (.A1(_21118_),
    .A2(_21121_),
    .B1(_21122_),
    .X(_21124_));
 sky130_fd_sc_hd__o2bb2ai_2 _50013_ (.A1_N(_21123_),
    .A2_N(_21124_),
    .B1(_20693_),
    .B2(_20698_),
    .Y(_21125_));
 sky130_fd_sc_hd__buf_2 _50014_ (.A(_20700_),
    .X(_21126_));
 sky130_fd_sc_hd__a21o_1 _50015_ (.A1(_20699_),
    .A2(_21126_),
    .B1(_20696_),
    .X(_21127_));
 sky130_fd_sc_hd__a21oi_2 _50016_ (.A1(_21127_),
    .A2(_20705_),
    .B1(_20697_),
    .Y(_21128_));
 sky130_fd_sc_hd__o22ai_1 _50017_ (.A1(_20693_),
    .A2(_20698_),
    .B1(_18672_),
    .B2(_21128_),
    .Y(_21129_));
 sky130_fd_sc_hd__nand3_2 _50018_ (.A(_21123_),
    .B(_21124_),
    .C(_21129_),
    .Y(_21130_));
 sky130_fd_sc_hd__o211a_1 _50019_ (.A1(_20703_),
    .A2(_21125_),
    .B1(_02106_),
    .C1(_21130_),
    .X(_21131_));
 sky130_fd_sc_hd__nand2_1 _50020_ (.A(_21123_),
    .B(_21124_),
    .Y(_21132_));
 sky130_fd_sc_hd__o221ai_4 _50021_ (.A1(_19611_),
    .A2(_21128_),
    .B1(_20698_),
    .B2(_20693_),
    .C1(_21132_),
    .Y(_21133_));
 sky130_fd_sc_hd__a21oi_1 _50022_ (.A1(_21130_),
    .A2(_21133_),
    .B1(_02117_),
    .Y(_21134_));
 sky130_fd_sc_hd__a21boi_1 _50023_ (.A1(_20709_),
    .A2(_24468_),
    .B1_N(_20712_),
    .Y(_21135_));
 sky130_fd_sc_hd__o21ai_1 _50024_ (.A1(_21131_),
    .A2(_21134_),
    .B1(_21135_),
    .Y(_21136_));
 sky130_fd_sc_hd__a21oi_1 _50025_ (.A1(_20710_),
    .A2(_20711_),
    .B1(_20708_),
    .Y(_21137_));
 sky130_fd_sc_hd__o21ai_2 _50026_ (.A1(_24545_),
    .A2(_21137_),
    .B1(_20714_),
    .Y(_21138_));
 sky130_fd_sc_hd__o211ai_4 _50027_ (.A1(_20703_),
    .A2(_21125_),
    .B1(_02117_),
    .C1(_21130_),
    .Y(_21139_));
 sky130_fd_sc_hd__a21o_1 _50028_ (.A1(_21130_),
    .A2(_21133_),
    .B1(_02117_),
    .X(_21140_));
 sky130_fd_sc_hd__nand3_2 _50029_ (.A(_21138_),
    .B(_21139_),
    .C(_21140_),
    .Y(_21141_));
 sky130_fd_sc_hd__nand4_1 _50030_ (.A(_21111_),
    .B(_20716_),
    .C(_21136_),
    .D(_21141_),
    .Y(_21142_));
 sky130_fd_sc_hd__nand2_1 _50031_ (.A(_20713_),
    .B(_20715_),
    .Y(_21143_));
 sky130_fd_sc_hd__o2bb2ai_2 _50032_ (.A1_N(_21136_),
    .A2_N(_21141_),
    .B1(_20720_),
    .B2(_21143_),
    .Y(_21144_));
 sky130_fd_sc_hd__a21o_1 _50033_ (.A1(_21142_),
    .A2(_21144_),
    .B1(_24501_),
    .X(_21145_));
 sky130_fd_sc_hd__o221a_1 _50034_ (.A1(_21137_),
    .A2(_24545_),
    .B1(_21134_),
    .B2(_21131_),
    .C1(_20714_),
    .X(_21146_));
 sky130_fd_sc_hd__nand4_2 _50035_ (.A(_20713_),
    .B(_20715_),
    .C(_20716_),
    .D(_21141_),
    .Y(_21147_));
 sky130_fd_sc_hd__o211ai_2 _50036_ (.A1(_21146_),
    .A2(_21147_),
    .B1(_21144_),
    .C1(_24512_),
    .Y(_21148_));
 sky130_fd_sc_hd__a21oi_1 _50037_ (.A1(_20713_),
    .A2(_20715_),
    .B1(_20716_),
    .Y(_21149_));
 sky130_fd_sc_hd__nand3_1 _50038_ (.A(_20717_),
    .B(_19616_),
    .C(_19613_),
    .Y(_21150_));
 sky130_fd_sc_hd__nor2_1 _50039_ (.A(_21149_),
    .B(_21150_),
    .Y(_21151_));
 sky130_fd_sc_hd__a21oi_1 _50040_ (.A1(_21145_),
    .A2(_21148_),
    .B1(_21151_),
    .Y(_21152_));
 sky130_fd_sc_hd__inv_2 _50041_ (.A(_19610_),
    .Y(_21153_));
 sky130_fd_sc_hd__o22ai_1 _50042_ (.A1(_20722_),
    .A2(_21153_),
    .B1(_20726_),
    .B2(_21151_),
    .Y(_21154_));
 sky130_fd_sc_hd__a21oi_1 _50043_ (.A1(_21154_),
    .A2(_19618_),
    .B1(_20728_),
    .Y(_21155_));
 sky130_fd_sc_hd__nor2_1 _50044_ (.A(_21152_),
    .B(_21155_),
    .Y(_21156_));
 sky130_fd_sc_hd__and3_1 _50045_ (.A(_21145_),
    .B(_21148_),
    .C(_21151_),
    .X(_21157_));
 sky130_fd_sc_hd__o221a_1 _50046_ (.A1(_20727_),
    .A2(_20726_),
    .B1(_21152_),
    .B2(_21157_),
    .C1(_20731_),
    .X(_21158_));
 sky130_fd_sc_hd__nand3b_1 _50047_ (.A_N(_02161_),
    .B(_20674_),
    .C(_00568_),
    .Y(_21159_));
 sky130_fd_sc_hd__a21oi_1 _50048_ (.A1(_19570_),
    .A2(_05337_),
    .B1(_20667_),
    .Y(_21160_));
 sky130_fd_sc_hd__clkbuf_2 _50049_ (.A(\delay_line[33][8] ),
    .X(_21161_));
 sky130_fd_sc_hd__xnor2_1 _50050_ (.A(_17822_),
    .B(_21161_),
    .Y(_21162_));
 sky130_fd_sc_hd__o21a_1 _50051_ (.A1(_20670_),
    .A2(_21160_),
    .B1(_21162_),
    .X(_21163_));
 sky130_fd_sc_hd__o22a_1 _50052_ (.A1(_02161_),
    .A2(_05337_),
    .B1(_21160_),
    .B2(_21162_),
    .X(_21164_));
 sky130_fd_sc_hd__nor2_1 _50053_ (.A(_20670_),
    .B(_21164_),
    .Y(_21165_));
 sky130_fd_sc_hd__o2bb2ai_2 _50054_ (.A1_N(_20673_),
    .A2_N(_21159_),
    .B1(_21163_),
    .B2(_21165_),
    .Y(_21166_));
 sky130_fd_sc_hd__o21ai_1 _50055_ (.A1(_20670_),
    .A2(_21160_),
    .B1(_21162_),
    .Y(_21167_));
 sky130_fd_sc_hd__o2111ai_2 _50056_ (.A1(_20670_),
    .A2(_21164_),
    .B1(_21167_),
    .C1(_20673_),
    .D1(_21159_),
    .Y(_21168_));
 sky130_fd_sc_hd__nand4_2 _50057_ (.A(_21166_),
    .B(_00579_),
    .C(_21168_),
    .D(_02172_),
    .Y(_21169_));
 sky130_fd_sc_hd__a22o_1 _50058_ (.A1(_00579_),
    .A2(_02172_),
    .B1(_21168_),
    .B2(_21166_),
    .X(_21170_));
 sky130_fd_sc_hd__nand2_1 _50059_ (.A(_20682_),
    .B(_20681_),
    .Y(_21171_));
 sky130_fd_sc_hd__nand3_1 _50060_ (.A(_21169_),
    .B(_21170_),
    .C(_21171_),
    .Y(_21172_));
 sky130_fd_sc_hd__a21o_1 _50061_ (.A1(_21169_),
    .A2(_21170_),
    .B1(_21171_),
    .X(_21173_));
 sky130_fd_sc_hd__nand2_1 _50062_ (.A(_21172_),
    .B(_21173_),
    .Y(_21174_));
 sky130_fd_sc_hd__a21oi_2 _50063_ (.A1(_21174_),
    .A2(_22534_),
    .B1(_20684_),
    .Y(_21175_));
 sky130_fd_sc_hd__xnor2_1 _50064_ (.A(_22534_),
    .B(_21174_),
    .Y(_21176_));
 sky130_fd_sc_hd__and2_1 _50065_ (.A(_20684_),
    .B(_21176_),
    .X(_21177_));
 sky130_fd_sc_hd__nor2_1 _50066_ (.A(_21175_),
    .B(_21177_),
    .Y(_21178_));
 sky130_fd_sc_hd__o21bai_1 _50067_ (.A1(_21156_),
    .A2(_21158_),
    .B1_N(_21178_),
    .Y(_21179_));
 sky130_fd_sc_hd__or3b_2 _50068_ (.A(_21156_),
    .B(_21158_),
    .C_N(_21178_),
    .X(_21180_));
 sky130_fd_sc_hd__and2_1 _50069_ (.A(_21179_),
    .B(_21180_),
    .X(_21181_));
 sky130_fd_sc_hd__nand2_1 _50070_ (.A(_21110_),
    .B(_21181_),
    .Y(_21182_));
 sky130_fd_sc_hd__or2_1 _50071_ (.A(_21110_),
    .B(_21181_),
    .X(_21183_));
 sky130_fd_sc_hd__nand2_1 _50072_ (.A(_21182_),
    .B(_21183_),
    .Y(_21184_));
 sky130_fd_sc_hd__and3_1 _50073_ (.A(_20366_),
    .B(_20369_),
    .C(_21184_),
    .X(_21185_));
 sky130_fd_sc_hd__a21oi_1 _50074_ (.A1(_20366_),
    .A2(_20369_),
    .B1(_21184_),
    .Y(_21186_));
 sky130_fd_sc_hd__nor2_1 _50075_ (.A(_21185_),
    .B(_21186_),
    .Y(_21187_));
 sky130_fd_sc_hd__nand2_1 _50076_ (.A(_20761_),
    .B(_20762_),
    .Y(_21188_));
 sky130_fd_sc_hd__xor2_1 _50077_ (.A(_21187_),
    .B(_21188_),
    .X(_21189_));
 sky130_fd_sc_hd__a211oi_1 _50078_ (.A1(_20766_),
    .A2(_20665_),
    .B1(_20765_),
    .C1(_21189_),
    .Y(_21190_));
 sky130_fd_sc_hd__and2_1 _50079_ (.A(_20766_),
    .B(_20665_),
    .X(_21191_));
 sky130_fd_sc_hd__o21ai_1 _50080_ (.A1(_20765_),
    .A2(_21191_),
    .B1(_21189_),
    .Y(_21192_));
 sky130_fd_sc_hd__or3b_1 _50081_ (.A(_21083_),
    .B(_21190_),
    .C_N(_21192_),
    .X(_21193_));
 sky130_fd_sc_hd__or2b_1 _50082_ (.A(_21190_),
    .B_N(_21192_),
    .X(_21194_));
 sky130_fd_sc_hd__nand2_1 _50083_ (.A(_21083_),
    .B(_21194_),
    .Y(_21195_));
 sky130_fd_sc_hd__nand2_1 _50084_ (.A(_21193_),
    .B(_21195_),
    .Y(_21196_));
 sky130_fd_sc_hd__o21a_1 _50085_ (.A1(_20301_),
    .A2(_20443_),
    .B1(_20448_),
    .X(_21197_));
 sky130_fd_sc_hd__xnor2_1 _50086_ (.A(_21196_),
    .B(_21197_),
    .Y(_21198_));
 sky130_fd_sc_hd__or2b_1 _50087_ (.A(_20984_),
    .B_N(_21198_),
    .X(_21199_));
 sky130_fd_sc_hd__or2b_1 _50088_ (.A(_21198_),
    .B_N(_20984_),
    .X(_21200_));
 sky130_fd_sc_hd__a21o_2 _50089_ (.A1(_20371_),
    .A2(_20442_),
    .B1(_20441_),
    .X(_21201_));
 sky130_fd_sc_hd__nand3_2 _50090_ (.A(_20426_),
    .B(_20432_),
    .C(_20434_),
    .Y(_21202_));
 sky130_fd_sc_hd__a21o_1 _50091_ (.A1(_19300_),
    .A2(_20410_),
    .B1(\delay_line[28][8] ),
    .X(_21203_));
 sky130_fd_sc_hd__buf_1 _50092_ (.A(\delay_line[28][8] ),
    .X(_21204_));
 sky130_fd_sc_hd__nand3_1 _50093_ (.A(_19301_),
    .B(_20407_),
    .C(_21204_),
    .Y(_21205_));
 sky130_fd_sc_hd__a21o_1 _50094_ (.A1(_21203_),
    .A2(_21205_),
    .B1(\delay_line[28][3] ),
    .X(_21206_));
 sky130_fd_sc_hd__nand3_1 _50095_ (.A(_21203_),
    .B(_21205_),
    .C(_06414_),
    .Y(_21207_));
 sky130_fd_sc_hd__a2bb2o_1 _50096_ (.A1_N(_20407_),
    .A2_N(_20408_),
    .B1(\delay_line[28][2] ),
    .B2(_20412_),
    .X(_21208_));
 sky130_fd_sc_hd__a21o_1 _50097_ (.A1(_21206_),
    .A2(_21207_),
    .B1(_21208_),
    .X(_21209_));
 sky130_fd_sc_hd__nand3_2 _50098_ (.A(_21208_),
    .B(_21206_),
    .C(_21207_),
    .Y(_21210_));
 sky130_fd_sc_hd__and3_1 _50099_ (.A(_21209_),
    .B(_21210_),
    .C(_01117_),
    .X(_21211_));
 sky130_fd_sc_hd__a21oi_2 _50100_ (.A1(_21209_),
    .A2(_21210_),
    .B1(_01128_),
    .Y(_21212_));
 sky130_fd_sc_hd__a211oi_4 _50101_ (.A1(_20418_),
    .A2(_20419_),
    .B1(_21211_),
    .C1(_21212_),
    .Y(_21213_));
 sky130_fd_sc_hd__a21oi_1 _50102_ (.A1(_20417_),
    .A2(_24380_),
    .B1(_20433_),
    .Y(_21214_));
 sky130_fd_sc_hd__o21ai_1 _50103_ (.A1(_21211_),
    .A2(_21212_),
    .B1(_21214_),
    .Y(_21215_));
 sky130_fd_sc_hd__inv_2 _50104_ (.A(_21215_),
    .Y(_21216_));
 sky130_fd_sc_hd__o21ai_4 _50105_ (.A1(_21213_),
    .A2(_21216_),
    .B1(_20425_),
    .Y(_21217_));
 sky130_fd_sc_hd__nor3_2 _50106_ (.A(_20425_),
    .B(_21213_),
    .C(_21216_),
    .Y(_21218_));
 sky130_fd_sc_hd__and2b_1 _50107_ (.A_N(_21218_),
    .B(_21217_),
    .X(_21219_));
 sky130_fd_sc_hd__nor2_1 _50108_ (.A(_21202_),
    .B(_21219_),
    .Y(_21220_));
 sky130_fd_sc_hd__a21oi_1 _50109_ (.A1(_21202_),
    .A2(_21217_),
    .B1(_21220_),
    .Y(_21221_));
 sky130_fd_sc_hd__o21a_1 _50110_ (.A1(_18485_),
    .A2(net339),
    .B1(_01161_),
    .X(_21222_));
 sky130_fd_sc_hd__inv_2 _50111_ (.A(_16009_),
    .Y(_21223_));
 sky130_fd_sc_hd__nor2_1 _50112_ (.A(net339),
    .B(_21223_),
    .Y(_21224_));
 sky130_fd_sc_hd__nor2_1 _50113_ (.A(_16009_),
    .B(_06469_),
    .Y(_21225_));
 sky130_fd_sc_hd__or3_1 _50114_ (.A(_21222_),
    .B(_21224_),
    .C(_21225_),
    .X(_21226_));
 sky130_fd_sc_hd__o21ai_1 _50115_ (.A1(_21224_),
    .A2(_21225_),
    .B1(_21222_),
    .Y(_21227_));
 sky130_fd_sc_hd__clkbuf_2 _50116_ (.A(\delay_line[26][7] ),
    .X(_21228_));
 sky130_fd_sc_hd__and3_2 _50117_ (.A(_21226_),
    .B(_21227_),
    .C(_21228_),
    .X(_21229_));
 sky130_fd_sc_hd__a21oi_2 _50118_ (.A1(_21226_),
    .A2(_21227_),
    .B1(_21228_),
    .Y(_21230_));
 sky130_fd_sc_hd__a211oi_4 _50119_ (.A1(_20399_),
    .A2(_20401_),
    .B1(_21229_),
    .C1(_21230_),
    .Y(_21231_));
 sky130_fd_sc_hd__o211a_1 _50120_ (.A1(_21229_),
    .A2(_21230_),
    .B1(_20399_),
    .C1(_20401_),
    .X(_21232_));
 sky130_fd_sc_hd__o21a_1 _50121_ (.A1(_20382_),
    .A2(_20383_),
    .B1(_20384_),
    .X(_21233_));
 sky130_fd_sc_hd__o21ai_1 _50122_ (.A1(_20372_),
    .A2(_21233_),
    .B1(_20389_),
    .Y(_21234_));
 sky130_fd_sc_hd__clkbuf_2 _50123_ (.A(\delay_line[27][8] ),
    .X(_21235_));
 sky130_fd_sc_hd__nand4b_2 _50124_ (.A_N(_20375_),
    .B(_20378_),
    .C(_21235_),
    .D(_19279_),
    .Y(_21236_));
 sky130_fd_sc_hd__nor2_1 _50125_ (.A(net332),
    .B(\delay_line[27][8] ),
    .Y(_21237_));
 sky130_fd_sc_hd__nand2_1 _50126_ (.A(_19273_),
    .B(_21235_),
    .Y(_21238_));
 sky130_fd_sc_hd__nand3b_1 _50127_ (.A_N(_21237_),
    .B(_21238_),
    .C(_20376_),
    .Y(_21239_));
 sky130_fd_sc_hd__and2_1 _50128_ (.A(net332),
    .B(\delay_line[27][8] ),
    .X(_21240_));
 sky130_fd_sc_hd__o21ai_2 _50129_ (.A1(_21237_),
    .A2(_21240_),
    .B1(_20378_),
    .Y(_21241_));
 sky130_fd_sc_hd__nand3_2 _50130_ (.A(_20379_),
    .B(_21239_),
    .C(_21241_),
    .Y(_21242_));
 sky130_fd_sc_hd__nand3b_2 _50131_ (.A_N(_01205_),
    .B(_21236_),
    .C(_21242_),
    .Y(_21243_));
 sky130_fd_sc_hd__a21bo_1 _50132_ (.A1(_21236_),
    .A2(_21242_),
    .B1_N(_01194_),
    .X(_21244_));
 sky130_fd_sc_hd__o211a_1 _50133_ (.A1(_20374_),
    .A2(_20382_),
    .B1(_21243_),
    .C1(_21244_),
    .X(_21245_));
 sky130_fd_sc_hd__a211oi_4 _50134_ (.A1(_21243_),
    .A2(_21244_),
    .B1(_20374_),
    .C1(_20382_),
    .Y(_21246_));
 sky130_fd_sc_hd__nor2_1 _50135_ (.A(_21245_),
    .B(_21246_),
    .Y(_21247_));
 sky130_fd_sc_hd__nand2_1 _50136_ (.A(_21234_),
    .B(_21247_),
    .Y(_21248_));
 sky130_fd_sc_hd__o221ai_1 _50137_ (.A1(_20372_),
    .A2(_21233_),
    .B1(_21245_),
    .B2(_21246_),
    .C1(_20389_),
    .Y(_21249_));
 sky130_fd_sc_hd__nand2_1 _50138_ (.A(_21248_),
    .B(_21249_),
    .Y(_21250_));
 sky130_fd_sc_hd__xnor2_1 _50139_ (.A(_20394_),
    .B(_21250_),
    .Y(_21251_));
 sky130_fd_sc_hd__o21ai_1 _50140_ (.A1(_21231_),
    .A2(_21232_),
    .B1(_21251_),
    .Y(_21252_));
 sky130_fd_sc_hd__o211ai_1 _50141_ (.A1(_21229_),
    .A2(_21230_),
    .B1(_20399_),
    .C1(_20401_),
    .Y(_21253_));
 sky130_fd_sc_hd__or3b_1 _50142_ (.A(_21231_),
    .B(_21251_),
    .C_N(_21253_),
    .X(_21254_));
 sky130_fd_sc_hd__nand2_2 _50143_ (.A(_21252_),
    .B(_21254_),
    .Y(_21255_));
 sky130_fd_sc_hd__xor2_2 _50144_ (.A(_21221_),
    .B(_21255_),
    .X(_21256_));
 sky130_fd_sc_hd__a21oi_2 _50145_ (.A1(_20404_),
    .A2(_20436_),
    .B1(_21256_),
    .Y(_21257_));
 sky130_fd_sc_hd__nand3_2 _50146_ (.A(_20404_),
    .B(_20436_),
    .C(_21256_),
    .Y(_21258_));
 sky130_fd_sc_hd__or2b_2 _50147_ (.A(_21257_),
    .B_N(_21258_),
    .X(_21259_));
 sky130_fd_sc_hd__nor2_1 _50148_ (.A(_19375_),
    .B(_20326_),
    .Y(_21260_));
 sky130_fd_sc_hd__nand2_1 _50149_ (.A(_19351_),
    .B(_20303_),
    .Y(_21261_));
 sky130_fd_sc_hd__inv_2 _50150_ (.A(\delay_line[31][8] ),
    .Y(_21262_));
 sky130_fd_sc_hd__nand2_1 _50151_ (.A(_20308_),
    .B(_21262_),
    .Y(_21263_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50152_ (.A(\delay_line[31][8] ),
    .X(_21264_));
 sky130_fd_sc_hd__nand2_1 _50153_ (.A(_20303_),
    .B(_21264_),
    .Y(_21265_));
 sky130_fd_sc_hd__nand4_2 _50154_ (.A(_21261_),
    .B(_20305_),
    .C(_21263_),
    .D(_21265_),
    .Y(_21266_));
 sky130_fd_sc_hd__nor2_1 _50155_ (.A(_20303_),
    .B(\delay_line[31][8] ),
    .Y(_21267_));
 sky130_fd_sc_hd__and2_1 _50156_ (.A(\delay_line[31][7] ),
    .B(\delay_line[31][8] ),
    .X(_21268_));
 sky130_fd_sc_hd__o2bb2ai_4 _50157_ (.A1_N(_21261_),
    .A2_N(_20305_),
    .B1(_21267_),
    .B2(_21268_),
    .Y(_21269_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50158_ (.A(_20302_),
    .X(_21270_));
 sky130_fd_sc_hd__and3_1 _50159_ (.A(_21266_),
    .B(_21269_),
    .C(_21270_),
    .X(_21271_));
 sky130_fd_sc_hd__a21oi_1 _50160_ (.A1(_21266_),
    .A2(_21269_),
    .B1(_20302_),
    .Y(_21272_));
 sky130_fd_sc_hd__o21ai_2 _50161_ (.A1(_21271_),
    .A2(_21272_),
    .B1(_20318_),
    .Y(_21273_));
 sky130_fd_sc_hd__nand3_2 _50162_ (.A(_21266_),
    .B(_21269_),
    .C(_21270_),
    .Y(_21274_));
 sky130_fd_sc_hd__nand3b_1 _50163_ (.A_N(_21272_),
    .B(_20312_),
    .C(_21274_),
    .Y(_21275_));
 sky130_fd_sc_hd__buf_1 _50164_ (.A(_21275_),
    .X(_21276_));
 sky130_fd_sc_hd__a21o_1 _50165_ (.A1(_21273_),
    .A2(_21276_),
    .B1(_15712_),
    .X(_21277_));
 sky130_fd_sc_hd__nand3_1 _50166_ (.A(_15712_),
    .B(_21273_),
    .C(_21276_),
    .Y(_21278_));
 sky130_fd_sc_hd__a21boi_1 _50167_ (.A1(_20316_),
    .A2(_20317_),
    .B1_N(_20319_),
    .Y(_21279_));
 sky130_fd_sc_hd__nand3_1 _50168_ (.A(_21277_),
    .B(_21278_),
    .C(_21279_),
    .Y(_21280_));
 sky130_fd_sc_hd__nand3_1 _50169_ (.A(_21273_),
    .B(_21276_),
    .C(_00985_),
    .Y(_21281_));
 sky130_fd_sc_hd__a21o_1 _50170_ (.A1(_21273_),
    .A2(_21275_),
    .B1(_00985_),
    .X(_21282_));
 sky130_fd_sc_hd__nand3b_2 _50171_ (.A_N(_21279_),
    .B(_21281_),
    .C(_21282_),
    .Y(_21283_));
 sky130_fd_sc_hd__nand2_1 _50172_ (.A(_20320_),
    .B(_20321_),
    .Y(_21284_));
 sky130_fd_sc_hd__o41a_1 _50173_ (.A1(_18473_),
    .A2(_19362_),
    .A3(_19364_),
    .A4(_19363_),
    .B1(_19367_),
    .X(_21285_));
 sky130_fd_sc_hd__o2bb2ai_2 _50174_ (.A1_N(_21280_),
    .A2_N(_21283_),
    .B1(_21284_),
    .B2(_21285_),
    .Y(_21286_));
 sky130_fd_sc_hd__nand3b_1 _50175_ (.A_N(_20323_),
    .B(_21280_),
    .C(_21283_),
    .Y(_21287_));
 sky130_fd_sc_hd__buf_1 _50176_ (.A(_21287_),
    .X(_21288_));
 sky130_fd_sc_hd__nand3b_1 _50177_ (.A_N(_19369_),
    .B(_20323_),
    .C(_20324_),
    .Y(_21289_));
 sky130_fd_sc_hd__a31oi_1 _50178_ (.A1(_21286_),
    .A2(_24567_),
    .A3(_21288_),
    .B1(_21289_),
    .Y(_21290_));
 sky130_fd_sc_hd__a21o_1 _50179_ (.A1(_21288_),
    .A2(_21286_),
    .B1(_24567_),
    .X(_21291_));
 sky130_fd_sc_hd__nor2_1 _50180_ (.A(_19369_),
    .B(_20326_),
    .Y(_21292_));
 sky130_fd_sc_hd__a31oi_1 _50181_ (.A1(_22237_),
    .A2(_21288_),
    .A3(_21286_),
    .B1(_21292_),
    .Y(_21293_));
 sky130_fd_sc_hd__a21o_1 _50182_ (.A1(_21287_),
    .A2(_21286_),
    .B1(_22226_),
    .X(_21294_));
 sky130_fd_sc_hd__a22o_1 _50183_ (.A1(_21290_),
    .A2(_21291_),
    .B1(_21293_),
    .B2(_21294_),
    .X(_21295_));
 sky130_fd_sc_hd__o21a_1 _50184_ (.A1(_20331_),
    .A2(_21260_),
    .B1(_21295_),
    .X(_21296_));
 sky130_fd_sc_hd__or3_1 _50185_ (.A(_20331_),
    .B(_21260_),
    .C(_21295_),
    .X(_21297_));
 sky130_fd_sc_hd__and2b_1 _50186_ (.A_N(_21296_),
    .B(_21297_),
    .X(_21298_));
 sky130_fd_sc_hd__or2b_1 _50187_ (.A(\delay_line[29][2] ),
    .B_N(\delay_line[29][6] ),
    .X(_21299_));
 sky130_fd_sc_hd__buf_1 _50188_ (.A(\delay_line[29][6] ),
    .X(_21300_));
 sky130_fd_sc_hd__or2b_1 _50189_ (.A(_21300_),
    .B_N(_15646_),
    .X(_21301_));
 sky130_fd_sc_hd__a221oi_2 _50190_ (.A1(_19322_),
    .A2(_20332_),
    .B1(_21299_),
    .B2(_21301_),
    .C1(_20335_),
    .Y(_21302_));
 sky130_fd_sc_hd__o211a_1 _50191_ (.A1(_20334_),
    .A2(_20335_),
    .B1(_21299_),
    .C1(_21301_),
    .X(_21303_));
 sky130_fd_sc_hd__nor3_1 _50192_ (.A(_21302_),
    .B(_21303_),
    .C(_20337_),
    .Y(_21304_));
 sky130_fd_sc_hd__o21a_1 _50193_ (.A1(_21302_),
    .A2(_21303_),
    .B1(_20337_),
    .X(_21305_));
 sky130_fd_sc_hd__nand2_1 _50194_ (.A(_24611_),
    .B(_06326_),
    .Y(_21306_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50195_ (.A(\delay_line[30][8] ),
    .X(_21307_));
 sky130_fd_sc_hd__inv_2 _50196_ (.A(_21307_),
    .Y(_21308_));
 sky130_fd_sc_hd__nand2_1 _50197_ (.A(_21308_),
    .B(\delay_line[30][5] ),
    .Y(_21309_));
 sky130_fd_sc_hd__inv_2 _50198_ (.A(\delay_line[30][5] ),
    .Y(_21310_));
 sky130_fd_sc_hd__nand2_1 _50199_ (.A(_21310_),
    .B(_21307_),
    .Y(_21311_));
 sky130_fd_sc_hd__o2111ai_4 _50200_ (.A1(_20346_),
    .A2(_20347_),
    .B1(_21309_),
    .C1(_21311_),
    .D1(_20348_),
    .Y(_21312_));
 sky130_fd_sc_hd__nand2_1 _50201_ (.A(_20341_),
    .B(_20344_),
    .Y(_21313_));
 sky130_fd_sc_hd__a22o_2 _50202_ (.A1(_21309_),
    .A2(_21311_),
    .B1(_21313_),
    .B2(_20348_),
    .X(_21314_));
 sky130_fd_sc_hd__a21oi_1 _50203_ (.A1(_20343_),
    .A2(_01018_),
    .B1(_06315_),
    .Y(_21315_));
 sky130_fd_sc_hd__and3_1 _50204_ (.A(_20343_),
    .B(_06304_),
    .C(_01018_),
    .X(_21316_));
 sky130_fd_sc_hd__o2bb2ai_2 _50205_ (.A1_N(_21312_),
    .A2_N(_21314_),
    .B1(_21315_),
    .B2(_21316_),
    .Y(_21317_));
 sky130_fd_sc_hd__and2_1 _50206_ (.A(_20344_),
    .B(_06304_),
    .X(_21318_));
 sky130_fd_sc_hd__nor2_1 _50207_ (.A(_06304_),
    .B(_20344_),
    .Y(_21319_));
 sky130_fd_sc_hd__o211ai_4 _50208_ (.A1(_21318_),
    .A2(_21319_),
    .B1(_21312_),
    .C1(_21314_),
    .Y(_21320_));
 sky130_fd_sc_hd__a21boi_1 _50209_ (.A1(_20345_),
    .A2(_20349_),
    .B1_N(_19337_),
    .Y(_21321_));
 sky130_fd_sc_hd__o21ai_2 _50210_ (.A1(_19330_),
    .A2(_21321_),
    .B1(_20353_),
    .Y(_21322_));
 sky130_fd_sc_hd__a21oi_1 _50211_ (.A1(_21317_),
    .A2(_21320_),
    .B1(_21322_),
    .Y(_21323_));
 sky130_fd_sc_hd__nand3_1 _50212_ (.A(_21322_),
    .B(_21317_),
    .C(_21320_),
    .Y(_21324_));
 sky130_fd_sc_hd__nor3b_1 _50213_ (.A(_21306_),
    .B(_21323_),
    .C_N(_21324_),
    .Y(_21325_));
 sky130_fd_sc_hd__a21o_1 _50214_ (.A1(_21317_),
    .A2(_21320_),
    .B1(_21322_),
    .X(_21326_));
 sky130_fd_sc_hd__a22o_1 _50215_ (.A1(_24611_),
    .A2(_06326_),
    .B1(_21326_),
    .B2(_21324_),
    .X(_21327_));
 sky130_fd_sc_hd__nand2_1 _50216_ (.A(_22281_),
    .B(_01029_),
    .Y(_21328_));
 sky130_fd_sc_hd__a21oi_1 _50217_ (.A1(_20354_),
    .A2(_20355_),
    .B1(_20356_),
    .Y(_21329_));
 sky130_fd_sc_hd__o21ai_1 _50218_ (.A1(_21328_),
    .A2(_21329_),
    .B1(_20358_),
    .Y(_21330_));
 sky130_fd_sc_hd__nand3b_1 _50219_ (.A_N(_21325_),
    .B(_21327_),
    .C(_21330_),
    .Y(_21331_));
 sky130_fd_sc_hd__a22oi_1 _50220_ (.A1(_24622_),
    .A2(_06326_),
    .B1(_21326_),
    .B2(_21324_),
    .Y(_21332_));
 sky130_fd_sc_hd__o21a_1 _50221_ (.A1(_21328_),
    .A2(_21329_),
    .B1(_20358_),
    .X(_21333_));
 sky130_fd_sc_hd__o21ai_1 _50222_ (.A1(_21325_),
    .A2(_21332_),
    .B1(_21333_),
    .Y(_21334_));
 sky130_fd_sc_hd__nand3_1 _50223_ (.A(_19327_),
    .B(_21331_),
    .C(_21334_),
    .Y(_21335_));
 sky130_fd_sc_hd__a21o_1 _50224_ (.A1(_21331_),
    .A2(_21334_),
    .B1(_19327_),
    .X(_21336_));
 sky130_fd_sc_hd__a2bb2oi_1 _50225_ (.A1_N(_19347_),
    .A2_N(_20360_),
    .B1(_21335_),
    .B2(_21336_),
    .Y(_21337_));
 sky130_fd_sc_hd__a2bb2o_1 _50226_ (.A1_N(_19347_),
    .A2_N(_20361_),
    .B1(_21335_),
    .B2(_21336_),
    .X(_21338_));
 sky130_fd_sc_hd__nor2_1 _50227_ (.A(_19344_),
    .B(_20360_),
    .Y(_21339_));
 sky130_fd_sc_hd__nand3_1 _50228_ (.A(_21336_),
    .B(_21339_),
    .C(_21335_),
    .Y(_21340_));
 sky130_fd_sc_hd__a2bb2o_1 _50229_ (.A1_N(_19345_),
    .A2_N(_20361_),
    .B1(_21338_),
    .B2(_21340_),
    .X(_21341_));
 sky130_fd_sc_hd__o31a_1 _50230_ (.A1(_19346_),
    .A2(_20361_),
    .A3(_21337_),
    .B1(_21341_),
    .X(_21342_));
 sky130_fd_sc_hd__o21bai_1 _50231_ (.A1(net235),
    .A2(_21305_),
    .B1_N(_21342_),
    .Y(_21343_));
 sky130_fd_sc_hd__or3b_4 _50232_ (.A(net235),
    .B(_21305_),
    .C_N(_21342_),
    .X(_21344_));
 sky130_fd_sc_hd__and2_1 _50233_ (.A(_21343_),
    .B(_21344_),
    .X(_21345_));
 sky130_fd_sc_hd__nand2_2 _50234_ (.A(_21298_),
    .B(_21345_),
    .Y(_21346_));
 sky130_fd_sc_hd__or2_1 _50235_ (.A(_21298_),
    .B(_21345_),
    .X(_21347_));
 sky130_fd_sc_hd__and2_2 _50236_ (.A(_21346_),
    .B(_21347_),
    .X(_21348_));
 sky130_fd_sc_hd__xnor2_4 _50237_ (.A(_21259_),
    .B(_21348_),
    .Y(_21349_));
 sky130_fd_sc_hd__o21a_1 _50238_ (.A1(_20507_),
    .A2(_20510_),
    .B1(_21349_),
    .X(_21350_));
 sky130_fd_sc_hd__a211oi_1 _50239_ (.A1(_20508_),
    .A2(_20509_),
    .B1(_20507_),
    .C1(_21349_),
    .Y(_21351_));
 sky130_fd_sc_hd__nor2_1 _50240_ (.A(_21350_),
    .B(_21351_),
    .Y(_21352_));
 sky130_fd_sc_hd__xnor2_2 _50241_ (.A(_21201_),
    .B(_21352_),
    .Y(_21353_));
 sky130_fd_sc_hd__buf_2 _50242_ (.A(_19391_),
    .X(_21354_));
 sky130_fd_sc_hd__inv_2 _50243_ (.A(net374),
    .Y(_21355_));
 sky130_fd_sc_hd__inv_2 _50244_ (.A(\delay_line[18][6] ),
    .Y(_21356_));
 sky130_fd_sc_hd__buf_1 _50245_ (.A(\delay_line[18][3] ),
    .X(_21357_));
 sky130_fd_sc_hd__buf_1 _50246_ (.A(\delay_line[18][7] ),
    .X(_21358_));
 sky130_fd_sc_hd__and2_1 _50247_ (.A(_21357_),
    .B(_21358_),
    .X(_21359_));
 sky130_fd_sc_hd__nor2_1 _50248_ (.A(_21357_),
    .B(_21358_),
    .Y(_21360_));
 sky130_fd_sc_hd__o22ai_2 _50249_ (.A1(_21355_),
    .A2(_21356_),
    .B1(_21359_),
    .B2(_21360_),
    .Y(_21361_));
 sky130_fd_sc_hd__buf_2 _50250_ (.A(\delay_line[18][6] ),
    .X(_21362_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50251_ (.A(\delay_line[18][7] ),
    .X(_21363_));
 sky130_fd_sc_hd__nand2_1 _50252_ (.A(_21357_),
    .B(_21363_),
    .Y(_21364_));
 sky130_fd_sc_hd__nand4b_4 _50253_ (.A_N(_21360_),
    .B(_21362_),
    .C(_07514_),
    .D(_21364_),
    .Y(_21365_));
 sky130_fd_sc_hd__nand3_1 _50254_ (.A(_21361_),
    .B(_23852_),
    .C(_21365_),
    .Y(_21366_));
 sky130_fd_sc_hd__clkbuf_2 _50255_ (.A(_21366_),
    .X(_21367_));
 sky130_fd_sc_hd__a21o_1 _50256_ (.A1(_21365_),
    .A2(_21361_),
    .B1(_23852_),
    .X(_21368_));
 sky130_fd_sc_hd__a32o_1 _50257_ (.A1(_01677_),
    .A2(_21354_),
    .A3(_20543_),
    .B1(_21367_),
    .B2(_21368_),
    .X(_21369_));
 sky130_fd_sc_hd__nand4_2 _50258_ (.A(_21368_),
    .B(_20543_),
    .C(_19396_),
    .D(_21367_),
    .Y(_21370_));
 sky130_fd_sc_hd__and4_1 _50259_ (.A(_21369_),
    .B(_20544_),
    .C(_20541_),
    .D(_21370_),
    .X(_21371_));
 sky130_fd_sc_hd__a22oi_2 _50260_ (.A1(_20541_),
    .A2(_20544_),
    .B1(_21370_),
    .B2(_21369_),
    .Y(_21372_));
 sky130_fd_sc_hd__a22o_1 _50261_ (.A1(_20553_),
    .A2(_19401_),
    .B1(_20551_),
    .B2(_07371_),
    .X(_21373_));
 sky130_fd_sc_hd__nor2_1 _50262_ (.A(_20547_),
    .B(\delay_line[19][7] ),
    .Y(_21374_));
 sky130_fd_sc_hd__and2_1 _50263_ (.A(\delay_line[19][6] ),
    .B(net370),
    .X(_21375_));
 sky130_fd_sc_hd__nand2_2 _50264_ (.A(_19402_),
    .B(_20560_),
    .Y(_21376_));
 sky130_fd_sc_hd__o21ai_2 _50265_ (.A1(_21374_),
    .A2(_21375_),
    .B1(_21376_),
    .Y(_21377_));
 sky130_fd_sc_hd__inv_2 _50266_ (.A(net370),
    .Y(_21378_));
 sky130_fd_sc_hd__nand2_1 _50267_ (.A(_20548_),
    .B(_21378_),
    .Y(_21379_));
 sky130_fd_sc_hd__a21o_1 _50268_ (.A1(_21377_),
    .A2(_21379_),
    .B1(_07448_),
    .X(_21380_));
 sky130_fd_sc_hd__buf_1 _50269_ (.A(net370),
    .X(_21381_));
 sky130_fd_sc_hd__buf_2 _50270_ (.A(_21381_),
    .X(_21382_));
 sky130_fd_sc_hd__o211ai_1 _50271_ (.A1(_21382_),
    .A2(_21376_),
    .B1(_07448_),
    .C1(_21377_),
    .Y(_21383_));
 sky130_fd_sc_hd__nand3_2 _50272_ (.A(_21373_),
    .B(_21380_),
    .C(_21383_),
    .Y(_21384_));
 sky130_fd_sc_hd__a21oi_1 _50273_ (.A1(_21377_),
    .A2(_21379_),
    .B1(_07448_),
    .Y(_21385_));
 sky130_fd_sc_hd__and3_1 _50274_ (.A(_21377_),
    .B(_21379_),
    .C(_07393_),
    .X(_21386_));
 sky130_fd_sc_hd__o2bb2a_1 _50275_ (.A1_N(_07371_),
    .A2_N(_20552_),
    .B1(_20550_),
    .B2(_20561_),
    .X(_21387_));
 sky130_fd_sc_hd__o21ai_2 _50276_ (.A1(_21385_),
    .A2(_21386_),
    .B1(_21387_),
    .Y(_21388_));
 sky130_fd_sc_hd__a2bb2o_1 _50277_ (.A1_N(_01633_),
    .A2_N(_01655_),
    .B1(_21384_),
    .B2(_21388_),
    .X(_21389_));
 sky130_fd_sc_hd__nand3b_1 _50278_ (.A_N(_01710_),
    .B(_21384_),
    .C(_21388_),
    .Y(_21390_));
 sky130_fd_sc_hd__a21boi_1 _50279_ (.A1(_20558_),
    .A2(_23896_),
    .B1_N(_20563_),
    .Y(_21391_));
 sky130_fd_sc_hd__nand3_1 _50280_ (.A(_21389_),
    .B(_21390_),
    .C(_21391_),
    .Y(_21392_));
 sky130_fd_sc_hd__nand2_1 _50281_ (.A(_20563_),
    .B(_20564_),
    .Y(_21393_));
 sky130_fd_sc_hd__o211ai_2 _50282_ (.A1(_01633_),
    .A2(_01655_),
    .B1(_21384_),
    .C1(_21388_),
    .Y(_21394_));
 sky130_fd_sc_hd__a21o_1 _50283_ (.A1(_21384_),
    .A2(_21388_),
    .B1(_01710_),
    .X(_21395_));
 sky130_fd_sc_hd__nand3_2 _50284_ (.A(_21393_),
    .B(_21394_),
    .C(_21395_),
    .Y(_21396_));
 sky130_fd_sc_hd__nand4_2 _50285_ (.A(_20567_),
    .B(_20571_),
    .C(_21392_),
    .D(_21396_),
    .Y(_21397_));
 sky130_fd_sc_hd__nand4_1 _50286_ (.A(_19400_),
    .B(_19407_),
    .C(_19408_),
    .D(_18377_),
    .Y(_21398_));
 sky130_fd_sc_hd__nand2_1 _50287_ (.A(_20565_),
    .B(_20566_),
    .Y(_21399_));
 sky130_fd_sc_hd__o2bb2ai_1 _50288_ (.A1_N(_21392_),
    .A2_N(_21396_),
    .B1(_21398_),
    .B2(_21399_),
    .Y(_21400_));
 sky130_fd_sc_hd__nand4_1 _50289_ (.A(_21397_),
    .B(_21400_),
    .C(_20571_),
    .D(_20570_),
    .Y(_21401_));
 sky130_fd_sc_hd__inv_2 _50290_ (.A(_21401_),
    .Y(_21402_));
 sky130_fd_sc_hd__a22oi_2 _50291_ (.A1(_20571_),
    .A2(_20570_),
    .B1(_21397_),
    .B2(_21400_),
    .Y(_21403_));
 sky130_fd_sc_hd__o21ai_1 _50292_ (.A1(_21402_),
    .A2(_21403_),
    .B1(_20573_),
    .Y(_21404_));
 sky130_fd_sc_hd__or2_1 _50293_ (.A(_20573_),
    .B(_21403_),
    .X(_21405_));
 sky130_fd_sc_hd__or4bb_4 _50294_ (.A(_21371_),
    .B(_21372_),
    .C_N(_21404_),
    .D_N(_21405_),
    .X(_21406_));
 sky130_fd_sc_hd__inv_2 _50295_ (.A(_21406_),
    .Y(_21407_));
 sky130_fd_sc_hd__a2bb2oi_2 _50296_ (.A1_N(_21371_),
    .A2_N(_21372_),
    .B1(_21404_),
    .B2(_21405_),
    .Y(_21408_));
 sky130_fd_sc_hd__a2bb2o_1 _50297_ (.A1_N(_20521_),
    .A2_N(_20517_),
    .B1(_01600_),
    .B2(_20518_),
    .X(_21409_));
 sky130_fd_sc_hd__nor2_1 _50298_ (.A(_20514_),
    .B(\delay_line[21][7] ),
    .Y(_21410_));
 sky130_fd_sc_hd__and2_1 _50299_ (.A(_20514_),
    .B(\delay_line[21][7] ),
    .X(_21411_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50300_ (.A(\delay_line[21][5] ),
    .X(_21412_));
 sky130_fd_sc_hd__nand2_1 _50301_ (.A(_21412_),
    .B(_20514_),
    .Y(_21413_));
 sky130_fd_sc_hd__o21ai_2 _50302_ (.A1(_21410_),
    .A2(_21411_),
    .B1(_21413_),
    .Y(_21414_));
 sky130_fd_sc_hd__buf_1 _50303_ (.A(\delay_line[21][7] ),
    .X(_21415_));
 sky130_fd_sc_hd__or2_1 _50304_ (.A(_21415_),
    .B(_21413_),
    .X(_21416_));
 sky130_fd_sc_hd__a21o_1 _50305_ (.A1(_21414_),
    .A2(_21416_),
    .B1(_07305_),
    .X(_21417_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50306_ (.A(_21415_),
    .X(_21418_));
 sky130_fd_sc_hd__buf_1 _50307_ (.A(net361),
    .X(_21419_));
 sky130_fd_sc_hd__o211ai_1 _50308_ (.A1(_21418_),
    .A2(_21413_),
    .B1(_21419_),
    .C1(_21414_),
    .Y(_21420_));
 sky130_fd_sc_hd__nand3_1 _50309_ (.A(_21409_),
    .B(_21417_),
    .C(_21420_),
    .Y(_21421_));
 sky130_fd_sc_hd__buf_2 _50310_ (.A(_21421_),
    .X(_21422_));
 sky130_fd_sc_hd__clkbuf_2 _50311_ (.A(_20521_),
    .X(_21423_));
 sky130_fd_sc_hd__a21oi_1 _50312_ (.A1(_21414_),
    .A2(_21416_),
    .B1(_21419_),
    .Y(_21424_));
 sky130_fd_sc_hd__and3_1 _50313_ (.A(_21414_),
    .B(_21416_),
    .C(_07305_),
    .X(_21425_));
 sky130_fd_sc_hd__o221ai_4 _50314_ (.A1(_21423_),
    .A2(_20517_),
    .B1(_21424_),
    .B2(_21425_),
    .C1(_20522_),
    .Y(_21426_));
 sky130_fd_sc_hd__a2bb2o_1 _50315_ (.A1_N(_01589_),
    .A2_N(_01611_),
    .B1(_21422_),
    .B2(_21426_),
    .X(_21427_));
 sky130_fd_sc_hd__nand3_1 _50316_ (.A(_21426_),
    .B(_01622_),
    .C(_21422_),
    .Y(_21428_));
 sky130_fd_sc_hd__a21boi_1 _50317_ (.A1(_20524_),
    .A2(_07338_),
    .B1_N(_20525_),
    .Y(_21429_));
 sky130_fd_sc_hd__nand3_2 _50318_ (.A(_21427_),
    .B(_21428_),
    .C(_21429_),
    .Y(_21430_));
 sky130_fd_sc_hd__nand2_1 _50319_ (.A(_20525_),
    .B(_20526_),
    .Y(_21431_));
 sky130_fd_sc_hd__o211ai_4 _50320_ (.A1(_01589_),
    .A2(_01611_),
    .B1(_21422_),
    .C1(_21426_),
    .Y(_21432_));
 sky130_fd_sc_hd__nand2_1 _50321_ (.A(_21421_),
    .B(_21426_),
    .Y(_21433_));
 sky130_fd_sc_hd__nand2_1 _50322_ (.A(_21433_),
    .B(_01622_),
    .Y(_21434_));
 sky130_fd_sc_hd__nand3_4 _50323_ (.A(_21431_),
    .B(_21432_),
    .C(_21434_),
    .Y(_21435_));
 sky130_fd_sc_hd__nand4_4 _50324_ (.A(_20529_),
    .B(_20534_),
    .C(_21430_),
    .D(_21435_),
    .Y(_21436_));
 sky130_fd_sc_hd__nand2_1 _50325_ (.A(_20526_),
    .B(_20527_),
    .Y(_21437_));
 sky130_fd_sc_hd__o2bb2ai_1 _50326_ (.A1_N(_21430_),
    .A2_N(_21435_),
    .B1(_19424_),
    .B2(_21437_),
    .Y(_21438_));
 sky130_fd_sc_hd__nand4_1 _50327_ (.A(_21436_),
    .B(_21438_),
    .C(_20530_),
    .D(_20534_),
    .Y(_21439_));
 sky130_fd_sc_hd__a32o_1 _50328_ (.A1(_20530_),
    .A2(_20526_),
    .A3(_20527_),
    .B1(_21436_),
    .B2(_21438_),
    .X(_21440_));
 sky130_fd_sc_hd__nand2_1 _50329_ (.A(_21439_),
    .B(_21440_),
    .Y(_21441_));
 sky130_fd_sc_hd__xnor2_1 _50330_ (.A(_20538_),
    .B(_21441_),
    .Y(_21442_));
 sky130_fd_sc_hd__or3b_4 _50331_ (.A(_21407_),
    .B(_21408_),
    .C_N(_21442_),
    .X(_21443_));
 sky130_fd_sc_hd__o21bai_1 _50332_ (.A1(_21407_),
    .A2(_21408_),
    .B1_N(_21442_),
    .Y(_21444_));
 sky130_fd_sc_hd__and2_1 _50333_ (.A(_21443_),
    .B(_21444_),
    .X(_21445_));
 sky130_fd_sc_hd__buf_1 _50334_ (.A(_20615_),
    .X(_21446_));
 sky130_fd_sc_hd__o211a_1 _50335_ (.A1(_19468_),
    .A2(_18420_),
    .B1(_19465_),
    .C1(_19466_),
    .X(_21447_));
 sky130_fd_sc_hd__nand3_2 _50336_ (.A(_20614_),
    .B(_21447_),
    .C(_20613_),
    .Y(_21448_));
 sky130_fd_sc_hd__nand2_1 _50337_ (.A(_20605_),
    .B(_20611_),
    .Y(_21449_));
 sky130_fd_sc_hd__and2_1 _50338_ (.A(\delay_line[15][6] ),
    .B(\delay_line[15][8] ),
    .X(_21450_));
 sky130_fd_sc_hd__clkbuf_2 _50339_ (.A(_21450_),
    .X(_21451_));
 sky130_fd_sc_hd__buf_2 _50340_ (.A(\delay_line[15][8] ),
    .X(_21452_));
 sky130_fd_sc_hd__o211ai_4 _50341_ (.A1(_19461_),
    .A2(_21452_),
    .B1(_20600_),
    .C1(_18416_),
    .Y(_21453_));
 sky130_fd_sc_hd__buf_2 _50342_ (.A(_20598_),
    .X(_21454_));
 sky130_fd_sc_hd__nor2_1 _50343_ (.A(_19461_),
    .B(_21452_),
    .Y(_21455_));
 sky130_fd_sc_hd__o22ai_4 _50344_ (.A1(_21454_),
    .A2(_20596_),
    .B1(_21450_),
    .B2(_21455_),
    .Y(_21456_));
 sky130_fd_sc_hd__o211ai_1 _50345_ (.A1(_21451_),
    .A2(_21453_),
    .B1(_07096_),
    .C1(_21456_),
    .Y(_21457_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50346_ (.A(_19461_),
    .X(_21458_));
 sky130_fd_sc_hd__clkbuf_2 _50347_ (.A(_21452_),
    .X(_21459_));
 sky130_fd_sc_hd__a21o_1 _50348_ (.A1(_21458_),
    .A2(_21459_),
    .B1(_21453_),
    .X(_21460_));
 sky130_fd_sc_hd__a21o_1 _50349_ (.A1(_21460_),
    .A2(_21456_),
    .B1(_16777_),
    .X(_21461_));
 sky130_fd_sc_hd__nand3_2 _50350_ (.A(_21449_),
    .B(_21457_),
    .C(_21461_),
    .Y(_21462_));
 sky130_fd_sc_hd__o211a_1 _50351_ (.A1(_21451_),
    .A2(_21453_),
    .B1(_16777_),
    .C1(_21456_),
    .X(_21463_));
 sky130_fd_sc_hd__a21oi_1 _50352_ (.A1(_21460_),
    .A2(_21456_),
    .B1(_16777_),
    .Y(_21464_));
 sky130_fd_sc_hd__a21boi_1 _50353_ (.A1(_01798_),
    .A2(_20602_),
    .B1_N(_20605_),
    .Y(_21465_));
 sky130_fd_sc_hd__o21ai_2 _50354_ (.A1(_21463_),
    .A2(_21464_),
    .B1(_21465_),
    .Y(_21466_));
 sky130_fd_sc_hd__and2_1 _50355_ (.A(_07063_),
    .B(_22391_),
    .X(_21467_));
 sky130_fd_sc_hd__nor2_1 _50356_ (.A(_22391_),
    .B(_07118_),
    .Y(_21468_));
 sky130_fd_sc_hd__or2_1 _50357_ (.A(_21467_),
    .B(_21468_),
    .X(_21469_));
 sky130_fd_sc_hd__a21oi_1 _50358_ (.A1(_21462_),
    .A2(_21466_),
    .B1(_21469_),
    .Y(_21470_));
 sky130_fd_sc_hd__and3_1 _50359_ (.A(_21462_),
    .B(_21466_),
    .C(_21469_),
    .X(_21471_));
 sky130_fd_sc_hd__o211ai_1 _50360_ (.A1(_21470_),
    .A2(_21471_),
    .B1(_20612_),
    .C1(_20613_),
    .Y(_21472_));
 sky130_fd_sc_hd__a21o_1 _50361_ (.A1(_21462_),
    .A2(_21466_),
    .B1(_21469_),
    .X(_21473_));
 sky130_fd_sc_hd__o211ai_4 _50362_ (.A1(_21467_),
    .A2(_21468_),
    .B1(_21462_),
    .C1(_21466_),
    .Y(_21474_));
 sky130_fd_sc_hd__nand2_1 _50363_ (.A(_20612_),
    .B(_20613_),
    .Y(_21475_));
 sky130_fd_sc_hd__nand3_4 _50364_ (.A(_21473_),
    .B(_21474_),
    .C(_21475_),
    .Y(_21476_));
 sky130_fd_sc_hd__nand3b_2 _50365_ (.A_N(_21448_),
    .B(_21472_),
    .C(_21476_),
    .Y(_21477_));
 sky130_fd_sc_hd__a21oi_2 _50366_ (.A1(_21473_),
    .A2(_21474_),
    .B1(_21475_),
    .Y(_21478_));
 sky130_fd_sc_hd__a211oi_2 _50367_ (.A1(_20612_),
    .A2(_20613_),
    .B1(_21470_),
    .C1(_21471_),
    .Y(_21479_));
 sky130_fd_sc_hd__o21ai_1 _50368_ (.A1(_21478_),
    .A2(_21479_),
    .B1(_21448_),
    .Y(_21480_));
 sky130_fd_sc_hd__a2bb2o_2 _50369_ (.A1_N(_20595_),
    .A2_N(_21446_),
    .B1(_21477_),
    .B2(_21480_),
    .X(_21481_));
 sky130_fd_sc_hd__o22a_1 _50370_ (.A1(_19470_),
    .A2(_21446_),
    .B1(_21478_),
    .B2(_21479_),
    .X(_21482_));
 sky130_fd_sc_hd__or4_2 _50371_ (.A(_18431_),
    .B(_19472_),
    .C(_21446_),
    .D(_21482_),
    .X(_21483_));
 sky130_fd_sc_hd__a21oi_2 _50372_ (.A1(_21481_),
    .A2(_21483_),
    .B1(_20619_),
    .Y(_21484_));
 sky130_fd_sc_hd__a2bb2oi_1 _50373_ (.A1_N(_20595_),
    .A2_N(_21446_),
    .B1(_21477_),
    .B2(_21480_),
    .Y(_21485_));
 sky130_fd_sc_hd__and2_1 _50374_ (.A(_20618_),
    .B(_20616_),
    .X(_21486_));
 sky130_fd_sc_hd__or4b_2 _50375_ (.A(_18432_),
    .B(_19472_),
    .C(_21485_),
    .D_N(_21486_),
    .X(_21487_));
 sky130_fd_sc_hd__inv_2 _50376_ (.A(_21487_),
    .Y(_21488_));
 sky130_fd_sc_hd__o211ai_4 _50377_ (.A1(_19449_),
    .A2(_20583_),
    .B1(_20588_),
    .C1(_20590_),
    .Y(_21489_));
 sky130_fd_sc_hd__nand2_1 _50378_ (.A(_01765_),
    .B(_07173_),
    .Y(_21490_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50379_ (.A(net392),
    .X(_21491_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50380_ (.A(\delay_line[14][7] ),
    .X(_21492_));
 sky130_fd_sc_hd__o21ai_1 _50381_ (.A1(\delay_line[14][3] ),
    .A2(_20584_),
    .B1(_21492_),
    .Y(_21493_));
 sky130_fd_sc_hd__a21oi_1 _50382_ (.A1(_21491_),
    .A2(_20584_),
    .B1(_21493_),
    .Y(_21494_));
 sky130_fd_sc_hd__and2_1 _50383_ (.A(_16821_),
    .B(_20584_),
    .X(_21495_));
 sky130_fd_sc_hd__nor2_1 _50384_ (.A(_21491_),
    .B(_07173_),
    .Y(_21496_));
 sky130_fd_sc_hd__buf_1 _50385_ (.A(_21492_),
    .X(_21497_));
 sky130_fd_sc_hd__o21ba_1 _50386_ (.A1(_21495_),
    .A2(_21496_),
    .B1_N(_21497_),
    .X(_21498_));
 sky130_fd_sc_hd__a211o_1 _50387_ (.A1(_21490_),
    .A2(_20588_),
    .B1(_21494_),
    .C1(_21498_),
    .X(_21499_));
 sky130_fd_sc_hd__inv_2 _50388_ (.A(_21499_),
    .Y(_21500_));
 sky130_fd_sc_hd__o211a_2 _50389_ (.A1(_21494_),
    .A2(_21498_),
    .B1(_21490_),
    .C1(_20588_),
    .X(_21501_));
 sky130_fd_sc_hd__nor2_1 _50390_ (.A(_21500_),
    .B(_21501_),
    .Y(_21502_));
 sky130_fd_sc_hd__o211a_1 _50391_ (.A1(_19455_),
    .A2(_20592_),
    .B1(_21489_),
    .C1(_21502_),
    .X(_21503_));
 sky130_fd_sc_hd__o22a_1 _50392_ (.A1(_20591_),
    .A2(_20593_),
    .B1(_21500_),
    .B2(_21501_),
    .X(_21504_));
 sky130_fd_sc_hd__nor2_2 _50393_ (.A(_21503_),
    .B(_21504_),
    .Y(_21505_));
 sky130_fd_sc_hd__o21ai_2 _50394_ (.A1(_21484_),
    .A2(_21488_),
    .B1(_21505_),
    .Y(_21506_));
 sky130_fd_sc_hd__a311o_1 _50395_ (.A1(_20617_),
    .A2(_21481_),
    .A3(_21486_),
    .B1(_21505_),
    .C1(_21484_),
    .X(_21507_));
 sky130_fd_sc_hd__nand2_1 _50396_ (.A(_19445_),
    .B(_20639_),
    .Y(_21508_));
 sky130_fd_sc_hd__buf_1 _50397_ (.A(_07206_),
    .X(_21509_));
 sky130_fd_sc_hd__o21a_1 _50398_ (.A1(_16590_),
    .A2(_21509_),
    .B1(_01864_),
    .X(_21510_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50399_ (.A(_21510_),
    .X(_21511_));
 sky130_fd_sc_hd__a21oi_1 _50400_ (.A1(_16590_),
    .A2(_21509_),
    .B1(_01875_),
    .Y(_21512_));
 sky130_fd_sc_hd__and2_2 _50401_ (.A(\delay_line[16][3] ),
    .B(\delay_line[16][4] ),
    .X(_21513_));
 sky130_fd_sc_hd__clkbuf_2 _50402_ (.A(\delay_line[16][4] ),
    .X(_21514_));
 sky130_fd_sc_hd__o21ai_4 _50403_ (.A1(_16656_),
    .A2(_21514_),
    .B1(_07206_),
    .Y(_21515_));
 sky130_fd_sc_hd__clkbuf_2 _50404_ (.A(\delay_line[16][7] ),
    .X(_21516_));
 sky130_fd_sc_hd__clkbuf_2 _50405_ (.A(_21516_),
    .X(_21517_));
 sky130_fd_sc_hd__clkbuf_2 _50406_ (.A(_21517_),
    .X(_21518_));
 sky130_fd_sc_hd__nor2_1 _50407_ (.A(_16656_),
    .B(_21514_),
    .Y(_21519_));
 sky130_fd_sc_hd__o21ai_2 _50408_ (.A1(_21513_),
    .A2(_21519_),
    .B1(_07217_),
    .Y(_21520_));
 sky130_fd_sc_hd__o211ai_2 _50409_ (.A1(_21513_),
    .A2(_21515_),
    .B1(_21518_),
    .C1(_21520_),
    .Y(_21521_));
 sky130_fd_sc_hd__a21o_1 _50410_ (.A1(_16590_),
    .A2(_18399_),
    .B1(_21515_),
    .X(_21522_));
 sky130_fd_sc_hd__a21o_1 _50411_ (.A1(_21520_),
    .A2(_21522_),
    .B1(_21517_),
    .X(_21523_));
 sky130_fd_sc_hd__nand3_1 _50412_ (.A(_20632_),
    .B(_21521_),
    .C(_21523_),
    .Y(_21524_));
 sky130_fd_sc_hd__and3_1 _50413_ (.A(_21520_),
    .B(_21522_),
    .C(_21517_),
    .X(_21525_));
 sky130_fd_sc_hd__a21oi_1 _50414_ (.A1(_21520_),
    .A2(_21522_),
    .B1(_21518_),
    .Y(_21526_));
 sky130_fd_sc_hd__o21bai_1 _50415_ (.A1(_21525_),
    .A2(_21526_),
    .B1_N(_20631_),
    .Y(_21527_));
 sky130_fd_sc_hd__o211ai_2 _50416_ (.A1(_21511_),
    .A2(_21512_),
    .B1(_21524_),
    .C1(_21527_),
    .Y(_21528_));
 sky130_fd_sc_hd__o21ai_1 _50417_ (.A1(_21525_),
    .A2(_21526_),
    .B1(_20632_),
    .Y(_21529_));
 sky130_fd_sc_hd__nor2_1 _50418_ (.A(_21510_),
    .B(_21512_),
    .Y(_21530_));
 sky130_fd_sc_hd__nand3b_1 _50419_ (.A_N(_20631_),
    .B(_21521_),
    .C(_21523_),
    .Y(_21531_));
 sky130_fd_sc_hd__nand3_2 _50420_ (.A(_21529_),
    .B(_21530_),
    .C(_21531_),
    .Y(_21532_));
 sky130_fd_sc_hd__nand3_1 _50421_ (.A(_19439_),
    .B(_20632_),
    .C(_20635_),
    .Y(_21533_));
 sky130_fd_sc_hd__o21ai_1 _50422_ (.A1(_20625_),
    .A2(_20637_),
    .B1(_21533_),
    .Y(_21534_));
 sky130_fd_sc_hd__a21oi_1 _50423_ (.A1(_21528_),
    .A2(_21532_),
    .B1(_21534_),
    .Y(_21535_));
 sky130_fd_sc_hd__clkbuf_2 _50424_ (.A(_21509_),
    .X(_21536_));
 sky130_fd_sc_hd__o21a_1 _50425_ (.A1(_01886_),
    .A2(_21536_),
    .B1(_24138_),
    .X(_21537_));
 sky130_fd_sc_hd__nand3_2 _50426_ (.A(_21528_),
    .B(_21532_),
    .C(_21534_),
    .Y(_21538_));
 sky130_fd_sc_hd__nand3b_2 _50427_ (.A_N(_21535_),
    .B(_21537_),
    .C(_21538_),
    .Y(_21539_));
 sky130_fd_sc_hd__and3_1 _50428_ (.A(_21528_),
    .B(_21532_),
    .C(_21534_),
    .X(_21540_));
 sky130_fd_sc_hd__o22ai_2 _50429_ (.A1(_19437_),
    .A2(_16645_),
    .B1(_21535_),
    .B2(_21540_),
    .Y(_21541_));
 sky130_fd_sc_hd__nand4_2 _50430_ (.A(_21539_),
    .B(_21541_),
    .C(_19446_),
    .D(_20639_),
    .Y(_21542_));
 sky130_fd_sc_hd__inv_2 _50431_ (.A(_21542_),
    .Y(_21543_));
 sky130_fd_sc_hd__a22oi_2 _50432_ (.A1(_19446_),
    .A2(_20639_),
    .B1(_21539_),
    .B2(_21541_),
    .Y(_21544_));
 sky130_fd_sc_hd__or2_1 _50433_ (.A(_21543_),
    .B(_21544_),
    .X(_21545_));
 sky130_fd_sc_hd__xor2_1 _50434_ (.A(_21508_),
    .B(_21545_),
    .X(_21546_));
 sky130_fd_sc_hd__and3_1 _50435_ (.A(_21506_),
    .B(_21507_),
    .C(_21546_),
    .X(_21547_));
 sky130_fd_sc_hd__a21oi_1 _50436_ (.A1(_21506_),
    .A2(_21507_),
    .B1(_21546_),
    .Y(_21548_));
 sky130_fd_sc_hd__o211a_1 _50437_ (.A1(_21547_),
    .A2(_21548_),
    .B1(_20621_),
    .C1(_20643_),
    .X(_21549_));
 sky130_fd_sc_hd__a211o_4 _50438_ (.A1(_20621_),
    .A2(_20643_),
    .B1(_21547_),
    .C1(_21548_),
    .X(_21550_));
 sky130_fd_sc_hd__and2b_2 _50439_ (.A_N(_21549_),
    .B(_21550_),
    .X(_21551_));
 sky130_fd_sc_hd__xor2_1 _50440_ (.A(_21445_),
    .B(_21551_),
    .X(_21552_));
 sky130_fd_sc_hd__a211oi_1 _50441_ (.A1(_20582_),
    .A2(_20648_),
    .B1(_21552_),
    .C1(_20647_),
    .Y(_21553_));
 sky130_fd_sc_hd__o21a_2 _50442_ (.A1(_20647_),
    .A2(_20649_),
    .B1(_21552_),
    .X(_21554_));
 sky130_fd_sc_hd__nor2_2 _50443_ (.A(_21553_),
    .B(_21554_),
    .Y(_21555_));
 sky130_fd_sc_hd__and4bb_1 _50444_ (.A_N(_20453_),
    .B_N(_20455_),
    .C(_20479_),
    .D(_20477_),
    .X(_21556_));
 sky130_fd_sc_hd__nor2_1 _50445_ (.A(_21556_),
    .B(_20504_),
    .Y(_21557_));
 sky130_fd_sc_hd__a21oi_1 _50446_ (.A1(_20484_),
    .A2(_20485_),
    .B1(_19491_),
    .Y(_21558_));
 sky130_fd_sc_hd__a21oi_1 _50447_ (.A1(_17139_),
    .A2(_20486_),
    .B1(_21558_),
    .Y(_21559_));
 sky130_fd_sc_hd__and2_1 _50448_ (.A(\delay_line[25][6] ),
    .B(\delay_line[25][8] ),
    .X(_21560_));
 sky130_fd_sc_hd__clkbuf_2 _50449_ (.A(_21560_),
    .X(_21561_));
 sky130_fd_sc_hd__clkbuf_2 _50450_ (.A(\delay_line[25][8] ),
    .X(_21562_));
 sky130_fd_sc_hd__clkbuf_2 _50451_ (.A(_21562_),
    .X(_21563_));
 sky130_fd_sc_hd__o211ai_2 _50452_ (.A1(\delay_line[25][6] ),
    .A2(_21563_),
    .B1(_20483_),
    .C1(_18323_),
    .Y(_21564_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50453_ (.A(_20483_),
    .X(_21565_));
 sky130_fd_sc_hd__nor2_1 _50454_ (.A(_19488_),
    .B(_21563_),
    .Y(_21566_));
 sky130_fd_sc_hd__o2bb2ai_2 _50455_ (.A1_N(_18323_),
    .A2_N(_21565_),
    .B1(_21561_),
    .B2(_21566_),
    .Y(_21567_));
 sky130_fd_sc_hd__o211ai_1 _50456_ (.A1(_21561_),
    .A2(_21564_),
    .B1(_06788_),
    .C1(_21567_),
    .Y(_21568_));
 sky130_fd_sc_hd__buf_1 _50457_ (.A(_19488_),
    .X(_21569_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50458_ (.A(_21562_),
    .X(_21570_));
 sky130_fd_sc_hd__a21o_1 _50459_ (.A1(_21569_),
    .A2(_21570_),
    .B1(_21564_),
    .X(_21571_));
 sky130_fd_sc_hd__a21o_1 _50460_ (.A1(_21571_),
    .A2(_21567_),
    .B1(_17171_),
    .X(_21572_));
 sky130_fd_sc_hd__nand3b_2 _50461_ (.A_N(_21559_),
    .B(_21568_),
    .C(_21572_),
    .Y(_21573_));
 sky130_fd_sc_hd__o211a_1 _50462_ (.A1(_21561_),
    .A2(_21564_),
    .B1(_17171_),
    .C1(_21567_),
    .X(_21574_));
 sky130_fd_sc_hd__a21oi_1 _50463_ (.A1(_21571_),
    .A2(_21567_),
    .B1(_06788_),
    .Y(_21575_));
 sky130_fd_sc_hd__o21ai_2 _50464_ (.A1(_21574_),
    .A2(_21575_),
    .B1(_21559_),
    .Y(_21576_));
 sky130_fd_sc_hd__nand2_1 _50465_ (.A(_22358_),
    .B(_23731_),
    .Y(_21577_));
 sky130_fd_sc_hd__or2_1 _50466_ (.A(\delay_line[25][0] ),
    .B(\delay_line[25][1] ),
    .X(_21578_));
 sky130_fd_sc_hd__and2_1 _50467_ (.A(_21577_),
    .B(_21578_),
    .X(_21579_));
 sky130_fd_sc_hd__a21oi_1 _50468_ (.A1(_21573_),
    .A2(_21576_),
    .B1(_21579_),
    .Y(_21580_));
 sky130_fd_sc_hd__and3_1 _50469_ (.A(_21573_),
    .B(_21576_),
    .C(_21579_),
    .X(_21581_));
 sky130_fd_sc_hd__a21boi_1 _50470_ (.A1(_22369_),
    .A2(_20493_),
    .B1_N(_20491_),
    .Y(_21582_));
 sky130_fd_sc_hd__o21a_1 _50471_ (.A1(_21580_),
    .A2(_21581_),
    .B1(_21582_),
    .X(_21583_));
 sky130_fd_sc_hd__a211oi_1 _50472_ (.A1(_20491_),
    .A2(_20494_),
    .B1(_21580_),
    .C1(_21581_),
    .Y(_21584_));
 sky130_fd_sc_hd__o22ai_2 _50473_ (.A1(_19496_),
    .A2(_20498_),
    .B1(_21583_),
    .B2(_21584_),
    .Y(_21585_));
 sky130_fd_sc_hd__nand3_1 _50474_ (.A(_20495_),
    .B(_20481_),
    .C(_20494_),
    .Y(_21586_));
 sky130_fd_sc_hd__o21ai_1 _50475_ (.A1(_21580_),
    .A2(_21581_),
    .B1(_21582_),
    .Y(_21587_));
 sky130_fd_sc_hd__a21o_1 _50476_ (.A1(_21573_),
    .A2(_21576_),
    .B1(_21579_),
    .X(_21588_));
 sky130_fd_sc_hd__nand3_1 _50477_ (.A(_21573_),
    .B(_21576_),
    .C(_21579_),
    .Y(_21589_));
 sky130_fd_sc_hd__nand2_1 _50478_ (.A(_20491_),
    .B(_20494_),
    .Y(_21590_));
 sky130_fd_sc_hd__nand3_2 _50479_ (.A(_21588_),
    .B(_21589_),
    .C(_21590_),
    .Y(_21591_));
 sky130_fd_sc_hd__nand3b_2 _50480_ (.A_N(_21586_),
    .B(_21587_),
    .C(_21591_),
    .Y(_21592_));
 sky130_fd_sc_hd__and4_1 _50481_ (.A(_21585_),
    .B(_20496_),
    .C(_21592_),
    .D(_20482_),
    .X(_21593_));
 sky130_fd_sc_hd__or3b_1 _50482_ (.A(_20481_),
    .B(_18332_),
    .C_N(_19495_),
    .X(_21594_));
 sky130_fd_sc_hd__a2bb2oi_2 _50483_ (.A1_N(_20498_),
    .A2_N(_21594_),
    .B1(_21592_),
    .B2(_21585_),
    .Y(_21595_));
 sky130_fd_sc_hd__o21a_1 _50484_ (.A1(_21593_),
    .A2(_21595_),
    .B1(_20502_),
    .X(_21596_));
 sky130_fd_sc_hd__nor2_2 _50485_ (.A(_20502_),
    .B(_21595_),
    .Y(_21597_));
 sky130_fd_sc_hd__nor2_1 _50486_ (.A(net354),
    .B(net352),
    .Y(_21598_));
 sky130_fd_sc_hd__inv_2 _50487_ (.A(\delay_line[22][6] ),
    .Y(_21599_));
 sky130_fd_sc_hd__buf_1 _50488_ (.A(\delay_line[22][2] ),
    .X(_21600_));
 sky130_fd_sc_hd__nand2_1 _50489_ (.A(net354),
    .B(net352),
    .Y(_21601_));
 sky130_fd_sc_hd__or4bb_2 _50490_ (.A(_21598_),
    .B(_21599_),
    .C_N(_21600_),
    .D_N(_21601_),
    .X(_21602_));
 sky130_fd_sc_hd__and2_1 _50491_ (.A(net354),
    .B(net352),
    .X(_21603_));
 sky130_fd_sc_hd__o2bb2ai_1 _50492_ (.A1_N(_06865_),
    .A2_N(_20449_),
    .B1(_21603_),
    .B2(_21598_),
    .Y(_21604_));
 sky130_fd_sc_hd__a21o_1 _50493_ (.A1(_21602_),
    .A2(_21604_),
    .B1(_23666_),
    .X(_21605_));
 sky130_fd_sc_hd__nand3_1 _50494_ (.A(_21602_),
    .B(_21604_),
    .C(_23666_),
    .Y(_21606_));
 sky130_fd_sc_hd__nand4_1 _50495_ (.A(_21605_),
    .B(_20451_),
    .C(_19504_),
    .D(_21606_),
    .Y(_21607_));
 sky130_fd_sc_hd__a32o_1 _50496_ (.A1(_01413_),
    .A2(_19502_),
    .A3(_20451_),
    .B1(_21606_),
    .B2(_21605_),
    .X(_21608_));
 sky130_fd_sc_hd__a22oi_1 _50497_ (.A1(_19507_),
    .A2(_20452_),
    .B1(_21607_),
    .B2(_21608_),
    .Y(_21609_));
 sky130_fd_sc_hd__and4_1 _50498_ (.A(_21608_),
    .B(_20452_),
    .C(_19506_),
    .D(_21607_),
    .X(_21610_));
 sky130_fd_sc_hd__and2_1 _50499_ (.A(_17018_),
    .B(_06898_),
    .X(_21611_));
 sky130_fd_sc_hd__o21ai_1 _50500_ (.A1(_17018_),
    .A2(_06909_),
    .B1(_01435_),
    .Y(_21612_));
 sky130_fd_sc_hd__o21ai_1 _50501_ (.A1(_01446_),
    .A2(_21611_),
    .B1(_21612_),
    .Y(_21613_));
 sky130_fd_sc_hd__nand2_1 _50502_ (.A(_20459_),
    .B(_20462_),
    .Y(_21614_));
 sky130_fd_sc_hd__and2_2 _50503_ (.A(\delay_line[24][3] ),
    .B(net343),
    .X(_21615_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50504_ (.A(net343),
    .X(_21616_));
 sky130_fd_sc_hd__o21ai_1 _50505_ (.A1(_20458_),
    .A2(_21616_),
    .B1(_06898_),
    .Y(_21617_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50506_ (.A(_21617_),
    .X(_21618_));
 sky130_fd_sc_hd__clkbuf_2 _50507_ (.A(\delay_line[24][7] ),
    .X(_21619_));
 sky130_fd_sc_hd__clkbuf_2 _50508_ (.A(_21619_),
    .X(_21620_));
 sky130_fd_sc_hd__nor2_1 _50509_ (.A(\delay_line[24][3] ),
    .B(_21616_),
    .Y(_21621_));
 sky130_fd_sc_hd__o21bai_2 _50510_ (.A1(_21615_),
    .A2(_21621_),
    .B1_N(_06898_),
    .Y(_21622_));
 sky130_fd_sc_hd__o211ai_2 _50511_ (.A1(_21615_),
    .A2(_21618_),
    .B1(_21620_),
    .C1(_21622_),
    .Y(_21623_));
 sky130_fd_sc_hd__a21o_1 _50512_ (.A1(_17007_),
    .A2(_18309_),
    .B1(_21617_),
    .X(_21624_));
 sky130_fd_sc_hd__a21o_1 _50513_ (.A1(_21624_),
    .A2(_21622_),
    .B1(_21620_),
    .X(_21625_));
 sky130_fd_sc_hd__o211ai_1 _50514_ (.A1(_20467_),
    .A2(_21614_),
    .B1(_21623_),
    .C1(_21625_),
    .Y(_21626_));
 sky130_fd_sc_hd__o211a_1 _50515_ (.A1(_21615_),
    .A2(_21617_),
    .B1(_21620_),
    .C1(_21622_),
    .X(_21627_));
 sky130_fd_sc_hd__clkbuf_2 _50516_ (.A(_21620_),
    .X(_21628_));
 sky130_fd_sc_hd__a21oi_1 _50517_ (.A1(_21624_),
    .A2(_21622_),
    .B1(_21628_),
    .Y(_21629_));
 sky130_fd_sc_hd__o21bai_1 _50518_ (.A1(_21627_),
    .A2(_21629_),
    .B1_N(_20466_),
    .Y(_21630_));
 sky130_fd_sc_hd__nand3_1 _50519_ (.A(_21613_),
    .B(_21626_),
    .C(_21630_),
    .Y(_21631_));
 sky130_fd_sc_hd__o21ai_1 _50520_ (.A1(_21627_),
    .A2(_21629_),
    .B1(_20466_),
    .Y(_21632_));
 sky130_fd_sc_hd__o21a_1 _50521_ (.A1(_01435_),
    .A2(_21611_),
    .B1(_21612_),
    .X(_21633_));
 sky130_fd_sc_hd__nand3b_1 _50522_ (.A_N(_20465_),
    .B(_21623_),
    .C(_21625_),
    .Y(_21634_));
 sky130_fd_sc_hd__nand3_1 _50523_ (.A(_21632_),
    .B(_21633_),
    .C(_21634_),
    .Y(_21635_));
 sky130_fd_sc_hd__nand3_1 _50524_ (.A(_19517_),
    .B(_20466_),
    .C(_20470_),
    .Y(_21636_));
 sky130_fd_sc_hd__o21ai_2 _50525_ (.A1(_20457_),
    .A2(_20472_),
    .B1(_21636_),
    .Y(_21637_));
 sky130_fd_sc_hd__nand3_1 _50526_ (.A(_21631_),
    .B(_21635_),
    .C(_21637_),
    .Y(_21638_));
 sky130_fd_sc_hd__a21o_1 _50527_ (.A1(_21631_),
    .A2(_21635_),
    .B1(_21637_),
    .X(_21639_));
 sky130_fd_sc_hd__o2111ai_4 _50528_ (.A1(_01446_),
    .A2(_06931_),
    .B1(_23687_),
    .C1(_21638_),
    .D1(_21639_),
    .Y(_21640_));
 sky130_fd_sc_hd__a21oi_1 _50529_ (.A1(_21631_),
    .A2(_21635_),
    .B1(_21637_),
    .Y(_21641_));
 sky130_fd_sc_hd__and3_1 _50530_ (.A(_21631_),
    .B(_21635_),
    .C(_21637_),
    .X(_21642_));
 sky130_fd_sc_hd__o22ai_4 _50531_ (.A1(_19514_),
    .A2(_18305_),
    .B1(_21641_),
    .B2(_21642_),
    .Y(_21643_));
 sky130_fd_sc_hd__a22oi_2 _50532_ (.A1(_20456_),
    .A2(_20474_),
    .B1(_21640_),
    .B2(_21643_),
    .Y(_21644_));
 sky130_fd_sc_hd__xor2_1 _50533_ (.A(_20457_),
    .B(_20473_),
    .X(_21645_));
 sky130_fd_sc_hd__and4_1 _50534_ (.A(_21643_),
    .B(_20456_),
    .C(_21640_),
    .D(_20475_),
    .X(_21646_));
 sky130_fd_sc_hd__or4_2 _50535_ (.A(_19527_),
    .B(_21644_),
    .C(_21645_),
    .D(_21646_),
    .X(_21647_));
 sky130_fd_sc_hd__a2bb2o_1 _50536_ (.A1_N(_21646_),
    .A2_N(_21644_),
    .B1(_19524_),
    .B2(_20475_),
    .X(_21648_));
 sky130_fd_sc_hd__and4bb_1 _50537_ (.A_N(_21609_),
    .B_N(_21610_),
    .C(_21647_),
    .D(_21648_),
    .X(_21649_));
 sky130_fd_sc_hd__a2bb2oi_1 _50538_ (.A1_N(_21609_),
    .A2_N(_21610_),
    .B1(_21647_),
    .B2(_21648_),
    .Y(_21650_));
 sky130_fd_sc_hd__nor4_1 _50539_ (.A(_21596_),
    .B(_21597_),
    .C(_21649_),
    .D(_21650_),
    .Y(_21651_));
 sky130_fd_sc_hd__o22a_1 _50540_ (.A1(_21596_),
    .A2(_21597_),
    .B1(_21649_),
    .B2(_21650_),
    .X(_21652_));
 sky130_fd_sc_hd__nand3_4 _50541_ (.A(_20580_),
    .B(_20540_),
    .C(_20579_),
    .Y(_21653_));
 sky130_fd_sc_hd__o211a_1 _50542_ (.A1(_21651_),
    .A2(_21652_),
    .B1(_20579_),
    .C1(_21653_),
    .X(_21654_));
 sky130_fd_sc_hd__a211o_1 _50543_ (.A1(_20579_),
    .A2(_21653_),
    .B1(net113),
    .C1(_21652_),
    .X(_21655_));
 sky130_fd_sc_hd__or2b_1 _50544_ (.A(_21654_),
    .B_N(_21655_),
    .X(_21656_));
 sky130_fd_sc_hd__xor2_1 _50545_ (.A(_21557_),
    .B(_21656_),
    .X(_21657_));
 sky130_fd_sc_hd__and2_1 _50546_ (.A(_21555_),
    .B(_21657_),
    .X(_21658_));
 sky130_fd_sc_hd__nor2_1 _50547_ (.A(_21555_),
    .B(_21657_),
    .Y(_21659_));
 sky130_fd_sc_hd__or2_1 _50548_ (.A(_21658_),
    .B(_21659_),
    .X(_21660_));
 sky130_fd_sc_hd__a21o_1 _50549_ (.A1(_20653_),
    .A2(_20655_),
    .B1(_21660_),
    .X(_21661_));
 sky130_fd_sc_hd__o211ai_1 _50550_ (.A1(_20512_),
    .A2(_20654_),
    .B1(_21660_),
    .C1(_20653_),
    .Y(_21662_));
 sky130_fd_sc_hd__nand2_1 _50551_ (.A(_21661_),
    .B(_21662_),
    .Y(_21663_));
 sky130_fd_sc_hd__xnor2_1 _50552_ (.A(_21353_),
    .B(_21663_),
    .Y(_21664_));
 sky130_fd_sc_hd__a21o_1 _50553_ (.A1(_20658_),
    .A2(_20659_),
    .B1(_21664_),
    .X(_21665_));
 sky130_fd_sc_hd__and2_1 _50554_ (.A(_20658_),
    .B(_20659_),
    .X(_21666_));
 sky130_fd_sc_hd__nand2_1 _50555_ (.A(_21664_),
    .B(_21666_),
    .Y(_21667_));
 sky130_fd_sc_hd__nand2_1 _50556_ (.A(_21665_),
    .B(_21667_),
    .Y(_21668_));
 sky130_fd_sc_hd__a21bo_1 _50557_ (.A1(_21199_),
    .A2(_21200_),
    .B1_N(_21668_),
    .X(_21669_));
 sky130_fd_sc_hd__nand3b_2 _50558_ (.A_N(_21668_),
    .B(_21199_),
    .C(_21200_),
    .Y(_21670_));
 sky130_fd_sc_hd__nand2_1 _50559_ (.A(_21669_),
    .B(_21670_),
    .Y(_21671_));
 sky130_fd_sc_hd__a21o_1 _50560_ (.A1(_20982_),
    .A2(_20983_),
    .B1(_21671_),
    .X(_21672_));
 sky130_fd_sc_hd__inv_2 _50561_ (.A(_21672_),
    .Y(_21673_));
 sky130_fd_sc_hd__and3_1 _50562_ (.A(_20982_),
    .B(_20983_),
    .C(_21671_),
    .X(_21674_));
 sky130_fd_sc_hd__a21oi_4 _50563_ (.A1(_20277_),
    .A2(_20279_),
    .B1(_20276_),
    .Y(_21675_));
 sky130_fd_sc_hd__inv_2 _50564_ (.A(_20813_),
    .Y(_21676_));
 sky130_fd_sc_hd__a32o_1 _50565_ (.A1(_20178_),
    .A2(_20168_),
    .A3(_20172_),
    .B1(_20182_),
    .B2(_20228_),
    .X(_21677_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50566_ (.A(_08393_),
    .X(_21678_));
 sky130_fd_sc_hd__clkbuf_2 _50567_ (.A(net404),
    .X(_21679_));
 sky130_fd_sc_hd__or2_1 _50568_ (.A(_21679_),
    .B(_20061_),
    .X(_21680_));
 sky130_fd_sc_hd__nor2_1 _50569_ (.A(net405),
    .B(net404),
    .Y(_21681_));
 sky130_fd_sc_hd__and2_1 _50570_ (.A(\delay_line[12][7] ),
    .B(net404),
    .X(_21682_));
 sky130_fd_sc_hd__a2bb2o_2 _50571_ (.A1_N(_21681_),
    .A2_N(_21682_),
    .B1(\delay_line[12][6] ),
    .B2(_20060_),
    .X(_21683_));
 sky130_fd_sc_hd__a21oi_2 _50572_ (.A1(_21680_),
    .A2(_21683_),
    .B1(_08470_),
    .Y(_21684_));
 sky130_fd_sc_hd__o211ai_4 _50573_ (.A1(_21679_),
    .A2(_20061_),
    .B1(_12152_),
    .C1(_21683_),
    .Y(_21685_));
 sky130_fd_sc_hd__nand3b_2 _50574_ (.A_N(_21684_),
    .B(\delay_line[13][0] ),
    .C(_21685_),
    .Y(_21686_));
 sky130_fd_sc_hd__and3_1 _50575_ (.A(_21683_),
    .B(_08470_),
    .C(_21680_),
    .X(_21687_));
 sky130_fd_sc_hd__o21ai_1 _50576_ (.A1(_21687_),
    .A2(_21684_),
    .B1(_23194_),
    .Y(_21688_));
 sky130_fd_sc_hd__nand2_1 _50577_ (.A(_21686_),
    .B(_21688_),
    .Y(_21689_));
 sky130_fd_sc_hd__xnor2_1 _50578_ (.A(_20052_),
    .B(_21689_),
    .Y(_21690_));
 sky130_fd_sc_hd__o21a_1 _50579_ (.A1(_21678_),
    .A2(_20064_),
    .B1(_21690_),
    .X(_21691_));
 sky130_fd_sc_hd__nor3_1 _50580_ (.A(_21678_),
    .B(_20064_),
    .C(_21690_),
    .Y(_21692_));
 sky130_fd_sc_hd__a21o_1 _50581_ (.A1(_20038_),
    .A2(_20040_),
    .B1(_20036_),
    .X(_21693_));
 sky130_fd_sc_hd__or2_1 _50582_ (.A(_12383_),
    .B(net396),
    .X(_21694_));
 sky130_fd_sc_hd__nand2_1 _50583_ (.A(_12383_),
    .B(\delay_line[13][8] ),
    .Y(_21695_));
 sky130_fd_sc_hd__and3_1 _50584_ (.A(_21694_),
    .B(_21695_),
    .C(_19988_),
    .X(_21696_));
 sky130_fd_sc_hd__clkbuf_2 _50585_ (.A(_21696_),
    .X(_21697_));
 sky130_fd_sc_hd__a21oi_2 _50586_ (.A1(_21694_),
    .A2(_21695_),
    .B1(_19988_),
    .Y(_21698_));
 sky130_fd_sc_hd__nor2b_1 _50587_ (.A(_17934_),
    .B_N(net434),
    .Y(_21699_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50588_ (.A(_21699_),
    .X(_21700_));
 sky130_fd_sc_hd__buf_6 _50589_ (.A(\delay_line[4][5] ),
    .X(_21701_));
 sky130_fd_sc_hd__nor2_2 _50590_ (.A(_18928_),
    .B(_21701_),
    .Y(_21702_));
 sky130_fd_sc_hd__and2_2 _50591_ (.A(_18928_),
    .B(_21701_),
    .X(_21703_));
 sky130_fd_sc_hd__and2b_1 _50592_ (.A_N(net434),
    .B(\delay_line[4][2] ),
    .X(_21704_));
 sky130_fd_sc_hd__o22ai_4 _50593_ (.A1(_21702_),
    .A2(_21703_),
    .B1(_18929_),
    .B2(_21704_),
    .Y(_21705_));
 sky130_fd_sc_hd__nor2b_2 _50594_ (.A(_18928_),
    .B_N(_21701_),
    .Y(_21706_));
 sky130_fd_sc_hd__and2b_2 _50595_ (.A_N(_21701_),
    .B(_18928_),
    .X(_21707_));
 sky130_fd_sc_hd__o2bb2ai_1 _50596_ (.A1_N(\delay_line[4][4] ),
    .A2_N(_17940_),
    .B1(\delay_line[4][1] ),
    .B2(_19990_),
    .Y(_21708_));
 sky130_fd_sc_hd__o211ai_4 _50597_ (.A1(_21706_),
    .A2(_21707_),
    .B1(_21708_),
    .C1(_19992_),
    .Y(_21709_));
 sky130_fd_sc_hd__o211ai_2 _50598_ (.A1(_18923_),
    .A2(_12339_),
    .B1(_17946_),
    .C1(_19994_),
    .Y(_21710_));
 sky130_fd_sc_hd__o21ai_1 _50599_ (.A1(_18925_),
    .A2(_21710_),
    .B1(_20015_),
    .Y(_21711_));
 sky130_fd_sc_hd__o211ai_2 _50600_ (.A1(_21700_),
    .A2(_21705_),
    .B1(_21709_),
    .C1(_21711_),
    .Y(_21712_));
 sky130_fd_sc_hd__o21ai_2 _50601_ (.A1(_21699_),
    .A2(_21705_),
    .B1(_21709_),
    .Y(_21713_));
 sky130_fd_sc_hd__buf_6 _50602_ (.A(_21713_),
    .X(_21714_));
 sky130_fd_sc_hd__o21a_1 _50603_ (.A1(_18925_),
    .A2(_21710_),
    .B1(_20015_),
    .X(_21715_));
 sky130_fd_sc_hd__nand2_1 _50604_ (.A(_21714_),
    .B(_21715_),
    .Y(_21716_));
 sky130_fd_sc_hd__inv_2 _50605_ (.A(\delay_line[11][6] ),
    .Y(_21717_));
 sky130_fd_sc_hd__buf_2 _50606_ (.A(_21717_),
    .X(_21718_));
 sky130_fd_sc_hd__o21bai_4 _50607_ (.A1(_18933_),
    .A2(_20005_),
    .B1_N(\delay_line[11][1] ),
    .Y(_21719_));
 sky130_fd_sc_hd__buf_6 _50608_ (.A(\delay_line[11][6] ),
    .X(_21720_));
 sky130_fd_sc_hd__o2bb2a_1 _50609_ (.A1_N(_18933_),
    .A2_N(_20005_),
    .B1(_21720_),
    .B2(\delay_line[11][2] ),
    .X(_21721_));
 sky130_fd_sc_hd__o211ai_4 _50610_ (.A1(_12350_),
    .A2(_21718_),
    .B1(_21719_),
    .C1(_21721_),
    .Y(_21722_));
 sky130_fd_sc_hd__and2_1 _50611_ (.A(_12262_),
    .B(_21720_),
    .X(_21723_));
 sky130_fd_sc_hd__nor2_1 _50612_ (.A(_12262_),
    .B(_21720_),
    .Y(_21724_));
 sky130_fd_sc_hd__o2bb2ai_2 _50613_ (.A1_N(_21719_),
    .A2_N(_20009_),
    .B1(_21723_),
    .B2(_21724_),
    .Y(_21725_));
 sky130_fd_sc_hd__clkbuf_2 _50614_ (.A(_21725_),
    .X(_21726_));
 sky130_fd_sc_hd__a21oi_1 _50615_ (.A1(_21722_),
    .A2(_21726_),
    .B1(_20018_),
    .Y(_21727_));
 sky130_fd_sc_hd__buf_2 _50616_ (.A(_21717_),
    .X(_21728_));
 sky130_fd_sc_hd__o21ai_1 _50617_ (.A1(_12361_),
    .A2(_21728_),
    .B1(_21721_),
    .Y(_21729_));
 sky130_fd_sc_hd__o211a_1 _50618_ (.A1(_20008_),
    .A2(_21729_),
    .B1(_21726_),
    .C1(_20018_),
    .X(_21730_));
 sky130_fd_sc_hd__o2bb2ai_2 _50619_ (.A1_N(_21712_),
    .A2_N(_21716_),
    .B1(_21727_),
    .B2(_21730_),
    .Y(_21731_));
 sky130_fd_sc_hd__nand2_1 _50620_ (.A(_21722_),
    .B(_21726_),
    .Y(_21732_));
 sky130_fd_sc_hd__o2111ai_2 _50621_ (.A1(_21719_),
    .A2(_20006_),
    .B1(_18936_),
    .C1(_20007_),
    .D1(_21732_),
    .Y(_21733_));
 sky130_fd_sc_hd__o211ai_2 _50622_ (.A1(_20008_),
    .A2(_21729_),
    .B1(_21726_),
    .C1(_20018_),
    .Y(_21734_));
 sky130_fd_sc_hd__nand4_1 _50623_ (.A(_21712_),
    .B(_21716_),
    .C(_21733_),
    .D(_21734_),
    .Y(_21735_));
 sky130_fd_sc_hd__buf_2 _50624_ (.A(net455),
    .X(_21736_));
 sky130_fd_sc_hd__a21oi_1 _50625_ (.A1(_21731_),
    .A2(_21735_),
    .B1(_21736_),
    .Y(_21737_));
 sky130_fd_sc_hd__o211a_1 _50626_ (.A1(_21710_),
    .A2(_18925_),
    .B1(_20016_),
    .C1(_21714_),
    .X(_21738_));
 sky130_fd_sc_hd__o211ai_1 _50627_ (.A1(_21715_),
    .A2(_21714_),
    .B1(_21734_),
    .C1(_21733_),
    .Y(_21739_));
 sky130_fd_sc_hd__o211a_2 _50628_ (.A1(_21738_),
    .A2(_21739_),
    .B1(net455),
    .C1(_21731_),
    .X(_21740_));
 sky130_fd_sc_hd__o21bai_1 _50629_ (.A1(_21737_),
    .A2(_21740_),
    .B1_N(_20025_),
    .Y(_21741_));
 sky130_fd_sc_hd__a21o_1 _50630_ (.A1(_21731_),
    .A2(_21735_),
    .B1(net455),
    .X(_21742_));
 sky130_fd_sc_hd__o211ai_1 _50631_ (.A1(_21738_),
    .A2(_21739_),
    .B1(net455),
    .C1(_21731_),
    .Y(_21743_));
 sky130_fd_sc_hd__nand3_2 _50632_ (.A(_20025_),
    .B(_21742_),
    .C(_21743_),
    .Y(_21744_));
 sky130_fd_sc_hd__a21o_1 _50633_ (.A1(_21741_),
    .A2(_21744_),
    .B1(_19986_),
    .X(_21745_));
 sky130_fd_sc_hd__clkbuf_2 _50634_ (.A(_19986_),
    .X(_21746_));
 sky130_fd_sc_hd__nand3_1 _50635_ (.A(_21741_),
    .B(_21744_),
    .C(_21746_),
    .Y(_21747_));
 sky130_fd_sc_hd__a21o_1 _50636_ (.A1(_20030_),
    .A2(_20031_),
    .B1(_20027_),
    .X(_21748_));
 sky130_fd_sc_hd__a21oi_2 _50637_ (.A1(_21745_),
    .A2(_21747_),
    .B1(_21748_),
    .Y(_21749_));
 sky130_fd_sc_hd__inv_2 _50638_ (.A(_21744_),
    .Y(_21750_));
 sky130_fd_sc_hd__nand2_1 _50639_ (.A(_21741_),
    .B(_21746_),
    .Y(_21751_));
 sky130_fd_sc_hd__o211a_1 _50640_ (.A1(_21750_),
    .A2(_21751_),
    .B1(_21748_),
    .C1(_21745_),
    .X(_21752_));
 sky130_fd_sc_hd__o22ai_4 _50641_ (.A1(_21697_),
    .A2(_21698_),
    .B1(_21749_),
    .B2(_21752_),
    .Y(_21753_));
 sky130_fd_sc_hd__or2_1 _50642_ (.A(_21697_),
    .B(_21698_),
    .X(_21754_));
 sky130_fd_sc_hd__a21o_1 _50643_ (.A1(_21745_),
    .A2(_21747_),
    .B1(_21748_),
    .X(_21755_));
 sky130_fd_sc_hd__o211ai_4 _50644_ (.A1(_21750_),
    .A2(_21751_),
    .B1(_21748_),
    .C1(_21745_),
    .Y(_21756_));
 sky130_fd_sc_hd__nand3b_2 _50645_ (.A_N(_21754_),
    .B(_21755_),
    .C(_21756_),
    .Y(_21757_));
 sky130_fd_sc_hd__nand3_2 _50646_ (.A(_21693_),
    .B(_21753_),
    .C(_21757_),
    .Y(_21758_));
 sky130_fd_sc_hd__o21bai_1 _50647_ (.A1(_21749_),
    .A2(_21752_),
    .B1_N(_21754_),
    .Y(_21759_));
 sky130_fd_sc_hd__o31a_1 _50648_ (.A1(_19984_),
    .A2(_19985_),
    .A3(_20034_),
    .B1(_20039_),
    .X(_21760_));
 sky130_fd_sc_hd__o211ai_1 _50649_ (.A1(_21697_),
    .A2(_21698_),
    .B1(_21755_),
    .C1(_21756_),
    .Y(_21761_));
 sky130_fd_sc_hd__nand3_1 _50650_ (.A(_21759_),
    .B(_21760_),
    .C(_21761_),
    .Y(_21762_));
 sky130_fd_sc_hd__nand2_2 _50651_ (.A(_18913_),
    .B(_20048_),
    .Y(_21763_));
 sky130_fd_sc_hd__a21o_1 _50652_ (.A1(\delay_line[13][5] ),
    .A2(_20046_),
    .B1(\delay_line[13][6] ),
    .X(_21764_));
 sky130_fd_sc_hd__a21o_1 _50653_ (.A1(_21763_),
    .A2(_21764_),
    .B1(\delay_line[13][2] ),
    .X(_21765_));
 sky130_fd_sc_hd__nand3_2 _50654_ (.A(_21763_),
    .B(_21764_),
    .C(\delay_line[13][2] ),
    .Y(_21766_));
 sky130_fd_sc_hd__nand4_1 _50655_ (.A(_21765_),
    .B(_18947_),
    .C(_12570_),
    .D(_21766_),
    .Y(_21767_));
 sky130_fd_sc_hd__a32o_1 _50656_ (.A1(_12570_),
    .A2(_17950_),
    .A3(_18948_),
    .B1(_21766_),
    .B2(_21765_),
    .X(_21768_));
 sky130_fd_sc_hd__o311a_1 _50657_ (.A1(_18914_),
    .A2(_20047_),
    .A3(_20048_),
    .B1(_21767_),
    .C1(_21768_),
    .X(_21769_));
 sky130_fd_sc_hd__a21oi_1 _50658_ (.A1(_21767_),
    .A2(_21768_),
    .B1(_20053_),
    .Y(_21770_));
 sky130_fd_sc_hd__o2bb2ai_1 _50659_ (.A1_N(_21758_),
    .A2_N(_21762_),
    .B1(_21769_),
    .B2(_21770_),
    .Y(_21771_));
 sky130_fd_sc_hd__nor2_1 _50660_ (.A(_20052_),
    .B(_20054_),
    .Y(_21772_));
 sky130_fd_sc_hd__a32oi_4 _50661_ (.A1(_19981_),
    .A2(_20037_),
    .A3(_20041_),
    .B1(_20045_),
    .B2(_21772_),
    .Y(_21773_));
 sky130_fd_sc_hd__nand2_1 _50662_ (.A(_21767_),
    .B(_21768_),
    .Y(_21774_));
 sky130_fd_sc_hd__nor2_1 _50663_ (.A(_20053_),
    .B(_21774_),
    .Y(_21775_));
 sky130_fd_sc_hd__o31a_1 _50664_ (.A1(_18914_),
    .A2(_20047_),
    .A3(_20048_),
    .B1(_21774_),
    .X(_21776_));
 sky130_fd_sc_hd__clkbuf_2 _50665_ (.A(_21762_),
    .X(_21777_));
 sky130_fd_sc_hd__o211ai_1 _50666_ (.A1(_21775_),
    .A2(_21776_),
    .B1(_21758_),
    .C1(_21777_),
    .Y(_21778_));
 sky130_fd_sc_hd__nand3_1 _50667_ (.A(_21771_),
    .B(_21773_),
    .C(_21778_),
    .Y(_21779_));
 sky130_fd_sc_hd__o21ai_1 _50668_ (.A1(_21691_),
    .A2(_21692_),
    .B1(_21779_),
    .Y(_21780_));
 sky130_fd_sc_hd__inv_2 _50669_ (.A(_21773_),
    .Y(_21781_));
 sky130_fd_sc_hd__o2bb2ai_1 _50670_ (.A1_N(_21758_),
    .A2_N(_21777_),
    .B1(_21775_),
    .B2(_21776_),
    .Y(_21782_));
 sky130_fd_sc_hd__o211ai_2 _50671_ (.A1(_21769_),
    .A2(_21770_),
    .B1(_21758_),
    .C1(_21777_),
    .Y(_21783_));
 sky130_fd_sc_hd__and3_1 _50672_ (.A(_21781_),
    .B(_21782_),
    .C(_21783_),
    .X(_21784_));
 sky130_fd_sc_hd__a32o_1 _50673_ (.A1(_19980_),
    .A2(_20055_),
    .A3(_20058_),
    .B1(_20074_),
    .B2(_20069_),
    .X(_21785_));
 sky130_fd_sc_hd__nand3_1 _50674_ (.A(_21781_),
    .B(_21782_),
    .C(_21783_),
    .Y(_21786_));
 sky130_fd_sc_hd__clkbuf_2 _50675_ (.A(_21779_),
    .X(_21787_));
 sky130_fd_sc_hd__nor3b_1 _50676_ (.A(_21678_),
    .B(_20064_),
    .C_N(_21690_),
    .Y(_21788_));
 sky130_fd_sc_hd__o21ba_1 _50677_ (.A1(_21678_),
    .A2(_20064_),
    .B1_N(_21690_),
    .X(_21789_));
 sky130_fd_sc_hd__o2bb2ai_1 _50678_ (.A1_N(_21786_),
    .A2_N(_21787_),
    .B1(net170),
    .B2(_21789_),
    .Y(_21790_));
 sky130_fd_sc_hd__o211ai_2 _50679_ (.A1(_21780_),
    .A2(_21784_),
    .B1(_21785_),
    .C1(_21790_),
    .Y(_21791_));
 sky130_fd_sc_hd__o2bb2ai_1 _50680_ (.A1_N(_21786_),
    .A2_N(_21787_),
    .B1(_21691_),
    .B2(_21692_),
    .Y(_21792_));
 sky130_fd_sc_hd__inv_2 _50681_ (.A(_21785_),
    .Y(_21793_));
 sky130_fd_sc_hd__o211ai_1 _50682_ (.A1(net170),
    .A2(_21789_),
    .B1(_21786_),
    .C1(_21787_),
    .Y(_21794_));
 sky130_fd_sc_hd__nand3_2 _50683_ (.A(_21792_),
    .B(_21793_),
    .C(_21794_),
    .Y(_21795_));
 sky130_fd_sc_hd__or3_1 _50684_ (.A(_19969_),
    .B(_19970_),
    .C(_18896_),
    .X(_21796_));
 sky130_fd_sc_hd__o21ai_1 _50685_ (.A1(_19973_),
    .A2(_19968_),
    .B1(_21796_),
    .Y(_21797_));
 sky130_fd_sc_hd__a21oi_2 _50686_ (.A1(_18920_),
    .A2(_20065_),
    .B1(_20067_),
    .Y(_21798_));
 sky130_fd_sc_hd__nand2_1 _50687_ (.A(_18987_),
    .B(_18984_),
    .Y(_21799_));
 sky130_fd_sc_hd__buf_2 _50688_ (.A(\delay_line[10][8] ),
    .X(_21800_));
 sky130_fd_sc_hd__buf_2 _50689_ (.A(_21800_),
    .X(_21801_));
 sky130_fd_sc_hd__a21oi_2 _50690_ (.A1(_02436_),
    .A2(_02425_),
    .B1(_21801_),
    .Y(_21802_));
 sky130_fd_sc_hd__and3_1 _50691_ (.A(_02436_),
    .B(_02414_),
    .C(_21800_),
    .X(_21803_));
 sky130_fd_sc_hd__or4_1 _50692_ (.A(_20062_),
    .B(_21799_),
    .C(_21802_),
    .D(_21803_),
    .X(_21804_));
 sky130_fd_sc_hd__clkbuf_4 _50693_ (.A(_20062_),
    .X(_21805_));
 sky130_fd_sc_hd__o22ai_4 _50694_ (.A1(_21805_),
    .A2(_21799_),
    .B1(_21802_),
    .B2(_21803_),
    .Y(_21806_));
 sky130_fd_sc_hd__nand2_1 _50695_ (.A(_21804_),
    .B(_21806_),
    .Y(_21807_));
 sky130_fd_sc_hd__or3b_1 _50696_ (.A(_08437_),
    .B(_02447_),
    .C_N(_23238_),
    .X(_21808_));
 sky130_fd_sc_hd__o31a_1 _50697_ (.A1(_18986_),
    .A2(_17995_),
    .A3(_02799_),
    .B1(_21808_),
    .X(_21809_));
 sky130_fd_sc_hd__xor2_1 _50698_ (.A(_21807_),
    .B(_21809_),
    .X(_21810_));
 sky130_fd_sc_hd__nand2_1 _50699_ (.A(_11691_),
    .B(net419),
    .Y(_21811_));
 sky130_fd_sc_hd__inv_2 _50700_ (.A(net419),
    .Y(_21812_));
 sky130_fd_sc_hd__nand2_1 _50701_ (.A(_21812_),
    .B(\delay_line[10][0] ),
    .Y(_21813_));
 sky130_fd_sc_hd__and3_1 _50702_ (.A(_21811_),
    .B(_21813_),
    .C(_19961_),
    .X(_21814_));
 sky130_fd_sc_hd__a21oi_1 _50703_ (.A1(_21811_),
    .A2(_21813_),
    .B1(_19961_),
    .Y(_21815_));
 sky130_fd_sc_hd__or2_2 _50704_ (.A(_21814_),
    .B(_21815_),
    .X(_21816_));
 sky130_fd_sc_hd__buf_1 _50705_ (.A(\delay_line[10][3] ),
    .X(_21817_));
 sky130_fd_sc_hd__nor2_1 _50706_ (.A(_02821_),
    .B(_21817_),
    .Y(_21818_));
 sky130_fd_sc_hd__and2_1 _50707_ (.A(_02821_),
    .B(_21817_),
    .X(_21819_));
 sky130_fd_sc_hd__o21bai_1 _50708_ (.A1(_21818_),
    .A2(_21819_),
    .B1_N(_17919_),
    .Y(_21820_));
 sky130_fd_sc_hd__buf_2 _50709_ (.A(_19956_),
    .X(_21821_));
 sky130_fd_sc_hd__nand2_1 _50710_ (.A(_02821_),
    .B(_08701_),
    .Y(_21822_));
 sky130_fd_sc_hd__nand3b_1 _50711_ (.A_N(_21818_),
    .B(_21822_),
    .C(_17919_),
    .Y(_21823_));
 sky130_fd_sc_hd__nand4_1 _50712_ (.A(_21820_),
    .B(_21821_),
    .C(_21823_),
    .D(_19959_),
    .Y(_21824_));
 sky130_fd_sc_hd__a22o_1 _50713_ (.A1(_21821_),
    .A2(_19959_),
    .B1(_21823_),
    .B2(_21820_),
    .X(_21825_));
 sky130_fd_sc_hd__nand2_1 _50714_ (.A(_21824_),
    .B(_21825_),
    .Y(_21826_));
 sky130_fd_sc_hd__xor2_2 _50715_ (.A(_21816_),
    .B(_21826_),
    .X(_21827_));
 sky130_fd_sc_hd__xnor2_1 _50716_ (.A(_21810_),
    .B(_21827_),
    .Y(_21828_));
 sky130_fd_sc_hd__xnor2_1 _50717_ (.A(_21798_),
    .B(_21828_),
    .Y(_21829_));
 sky130_fd_sc_hd__and2_1 _50718_ (.A(_21797_),
    .B(_21829_),
    .X(_21830_));
 sky130_fd_sc_hd__nor2_1 _50719_ (.A(_21797_),
    .B(_21829_),
    .Y(_21831_));
 sky130_fd_sc_hd__o2bb2ai_1 _50720_ (.A1_N(_21791_),
    .A2_N(_21795_),
    .B1(_21830_),
    .B2(_21831_),
    .Y(_21832_));
 sky130_fd_sc_hd__o21ai_2 _50721_ (.A1(_20155_),
    .A2(_20081_),
    .B1(_20096_),
    .Y(_21833_));
 sky130_fd_sc_hd__inv_2 _50722_ (.A(_21833_),
    .Y(_21834_));
 sky130_fd_sc_hd__or2b_1 _50723_ (.A(_21829_),
    .B_N(_21797_),
    .X(_21835_));
 sky130_fd_sc_hd__inv_2 _50724_ (.A(_21835_),
    .Y(_21836_));
 sky130_fd_sc_hd__o211a_1 _50725_ (.A1(_19973_),
    .A2(_19968_),
    .B1(_21796_),
    .C1(_21829_),
    .X(_21837_));
 sky130_fd_sc_hd__o211ai_1 _50726_ (.A1(_21836_),
    .A2(_21837_),
    .B1(_21791_),
    .C1(_21795_),
    .Y(_21838_));
 sky130_fd_sc_hd__nand3_1 _50727_ (.A(_21832_),
    .B(_21834_),
    .C(_21838_),
    .Y(_21839_));
 sky130_fd_sc_hd__clkbuf_2 _50728_ (.A(_21839_),
    .X(_21840_));
 sky130_fd_sc_hd__nor2_1 _50729_ (.A(_20138_),
    .B(_20139_),
    .Y(_21841_));
 sky130_fd_sc_hd__a21o_1 _50730_ (.A1(_20140_),
    .A2(_21841_),
    .B1(_20138_),
    .X(_21842_));
 sky130_fd_sc_hd__clkbuf_2 _50731_ (.A(_20125_),
    .X(_21843_));
 sky130_fd_sc_hd__a21bo_1 _50732_ (.A1(_18867_),
    .A2(net420),
    .B1_N(_17912_),
    .X(_21844_));
 sky130_fd_sc_hd__o211ai_4 _50733_ (.A1(_20122_),
    .A2(_21843_),
    .B1(_02843_),
    .C1(_21844_),
    .Y(_21845_));
 sky130_fd_sc_hd__o21bai_2 _50734_ (.A1(_20128_),
    .A2(_20126_),
    .B1_N(_02843_),
    .Y(_21846_));
 sky130_fd_sc_hd__a22o_1 _50735_ (.A1(_25040_),
    .A2(_08712_),
    .B1(_21845_),
    .B2(_21846_),
    .X(_21847_));
 sky130_fd_sc_hd__nand4_1 _50736_ (.A(_21845_),
    .B(_21846_),
    .C(_25051_),
    .D(_08712_),
    .Y(_21848_));
 sky130_fd_sc_hd__o2111a_1 _50737_ (.A1(_17915_),
    .A2(_20123_),
    .B1(_20124_),
    .C1(_20127_),
    .D1(_20130_),
    .X(_21849_));
 sky130_fd_sc_hd__and3_1 _50738_ (.A(_21847_),
    .B(_21848_),
    .C(_21849_),
    .X(_21850_));
 sky130_fd_sc_hd__a21oi_1 _50739_ (.A1(_21847_),
    .A2(_21848_),
    .B1(_21849_),
    .Y(_21851_));
 sky130_fd_sc_hd__a21boi_2 _50740_ (.A1(_19963_),
    .A2(_18901_),
    .B1_N(_19965_),
    .Y(_21852_));
 sky130_fd_sc_hd__o21a_1 _50741_ (.A1(_21850_),
    .A2(_21851_),
    .B1(_21852_),
    .X(_21853_));
 sky130_fd_sc_hd__nor3_1 _50742_ (.A(_21852_),
    .B(_21850_),
    .C(_21851_),
    .Y(_21854_));
 sky130_fd_sc_hd__or3_1 _50743_ (.A(_20137_),
    .B(_21853_),
    .C(net207),
    .X(_21855_));
 sky130_fd_sc_hd__o21ai_1 _50744_ (.A1(_21853_),
    .A2(net207),
    .B1(_20137_),
    .Y(_21856_));
 sky130_fd_sc_hd__and3_1 _50745_ (.A(_21842_),
    .B(_21855_),
    .C(_21856_),
    .X(_21857_));
 sky130_fd_sc_hd__a221oi_2 _50746_ (.A1(_20140_),
    .A2(_21841_),
    .B1(_21855_),
    .B2(_21856_),
    .C1(_20138_),
    .Y(_21858_));
 sky130_fd_sc_hd__nor2_1 _50747_ (.A(_21857_),
    .B(_21858_),
    .Y(_21859_));
 sky130_fd_sc_hd__o221a_1 _50748_ (.A1(_11822_),
    .A2(_18850_),
    .B1(_20100_),
    .B2(_20103_),
    .C1(_18847_),
    .X(_21860_));
 sky130_fd_sc_hd__o21ai_2 _50749_ (.A1(_11833_),
    .A2(_21860_),
    .B1(_20107_),
    .Y(_21861_));
 sky130_fd_sc_hd__clkbuf_2 _50750_ (.A(\delay_line[7][8] ),
    .X(_21862_));
 sky130_fd_sc_hd__xnor2_1 _50751_ (.A(_23040_),
    .B(_21862_),
    .Y(_21863_));
 sky130_fd_sc_hd__nand2_1 _50752_ (.A(_21861_),
    .B(_21863_),
    .Y(_21864_));
 sky130_fd_sc_hd__or2_1 _50753_ (.A(_21863_),
    .B(_21861_),
    .X(_21865_));
 sky130_fd_sc_hd__and2_1 _50754_ (.A(_21864_),
    .B(_21865_),
    .X(_21866_));
 sky130_fd_sc_hd__clkbuf_2 _50755_ (.A(\delay_line[8][8] ),
    .X(_21867_));
 sky130_fd_sc_hd__nand2b_2 _50756_ (.A_N(\delay_line[9][0] ),
    .B(_21867_),
    .Y(_21868_));
 sky130_fd_sc_hd__clkbuf_2 _50757_ (.A(net424),
    .X(_21869_));
 sky130_fd_sc_hd__or2b_1 _50758_ (.A(_21869_),
    .B_N(\delay_line[9][0] ),
    .X(_21870_));
 sky130_fd_sc_hd__and3_1 _50759_ (.A(_18040_),
    .B(_20099_),
    .C(_20104_),
    .X(_21871_));
 sky130_fd_sc_hd__or3b_2 _50760_ (.A(_21871_),
    .B(_20100_),
    .C_N(_03183_),
    .X(_21872_));
 sky130_fd_sc_hd__o21bai_1 _50761_ (.A1(_21871_),
    .A2(_20100_),
    .B1_N(_09009_),
    .Y(_21873_));
 sky130_fd_sc_hd__and4_1 _50762_ (.A(_21868_),
    .B(_21870_),
    .C(_21872_),
    .D(_21873_),
    .X(_21874_));
 sky130_fd_sc_hd__buf_1 _50763_ (.A(_21874_),
    .X(_21875_));
 sky130_fd_sc_hd__a22oi_2 _50764_ (.A1(_21868_),
    .A2(_21870_),
    .B1(_21872_),
    .B2(_21873_),
    .Y(_21876_));
 sky130_fd_sc_hd__nand3_1 _50765_ (.A(_20109_),
    .B(_20110_),
    .C(_08877_),
    .Y(_21877_));
 sky130_fd_sc_hd__o21a_1 _50766_ (.A1(_21875_),
    .A2(_21876_),
    .B1(_21877_),
    .X(_21878_));
 sky130_fd_sc_hd__nor3_1 _50767_ (.A(_21874_),
    .B(_21876_),
    .C(_21877_),
    .Y(_21879_));
 sky130_fd_sc_hd__nor2_1 _50768_ (.A(_21878_),
    .B(_21879_),
    .Y(_21880_));
 sky130_fd_sc_hd__xor2_2 _50769_ (.A(_21866_),
    .B(_21880_),
    .X(_21881_));
 sky130_fd_sc_hd__o21a_1 _50770_ (.A1(_21859_),
    .A2(_21881_),
    .B1(_20091_),
    .X(_21882_));
 sky130_fd_sc_hd__or3b_1 _50771_ (.A(_21857_),
    .B(_21858_),
    .C_N(_21881_),
    .X(_21883_));
 sky130_fd_sc_hd__or2_1 _50772_ (.A(_21859_),
    .B(_21881_),
    .X(_21884_));
 sky130_fd_sc_hd__a21oi_1 _50773_ (.A1(_21883_),
    .A2(_21884_),
    .B1(_20091_),
    .Y(_21885_));
 sky130_fd_sc_hd__a21o_1 _50774_ (.A1(_21882_),
    .A2(_21883_),
    .B1(_21885_),
    .X(_21886_));
 sky130_fd_sc_hd__a21oi_1 _50775_ (.A1(_20120_),
    .A2(_20142_),
    .B1(_20145_),
    .Y(_21887_));
 sky130_fd_sc_hd__and2_1 _50776_ (.A(_21886_),
    .B(_21887_),
    .X(_21888_));
 sky130_fd_sc_hd__nor2_1 _50777_ (.A(_21887_),
    .B(_21886_),
    .Y(_21889_));
 sky130_fd_sc_hd__nor2_1 _50778_ (.A(_21888_),
    .B(_21889_),
    .Y(_21890_));
 sky130_fd_sc_hd__nand2_1 _50779_ (.A(_21840_),
    .B(_21890_),
    .Y(_21891_));
 sky130_fd_sc_hd__or2_1 _50780_ (.A(_21830_),
    .B(_21831_),
    .X(_21892_));
 sky130_fd_sc_hd__nand2_1 _50781_ (.A(_21795_),
    .B(_21892_),
    .Y(_21893_));
 sky130_fd_sc_hd__o211a_1 _50782_ (.A1(_21780_),
    .A2(_21784_),
    .B1(_21785_),
    .C1(_21790_),
    .X(_21894_));
 sky130_fd_sc_hd__o2bb2ai_1 _50783_ (.A1_N(_21791_),
    .A2_N(_21795_),
    .B1(_21836_),
    .B2(_21837_),
    .Y(_21895_));
 sky130_fd_sc_hd__o211a_2 _50784_ (.A1(_21893_),
    .A2(_21894_),
    .B1(_21833_),
    .C1(_21895_),
    .X(_21896_));
 sky130_fd_sc_hd__a21o_1 _50785_ (.A1(_20098_),
    .A2(_20153_),
    .B1(_20159_),
    .X(_21897_));
 sky130_fd_sc_hd__o211ai_2 _50786_ (.A1(_21893_),
    .A2(_21894_),
    .B1(_21833_),
    .C1(_21895_),
    .Y(_21898_));
 sky130_fd_sc_hd__o2bb2ai_1 _50787_ (.A1_N(_21898_),
    .A2_N(_21839_),
    .B1(_21888_),
    .B2(_21889_),
    .Y(_21899_));
 sky130_fd_sc_hd__o211ai_4 _50788_ (.A1(_21891_),
    .A2(_21896_),
    .B1(_21897_),
    .C1(_21899_),
    .Y(_21900_));
 sky130_fd_sc_hd__a21bo_1 _50789_ (.A1(_21898_),
    .A2(_21840_),
    .B1_N(_21890_),
    .X(_21901_));
 sky130_fd_sc_hd__o211ai_2 _50790_ (.A1(_21888_),
    .A2(_21889_),
    .B1(_21898_),
    .C1(_21840_),
    .Y(_21902_));
 sky130_fd_sc_hd__inv_2 _50791_ (.A(_21897_),
    .Y(_21903_));
 sky130_fd_sc_hd__nand3_2 _50792_ (.A(_21901_),
    .B(_21902_),
    .C(_21903_),
    .Y(_21904_));
 sky130_fd_sc_hd__a21oi_1 _50793_ (.A1(_19881_),
    .A2(_19945_),
    .B1(_19947_),
    .Y(_21905_));
 sky130_fd_sc_hd__buf_2 _50794_ (.A(_19857_),
    .X(_21906_));
 sky130_fd_sc_hd__o21ai_2 _50795_ (.A1(_11954_),
    .A2(_08954_),
    .B1(_21906_),
    .Y(_21907_));
 sky130_fd_sc_hd__a21o_1 _50796_ (.A1(_11965_),
    .A2(_08965_),
    .B1(_21907_),
    .X(_21908_));
 sky130_fd_sc_hd__nand2_2 _50797_ (.A(_11954_),
    .B(_08954_),
    .Y(_21909_));
 sky130_fd_sc_hd__inv_2 _50798_ (.A(\delay_line[7][4] ),
    .Y(_21910_));
 sky130_fd_sc_hd__inv_2 _50799_ (.A(\delay_line[7][3] ),
    .Y(_21911_));
 sky130_fd_sc_hd__nand2_1 _50800_ (.A(_21910_),
    .B(_21911_),
    .Y(_21912_));
 sky130_fd_sc_hd__a21o_1 _50801_ (.A1(_21909_),
    .A2(_21912_),
    .B1(_21906_),
    .X(_21913_));
 sky130_fd_sc_hd__and4bb_1 _50802_ (.A_N(_19858_),
    .B_N(_19861_),
    .C(_21908_),
    .D(_21913_),
    .X(_21914_));
 sky130_fd_sc_hd__a2bb2o_1 _50803_ (.A1_N(_19858_),
    .A2_N(_19861_),
    .B1(_21908_),
    .B2(_21913_),
    .X(_21915_));
 sky130_fd_sc_hd__and2b_1 _50804_ (.A_N(\delay_line[7][0] ),
    .B(\delay_line[6][8] ),
    .X(_21916_));
 sky130_fd_sc_hd__nor2_1 _50805_ (.A(\delay_line[6][8] ),
    .B(_22963_),
    .Y(_21917_));
 sky130_fd_sc_hd__o22a_1 _50806_ (.A1(_03139_),
    .A2(_21911_),
    .B1(_21916_),
    .B2(_21917_),
    .X(_21918_));
 sky130_fd_sc_hd__nor4_1 _50807_ (.A(_03139_),
    .B(_21911_),
    .C(_21916_),
    .D(_21917_),
    .Y(_21919_));
 sky130_fd_sc_hd__nor2_1 _50808_ (.A(_21918_),
    .B(_21919_),
    .Y(_21920_));
 sky130_fd_sc_hd__nand3b_1 _50809_ (.A_N(_21914_),
    .B(_21915_),
    .C(_21920_),
    .Y(_21921_));
 sky130_fd_sc_hd__o2bb2a_1 _50810_ (.A1_N(_21908_),
    .A2_N(_21913_),
    .B1(_19858_),
    .B2(_19861_),
    .X(_21922_));
 sky130_fd_sc_hd__o22ai_2 _50811_ (.A1(_21918_),
    .A2(_21919_),
    .B1(_21914_),
    .B2(_21922_),
    .Y(_21923_));
 sky130_fd_sc_hd__nand4_1 _50812_ (.A(_20115_),
    .B(_21921_),
    .C(_21923_),
    .D(_11943_),
    .Y(_21924_));
 sky130_fd_sc_hd__a22o_1 _50813_ (.A1(_11943_),
    .A2(_20115_),
    .B1(_21921_),
    .B2(_21923_),
    .X(_21925_));
 sky130_fd_sc_hd__a31o_1 _50814_ (.A1(_19864_),
    .A2(_03458_),
    .A3(_03238_),
    .B1(_19863_),
    .X(_21926_));
 sky130_fd_sc_hd__a21o_1 _50815_ (.A1(_21924_),
    .A2(_21925_),
    .B1(_21926_),
    .X(_21927_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50816_ (.A(_21924_),
    .X(_21928_));
 sky130_fd_sc_hd__nand3_2 _50817_ (.A(_21926_),
    .B(_21928_),
    .C(_21925_),
    .Y(_21929_));
 sky130_fd_sc_hd__nand2_1 _50818_ (.A(_21927_),
    .B(_21929_),
    .Y(_21930_));
 sky130_fd_sc_hd__a21oi_1 _50819_ (.A1(_20114_),
    .A2(_20118_),
    .B1(_21930_),
    .Y(_21931_));
 sky130_fd_sc_hd__o311a_1 _50820_ (.A1(_18859_),
    .A2(_20111_),
    .A3(_20112_),
    .B1(_20118_),
    .C1(_21930_),
    .X(_21932_));
 sky130_fd_sc_hd__o211ai_2 _50821_ (.A1(_21931_),
    .A2(_21932_),
    .B1(_19869_),
    .C1(_19872_),
    .Y(_21933_));
 sky130_fd_sc_hd__a211o_1 _50822_ (.A1(_19869_),
    .A2(_19872_),
    .B1(_21931_),
    .C1(_21932_),
    .X(_21934_));
 sky130_fd_sc_hd__o211ai_2 _50823_ (.A1(_19874_),
    .A2(_19877_),
    .B1(_21933_),
    .C1(_21934_),
    .Y(_21935_));
 sky130_fd_sc_hd__a211oi_1 _50824_ (.A1(_21933_),
    .A2(_21934_),
    .B1(_19874_),
    .C1(_19877_),
    .Y(_21936_));
 sky130_fd_sc_hd__inv_2 _50825_ (.A(_21936_),
    .Y(_21937_));
 sky130_fd_sc_hd__a31o_1 _50826_ (.A1(_19920_),
    .A2(_19921_),
    .A3(_19922_),
    .B1(_03590_),
    .X(_21938_));
 sky130_fd_sc_hd__or2b_1 _50827_ (.A(_19047_),
    .B_N(net442),
    .X(_21939_));
 sky130_fd_sc_hd__or2b_1 _50828_ (.A(net442),
    .B_N(_19047_),
    .X(_21940_));
 sky130_fd_sc_hd__and2b_1 _50829_ (.A_N(_18099_),
    .B(_19885_),
    .X(_21941_));
 sky130_fd_sc_hd__nand3_1 _50830_ (.A(_21939_),
    .B(_21940_),
    .C(_21941_),
    .Y(_21942_));
 sky130_fd_sc_hd__a21o_1 _50831_ (.A1(_21939_),
    .A2(_21940_),
    .B1(_21941_),
    .X(_21943_));
 sky130_fd_sc_hd__nand2_1 _50832_ (.A(_21942_),
    .B(_21943_),
    .Y(_21944_));
 sky130_fd_sc_hd__a21o_1 _50833_ (.A1(_19924_),
    .A2(_21938_),
    .B1(_21944_),
    .X(_21945_));
 sky130_fd_sc_hd__o211ai_1 _50834_ (.A1(_19920_),
    .A2(_19883_),
    .B1(_21938_),
    .C1(_21944_),
    .Y(_21946_));
 sky130_fd_sc_hd__nand3b_1 _50835_ (.A_N(_19890_),
    .B(_21945_),
    .C(_21946_),
    .Y(_21947_));
 sky130_fd_sc_hd__a32o_1 _50836_ (.A1(_19888_),
    .A2(_19886_),
    .A3(_19887_),
    .B1(_21945_),
    .B2(_21946_),
    .X(_21948_));
 sky130_fd_sc_hd__and4b_1 _50837_ (.A_N(_19930_),
    .B(_19932_),
    .C(_19883_),
    .D(_18107_),
    .X(_21949_));
 sky130_fd_sc_hd__a211oi_2 _50838_ (.A1(_21947_),
    .A2(_21948_),
    .B1(_21949_),
    .C1(_19936_),
    .Y(_21950_));
 sky130_fd_sc_hd__o211a_1 _50839_ (.A1(_21949_),
    .A2(_19936_),
    .B1(_21947_),
    .C1(_21948_),
    .X(_21951_));
 sky130_fd_sc_hd__a211oi_1 _50840_ (.A1(_19891_),
    .A2(_19893_),
    .B1(_21950_),
    .C1(_21951_),
    .Y(_21952_));
 sky130_fd_sc_hd__o211a_1 _50841_ (.A1(_21950_),
    .A2(_21951_),
    .B1(_19891_),
    .C1(_19893_),
    .X(_21953_));
 sky130_fd_sc_hd__or2_2 _50842_ (.A(_21952_),
    .B(_21953_),
    .X(_21954_));
 sky130_fd_sc_hd__a31o_1 _50843_ (.A1(_19929_),
    .A2(_19081_),
    .A3(_03414_),
    .B1(_19928_),
    .X(_21955_));
 sky130_fd_sc_hd__clkbuf_2 _50844_ (.A(_13449_),
    .X(_21956_));
 sky130_fd_sc_hd__and2b_1 _50845_ (.A_N(_13680_),
    .B(\delay_line[5][8] ),
    .X(_21957_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _50846_ (.A(\delay_line[5][8] ),
    .X(_21958_));
 sky130_fd_sc_hd__and2b_1 _50847_ (.A_N(_21958_),
    .B(_13680_),
    .X(_21959_));
 sky130_fd_sc_hd__o21ai_2 _50848_ (.A1(_21957_),
    .A2(_21959_),
    .B1(_19927_),
    .Y(_21960_));
 sky130_fd_sc_hd__or2b_1 _50849_ (.A(_13680_),
    .B_N(_21958_),
    .X(_21961_));
 sky130_fd_sc_hd__inv_2 _50850_ (.A(\delay_line[5][8] ),
    .Y(_21962_));
 sky130_fd_sc_hd__nand2_1 _50851_ (.A(_21962_),
    .B(_09437_),
    .Y(_21963_));
 sky130_fd_sc_hd__nand3_2 _50852_ (.A(_21961_),
    .B(_21963_),
    .C(\delay_line[5][7] ),
    .Y(_21964_));
 sky130_fd_sc_hd__a22o_1 _50853_ (.A1(_21956_),
    .A2(_19081_),
    .B1(_21960_),
    .B2(_21964_),
    .X(_21965_));
 sky130_fd_sc_hd__nand4_1 _50854_ (.A(_21960_),
    .B(_21964_),
    .C(_21956_),
    .D(_18095_),
    .Y(_21966_));
 sky130_fd_sc_hd__nand3b_1 _50855_ (.A_N(_21955_),
    .B(_21965_),
    .C(_21966_),
    .Y(_21967_));
 sky130_fd_sc_hd__a21oi_2 _50856_ (.A1(_21960_),
    .A2(_21964_),
    .B1(_19902_),
    .Y(_21968_));
 sky130_fd_sc_hd__and3_1 _50857_ (.A(_21960_),
    .B(_21964_),
    .C(_19902_),
    .X(_21969_));
 sky130_fd_sc_hd__o21ai_2 _50858_ (.A1(_21968_),
    .A2(_21969_),
    .B1(_21955_),
    .Y(_21970_));
 sky130_fd_sc_hd__clkbuf_2 _50859_ (.A(\delay_line[3][8] ),
    .X(_21971_));
 sky130_fd_sc_hd__xnor2_1 _50860_ (.A(_03546_),
    .B(_21971_),
    .Y(_21972_));
 sky130_fd_sc_hd__xor2_1 _50861_ (.A(_19921_),
    .B(_21972_),
    .X(_21973_));
 sky130_fd_sc_hd__nand3_1 _50862_ (.A(_21967_),
    .B(_21970_),
    .C(_21973_),
    .Y(_21974_));
 sky130_fd_sc_hd__a21o_1 _50863_ (.A1(_21967_),
    .A2(_21970_),
    .B1(_21973_),
    .X(_21975_));
 sky130_fd_sc_hd__nand2_1 _50864_ (.A(_21974_),
    .B(_21975_),
    .Y(_21976_));
 sky130_fd_sc_hd__nand2_1 _50865_ (.A(_19906_),
    .B(_19911_),
    .Y(_21977_));
 sky130_fd_sc_hd__clkbuf_2 _50866_ (.A(net428),
    .X(_21978_));
 sky130_fd_sc_hd__clkbuf_2 _50867_ (.A(_19904_),
    .X(_21979_));
 sky130_fd_sc_hd__nand3b_2 _50868_ (.A_N(_21978_),
    .B(_21979_),
    .C(_18082_),
    .Y(_21980_));
 sky130_fd_sc_hd__or2b_1 _50869_ (.A(\delay_line[6][6] ),
    .B_N(_18080_),
    .X(_21981_));
 sky130_fd_sc_hd__or2b_1 _50870_ (.A(net429),
    .B_N(_21978_),
    .X(_21982_));
 sky130_fd_sc_hd__nand3_1 _50871_ (.A(_19905_),
    .B(_21981_),
    .C(_21982_),
    .Y(_21983_));
 sky130_fd_sc_hd__a21o_1 _50872_ (.A1(_21980_),
    .A2(_21983_),
    .B1(_21956_),
    .X(_21984_));
 sky130_fd_sc_hd__nand3_2 _50873_ (.A(_21983_),
    .B(_21956_),
    .C(_21980_),
    .Y(_21985_));
 sky130_fd_sc_hd__nand4_4 _50874_ (.A(_21984_),
    .B(_21906_),
    .C(_03458_),
    .D(_21985_),
    .Y(_21986_));
 sky130_fd_sc_hd__o2bb2ai_1 _50875_ (.A1_N(_21985_),
    .A2_N(_21984_),
    .B1(_00073_),
    .B2(_03238_),
    .Y(_21987_));
 sky130_fd_sc_hd__nand3_2 _50876_ (.A(_21977_),
    .B(_21986_),
    .C(_21987_),
    .Y(_21988_));
 sky130_fd_sc_hd__a21o_1 _50877_ (.A1(_21986_),
    .A2(_21987_),
    .B1(_21977_),
    .X(_21989_));
 sky130_fd_sc_hd__o21a_1 _50878_ (.A1(_03425_),
    .A2(_19081_),
    .B1(_19916_),
    .X(_21990_));
 sky130_fd_sc_hd__a32o_1 _50879_ (.A1(_18078_),
    .A2(_19909_),
    .A3(_19911_),
    .B1(_19915_),
    .B2(_21990_),
    .X(_21991_));
 sky130_fd_sc_hd__a21o_1 _50880_ (.A1(_21988_),
    .A2(_21989_),
    .B1(_21991_),
    .X(_21992_));
 sky130_fd_sc_hd__nand3_2 _50881_ (.A(_21991_),
    .B(_21988_),
    .C(_21989_),
    .Y(_21993_));
 sky130_fd_sc_hd__nand3b_2 _50882_ (.A_N(_21976_),
    .B(_21992_),
    .C(_21993_),
    .Y(_21994_));
 sky130_fd_sc_hd__a22o_1 _50883_ (.A1(_21993_),
    .A2(_21992_),
    .B1(_21974_),
    .B2(_21975_),
    .X(_21995_));
 sky130_fd_sc_hd__o221a_1 _50884_ (.A1(_03425_),
    .A2(_19081_),
    .B1(_19064_),
    .B2(_19066_),
    .C1(_24820_),
    .X(_21996_));
 sky130_fd_sc_hd__a32o_1 _50885_ (.A1(_19912_),
    .A2(_19915_),
    .A3(_21996_),
    .B1(_19939_),
    .B2(_19938_),
    .X(_21997_));
 sky130_fd_sc_hd__a21o_1 _50886_ (.A1(_21994_),
    .A2(_21995_),
    .B1(_21997_),
    .X(_21998_));
 sky130_fd_sc_hd__nand3_2 _50887_ (.A(_21997_),
    .B(_21994_),
    .C(_21995_),
    .Y(_21999_));
 sky130_fd_sc_hd__nand2_2 _50888_ (.A(_21998_),
    .B(_21999_),
    .Y(_22000_));
 sky130_fd_sc_hd__xor2_2 _50889_ (.A(_21954_),
    .B(_22000_),
    .X(_22001_));
 sky130_fd_sc_hd__a21o_1 _50890_ (.A1(_21935_),
    .A2(_21937_),
    .B1(_22001_),
    .X(_22002_));
 sky130_fd_sc_hd__nand3_1 _50891_ (.A(_21937_),
    .B(_22001_),
    .C(_21935_),
    .Y(_22003_));
 sky130_fd_sc_hd__nand2_1 _50892_ (.A(_20148_),
    .B(_20151_),
    .Y(_22004_));
 sky130_fd_sc_hd__a21oi_4 _50893_ (.A1(_22002_),
    .A2(_22003_),
    .B1(_22004_),
    .Y(_22005_));
 sky130_fd_sc_hd__dfxtp_1 _50894_ (.CLK(clk),
    .D(_00000_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _50895_ (.CLK(clk),
    .D(_00001_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _50896_ (.CLK(clk),
    .D(_00002_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _50897_ (.CLK(clk),
    .D(_00003_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _50898_ (.CLK(clk),
    .D(_00035_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _50899_ (.CLK(clk),
    .D(_00036_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _50900_ (.CLK(clk),
    .D(_00037_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _50901_ (.CLK(clk),
    .D(_00038_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _50902_ (.CLK(clk),
    .D(_00039_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _50903_ (.CLK(clk),
    .D(_00040_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _50904_ (.CLK(clk),
    .D(_00004_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _50905_ (.CLK(clk),
    .D(_00005_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _50906_ (.CLK(clk),
    .D(_00006_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _50907_ (.CLK(clk),
    .D(_00007_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _50908_ (.CLK(clk),
    .D(_00008_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _50909_ (.CLK(clk),
    .D(_00009_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _50910_ (.CLK(clk),
    .D(_00010_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _50911_ (.CLK(clk),
    .D(_00011_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _50912_ (.CLK(clk),
    .D(_00012_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _50913_ (.CLK(clk),
    .D(_00013_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _50914_ (.CLK(clk),
    .D(_00014_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _50915_ (.CLK(clk),
    .D(_00015_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _50916_ (.CLK(clk),
    .D(_00016_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_2 _50917_ (.CLK(clk),
    .D(_00017_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _50918_ (.CLK(clk),
    .D(_00018_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_2 _50919_ (.CLK(clk),
    .D(_00019_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_2 _50920_ (.CLK(clk),
    .D(_00020_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_2 _50921_ (.CLK(clk),
    .D(_00021_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_2 _50922_ (.CLK(clk),
    .D(_00022_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_2 _50923_ (.CLK(clk),
    .D(_00023_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _50924_ (.CLK(clk),
    .D(_00024_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_2 _50925_ (.CLK(clk),
    .D(_00025_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_2 _50926_ (.CLK(clk),
    .D(_00026_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_2 _50927_ (.CLK(clk),
    .D(_00027_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _50928_ (.CLK(clk),
    .D(_00028_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _50929_ (.CLK(clk),
    .D(_00029_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _50930_ (.CLK(clk),
    .D(_00030_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _50931_ (.CLK(clk),
    .D(_00031_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _50932_ (.CLK(clk),
    .D(_00032_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _50933_ (.CLK(clk),
    .D(_00033_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _50934_ (.CLK(clk),
    .D(_00034_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_2 _50935_ (.CLK(clk),
    .D(net1),
    .Q(\delay_line[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _50936_ (.CLK(clk),
    .D(net8),
    .Q(\delay_line[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _50937_ (.CLK(clk),
    .D(net9),
    .Q(\delay_line[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _50938_ (.CLK(clk),
    .D(net10),
    .Q(\delay_line[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _50939_ (.CLK(clk),
    .D(net11),
    .Q(\delay_line[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _50940_ (.CLK(clk),
    .D(net12),
    .Q(\delay_line[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _50941_ (.CLK(clk),
    .D(net13),
    .Q(\delay_line[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _50942_ (.CLK(clk),
    .D(net14),
    .Q(\delay_line[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _50943_ (.CLK(clk),
    .D(net15),
    .Q(\delay_line[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _50944_ (.CLK(clk),
    .D(net16),
    .Q(\delay_line[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _50945_ (.CLK(clk),
    .D(net2),
    .Q(\delay_line[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _50946_ (.CLK(clk),
    .D(net3),
    .Q(\delay_line[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _50947_ (.CLK(clk),
    .D(net4),
    .Q(\delay_line[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _50948_ (.CLK(clk),
    .D(net5),
    .Q(\delay_line[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _50949_ (.CLK(clk),
    .D(net6),
    .Q(\delay_line[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _50950_ (.CLK(clk),
    .D(net7),
    .Q(\delay_line[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _50951_ (.CLK(clk),
    .D(\delay_line[0][0] ),
    .Q(\delay_line[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _50952_ (.CLK(clk),
    .D(\delay_line[0][1] ),
    .Q(\delay_line[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _50953_ (.CLK(clk),
    .D(\delay_line[0][2] ),
    .Q(\delay_line[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _50954_ (.CLK(clk),
    .D(\delay_line[0][3] ),
    .Q(\delay_line[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _50955_ (.CLK(clk),
    .D(\delay_line[0][4] ),
    .Q(\delay_line[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _50956_ (.CLK(clk),
    .D(\delay_line[0][5] ),
    .Q(\delay_line[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _50957_ (.CLK(clk),
    .D(\delay_line[0][6] ),
    .Q(\delay_line[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _50958_ (.CLK(clk),
    .D(\delay_line[0][7] ),
    .Q(\delay_line[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _50959_ (.CLK(clk),
    .D(net455),
    .Q(\delay_line[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _50960_ (.CLK(clk),
    .D(\delay_line[0][9] ),
    .Q(\delay_line[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _50961_ (.CLK(clk),
    .D(\delay_line[0][10] ),
    .Q(\delay_line[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _50962_ (.CLK(clk),
    .D(\delay_line[0][11] ),
    .Q(\delay_line[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _50963_ (.CLK(clk),
    .D(net454),
    .Q(\delay_line[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _50964_ (.CLK(clk),
    .D(\delay_line[0][13] ),
    .Q(\delay_line[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _50965_ (.CLK(clk),
    .D(\delay_line[0][14] ),
    .Q(\delay_line[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _50966_ (.CLK(clk),
    .D(\delay_line[0][15] ),
    .Q(\delay_line[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _50967_ (.CLK(clk),
    .D(\delay_line[1][0] ),
    .Q(\delay_line[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _50968_ (.CLK(clk),
    .D(\delay_line[1][1] ),
    .Q(\delay_line[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _50969_ (.CLK(clk),
    .D(\delay_line[1][2] ),
    .Q(\delay_line[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _50970_ (.CLK(clk),
    .D(\delay_line[1][3] ),
    .Q(\delay_line[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _50971_ (.CLK(clk),
    .D(\delay_line[1][4] ),
    .Q(\delay_line[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _50972_ (.CLK(clk),
    .D(\delay_line[1][5] ),
    .Q(\delay_line[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _50973_ (.CLK(clk),
    .D(\delay_line[1][6] ),
    .Q(\delay_line[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _50974_ (.CLK(clk),
    .D(\delay_line[1][7] ),
    .Q(\delay_line[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _50975_ (.CLK(clk),
    .D(net450),
    .Q(\delay_line[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _50976_ (.CLK(clk),
    .D(\delay_line[1][9] ),
    .Q(\delay_line[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _50977_ (.CLK(clk),
    .D(net449),
    .Q(\delay_line[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _50978_ (.CLK(clk),
    .D(\delay_line[1][11] ),
    .Q(\delay_line[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _50979_ (.CLK(clk),
    .D(\delay_line[1][12] ),
    .Q(\delay_line[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _50980_ (.CLK(clk),
    .D(net447),
    .Q(\delay_line[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _50981_ (.CLK(clk),
    .D(net446),
    .Q(\delay_line[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _50982_ (.CLK(clk),
    .D(net445),
    .Q(\delay_line[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _50983_ (.CLK(clk),
    .D(\delay_line[2][0] ),
    .Q(\delay_line[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _50984_ (.CLK(clk),
    .D(\delay_line[2][1] ),
    .Q(\delay_line[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _50985_ (.CLK(clk),
    .D(\delay_line[2][2] ),
    .Q(\delay_line[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _50986_ (.CLK(clk),
    .D(\delay_line[2][3] ),
    .Q(\delay_line[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _50987_ (.CLK(clk),
    .D(net444),
    .Q(\delay_line[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _50988_ (.CLK(clk),
    .D(net443),
    .Q(\delay_line[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _50989_ (.CLK(clk),
    .D(\delay_line[2][6] ),
    .Q(\delay_line[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _50990_ (.CLK(clk),
    .D(\delay_line[2][7] ),
    .Q(\delay_line[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _50991_ (.CLK(clk),
    .D(\delay_line[2][8] ),
    .Q(\delay_line[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _50992_ (.CLK(clk),
    .D(\delay_line[2][9] ),
    .Q(\delay_line[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _50993_ (.CLK(clk),
    .D(\delay_line[2][10] ),
    .Q(\delay_line[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _50994_ (.CLK(clk),
    .D(\delay_line[2][11] ),
    .Q(\delay_line[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _50995_ (.CLK(clk),
    .D(\delay_line[2][12] ),
    .Q(\delay_line[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _50996_ (.CLK(clk),
    .D(\delay_line[2][13] ),
    .Q(\delay_line[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _50997_ (.CLK(clk),
    .D(\delay_line[2][14] ),
    .Q(\delay_line[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _50998_ (.CLK(clk),
    .D(\delay_line[2][15] ),
    .Q(\delay_line[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _50999_ (.CLK(clk),
    .D(\delay_line[3][0] ),
    .Q(\delay_line[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _51000_ (.CLK(clk),
    .D(\delay_line[3][1] ),
    .Q(\delay_line[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _51001_ (.CLK(clk),
    .D(\delay_line[3][2] ),
    .Q(\delay_line[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51002_ (.CLK(clk),
    .D(\delay_line[3][3] ),
    .Q(\delay_line[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51003_ (.CLK(clk),
    .D(\delay_line[3][4] ),
    .Q(\delay_line[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51004_ (.CLK(clk),
    .D(\delay_line[3][5] ),
    .Q(\delay_line[4][5] ));
 sky130_fd_sc_hd__dfxtp_4 _51005_ (.CLK(clk),
    .D(\delay_line[3][6] ),
    .Q(\delay_line[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _51006_ (.CLK(clk),
    .D(\delay_line[3][7] ),
    .Q(\delay_line[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _51007_ (.CLK(clk),
    .D(\delay_line[3][8] ),
    .Q(\delay_line[4][8] ));
 sky130_fd_sc_hd__dfxtp_4 _51008_ (.CLK(clk),
    .D(\delay_line[3][9] ),
    .Q(\delay_line[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51009_ (.CLK(clk),
    .D(\delay_line[3][10] ),
    .Q(\delay_line[4][10] ));
 sky130_fd_sc_hd__dfxtp_4 _51010_ (.CLK(clk),
    .D(\delay_line[3][11] ),
    .Q(\delay_line[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51011_ (.CLK(clk),
    .D(\delay_line[3][12] ),
    .Q(\delay_line[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _51012_ (.CLK(clk),
    .D(\delay_line[3][13] ),
    .Q(\delay_line[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _51013_ (.CLK(clk),
    .D(net435),
    .Q(\delay_line[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _51014_ (.CLK(clk),
    .D(\delay_line[3][15] ),
    .Q(\delay_line[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _51015_ (.CLK(clk),
    .D(\delay_line[4][0] ),
    .Q(\delay_line[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51016_ (.CLK(clk),
    .D(\delay_line[4][1] ),
    .Q(\delay_line[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51017_ (.CLK(clk),
    .D(\delay_line[4][2] ),
    .Q(\delay_line[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51018_ (.CLK(clk),
    .D(\delay_line[4][3] ),
    .Q(\delay_line[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _51019_ (.CLK(clk),
    .D(net434),
    .Q(\delay_line[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51020_ (.CLK(clk),
    .D(\delay_line[4][5] ),
    .Q(\delay_line[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51021_ (.CLK(clk),
    .D(\delay_line[4][6] ),
    .Q(\delay_line[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51022_ (.CLK(clk),
    .D(\delay_line[4][7] ),
    .Q(\delay_line[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51023_ (.CLK(clk),
    .D(\delay_line[4][8] ),
    .Q(\delay_line[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _51024_ (.CLK(clk),
    .D(\delay_line[4][9] ),
    .Q(\delay_line[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51025_ (.CLK(clk),
    .D(\delay_line[4][10] ),
    .Q(\delay_line[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51026_ (.CLK(clk),
    .D(\delay_line[4][11] ),
    .Q(\delay_line[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51027_ (.CLK(clk),
    .D(net433),
    .Q(\delay_line[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51028_ (.CLK(clk),
    .D(\delay_line[4][13] ),
    .Q(\delay_line[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51029_ (.CLK(clk),
    .D(net432),
    .Q(\delay_line[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51030_ (.CLK(clk),
    .D(\delay_line[4][15] ),
    .Q(\delay_line[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51031_ (.CLK(clk),
    .D(\delay_line[5][0] ),
    .Q(\delay_line[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51032_ (.CLK(clk),
    .D(\delay_line[5][1] ),
    .Q(\delay_line[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51033_ (.CLK(clk),
    .D(\delay_line[5][2] ),
    .Q(\delay_line[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51034_ (.CLK(clk),
    .D(\delay_line[5][3] ),
    .Q(\delay_line[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51035_ (.CLK(clk),
    .D(\delay_line[5][4] ),
    .Q(\delay_line[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51036_ (.CLK(clk),
    .D(\delay_line[5][5] ),
    .Q(\delay_line[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51037_ (.CLK(clk),
    .D(\delay_line[5][6] ),
    .Q(\delay_line[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51038_ (.CLK(clk),
    .D(\delay_line[5][7] ),
    .Q(\delay_line[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51039_ (.CLK(clk),
    .D(\delay_line[5][8] ),
    .Q(\delay_line[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51040_ (.CLK(clk),
    .D(\delay_line[5][9] ),
    .Q(\delay_line[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51041_ (.CLK(clk),
    .D(net430),
    .Q(\delay_line[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51042_ (.CLK(clk),
    .D(\delay_line[5][11] ),
    .Q(\delay_line[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51043_ (.CLK(clk),
    .D(\delay_line[5][12] ),
    .Q(\delay_line[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51044_ (.CLK(clk),
    .D(\delay_line[5][13] ),
    .Q(\delay_line[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51045_ (.CLK(clk),
    .D(\delay_line[5][14] ),
    .Q(\delay_line[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51046_ (.CLK(clk),
    .D(\delay_line[5][15] ),
    .Q(\delay_line[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51047_ (.CLK(clk),
    .D(\delay_line[6][0] ),
    .Q(\delay_line[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51048_ (.CLK(clk),
    .D(\delay_line[6][1] ),
    .Q(\delay_line[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51049_ (.CLK(clk),
    .D(\delay_line[6][2] ),
    .Q(\delay_line[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51050_ (.CLK(clk),
    .D(\delay_line[6][3] ),
    .Q(\delay_line[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51051_ (.CLK(clk),
    .D(\delay_line[6][4] ),
    .Q(\delay_line[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51052_ (.CLK(clk),
    .D(\delay_line[6][5] ),
    .Q(\delay_line[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51053_ (.CLK(clk),
    .D(net428),
    .Q(\delay_line[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51054_ (.CLK(clk),
    .D(\delay_line[6][7] ),
    .Q(\delay_line[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51055_ (.CLK(clk),
    .D(\delay_line[6][8] ),
    .Q(\delay_line[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51056_ (.CLK(clk),
    .D(\delay_line[6][9] ),
    .Q(\delay_line[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51057_ (.CLK(clk),
    .D(\delay_line[6][10] ),
    .Q(\delay_line[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51058_ (.CLK(clk),
    .D(\delay_line[6][11] ),
    .Q(\delay_line[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51059_ (.CLK(clk),
    .D(\delay_line[6][12] ),
    .Q(\delay_line[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51060_ (.CLK(clk),
    .D(\delay_line[6][13] ),
    .Q(\delay_line[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51061_ (.CLK(clk),
    .D(\delay_line[6][14] ),
    .Q(\delay_line[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51062_ (.CLK(clk),
    .D(\delay_line[6][15] ),
    .Q(\delay_line[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51063_ (.CLK(clk),
    .D(\delay_line[7][0] ),
    .Q(\delay_line[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51064_ (.CLK(clk),
    .D(\delay_line[7][1] ),
    .Q(\delay_line[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51065_ (.CLK(clk),
    .D(\delay_line[7][2] ),
    .Q(\delay_line[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51066_ (.CLK(clk),
    .D(\delay_line[7][3] ),
    .Q(\delay_line[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51067_ (.CLK(clk),
    .D(\delay_line[7][4] ),
    .Q(\delay_line[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51068_ (.CLK(clk),
    .D(\delay_line[7][5] ),
    .Q(\delay_line[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51069_ (.CLK(clk),
    .D(\delay_line[7][6] ),
    .Q(\delay_line[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51070_ (.CLK(clk),
    .D(\delay_line[7][7] ),
    .Q(\delay_line[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51071_ (.CLK(clk),
    .D(\delay_line[7][8] ),
    .Q(\delay_line[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51072_ (.CLK(clk),
    .D(net425),
    .Q(\delay_line[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51073_ (.CLK(clk),
    .D(\delay_line[7][10] ),
    .Q(\delay_line[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51074_ (.CLK(clk),
    .D(\delay_line[7][11] ),
    .Q(\delay_line[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51075_ (.CLK(clk),
    .D(\delay_line[7][12] ),
    .Q(\delay_line[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51076_ (.CLK(clk),
    .D(\delay_line[7][13] ),
    .Q(\delay_line[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51077_ (.CLK(clk),
    .D(\delay_line[7][14] ),
    .Q(\delay_line[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51078_ (.CLK(clk),
    .D(\delay_line[7][15] ),
    .Q(\delay_line[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51079_ (.CLK(clk),
    .D(\delay_line[8][0] ),
    .Q(\delay_line[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _51080_ (.CLK(clk),
    .D(\delay_line[8][1] ),
    .Q(\delay_line[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51081_ (.CLK(clk),
    .D(\delay_line[8][2] ),
    .Q(\delay_line[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51082_ (.CLK(clk),
    .D(\delay_line[8][3] ),
    .Q(\delay_line[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51083_ (.CLK(clk),
    .D(\delay_line[8][4] ),
    .Q(\delay_line[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51084_ (.CLK(clk),
    .D(\delay_line[8][5] ),
    .Q(\delay_line[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51085_ (.CLK(clk),
    .D(\delay_line[8][6] ),
    .Q(\delay_line[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51086_ (.CLK(clk),
    .D(\delay_line[8][7] ),
    .Q(\delay_line[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51087_ (.CLK(clk),
    .D(net424),
    .Q(\delay_line[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51088_ (.CLK(clk),
    .D(\delay_line[8][9] ),
    .Q(\delay_line[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51089_ (.CLK(clk),
    .D(\delay_line[8][10] ),
    .Q(\delay_line[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51090_ (.CLK(clk),
    .D(\delay_line[8][11] ),
    .Q(\delay_line[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51091_ (.CLK(clk),
    .D(\delay_line[8][12] ),
    .Q(\delay_line[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51092_ (.CLK(clk),
    .D(\delay_line[8][13] ),
    .Q(\delay_line[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51093_ (.CLK(clk),
    .D(net423),
    .Q(\delay_line[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51094_ (.CLK(clk),
    .D(\delay_line[8][15] ),
    .Q(\delay_line[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51095_ (.CLK(clk),
    .D(\delay_line[9][0] ),
    .Q(\delay_line[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51096_ (.CLK(clk),
    .D(\delay_line[9][1] ),
    .Q(\delay_line[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51097_ (.CLK(clk),
    .D(\delay_line[9][2] ),
    .Q(\delay_line[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51098_ (.CLK(clk),
    .D(\delay_line[9][3] ),
    .Q(\delay_line[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51099_ (.CLK(clk),
    .D(\delay_line[9][4] ),
    .Q(\delay_line[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51100_ (.CLK(clk),
    .D(\delay_line[9][5] ),
    .Q(\delay_line[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51101_ (.CLK(clk),
    .D(net421),
    .Q(\delay_line[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51102_ (.CLK(clk),
    .D(\delay_line[9][7] ),
    .Q(\delay_line[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51103_ (.CLK(clk),
    .D(\delay_line[9][8] ),
    .Q(\delay_line[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51104_ (.CLK(clk),
    .D(\delay_line[9][9] ),
    .Q(\delay_line[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51105_ (.CLK(clk),
    .D(\delay_line[9][10] ),
    .Q(\delay_line[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51106_ (.CLK(clk),
    .D(\delay_line[9][11] ),
    .Q(\delay_line[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51107_ (.CLK(clk),
    .D(net417),
    .Q(\delay_line[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51108_ (.CLK(clk),
    .D(net416),
    .Q(\delay_line[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51109_ (.CLK(clk),
    .D(\delay_line[9][14] ),
    .Q(\delay_line[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51110_ (.CLK(clk),
    .D(\delay_line[9][15] ),
    .Q(\delay_line[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _51111_ (.CLK(clk),
    .D(net415),
    .Q(\delay_line[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51112_ (.CLK(clk),
    .D(\delay_line[10][1] ),
    .Q(\delay_line[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51113_ (.CLK(clk),
    .D(\delay_line[10][2] ),
    .Q(\delay_line[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51114_ (.CLK(clk),
    .D(\delay_line[10][3] ),
    .Q(\delay_line[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51115_ (.CLK(clk),
    .D(net413),
    .Q(\delay_line[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51116_ (.CLK(clk),
    .D(\delay_line[10][5] ),
    .Q(\delay_line[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51117_ (.CLK(clk),
    .D(\delay_line[10][6] ),
    .Q(\delay_line[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51118_ (.CLK(clk),
    .D(net412),
    .Q(\delay_line[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51119_ (.CLK(clk),
    .D(\delay_line[10][8] ),
    .Q(\delay_line[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51120_ (.CLK(clk),
    .D(\delay_line[10][9] ),
    .Q(\delay_line[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51121_ (.CLK(clk),
    .D(\delay_line[10][10] ),
    .Q(\delay_line[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51122_ (.CLK(clk),
    .D(\delay_line[10][11] ),
    .Q(\delay_line[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51123_ (.CLK(clk),
    .D(\delay_line[10][12] ),
    .Q(\delay_line[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _51124_ (.CLK(clk),
    .D(net411),
    .Q(\delay_line[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51125_ (.CLK(clk),
    .D(\delay_line[10][14] ),
    .Q(\delay_line[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51126_ (.CLK(clk),
    .D(\delay_line[10][15] ),
    .Q(\delay_line[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51127_ (.CLK(clk),
    .D(\delay_line[11][0] ),
    .Q(\delay_line[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51128_ (.CLK(clk),
    .D(\delay_line[11][1] ),
    .Q(\delay_line[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _51129_ (.CLK(clk),
    .D(\delay_line[11][2] ),
    .Q(\delay_line[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51130_ (.CLK(clk),
    .D(\delay_line[11][3] ),
    .Q(\delay_line[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _51131_ (.CLK(clk),
    .D(\delay_line[11][4] ),
    .Q(\delay_line[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51132_ (.CLK(clk),
    .D(\delay_line[11][5] ),
    .Q(\delay_line[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51133_ (.CLK(clk),
    .D(\delay_line[11][6] ),
    .Q(\delay_line[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51134_ (.CLK(clk),
    .D(\delay_line[11][7] ),
    .Q(\delay_line[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51135_ (.CLK(clk),
    .D(\delay_line[11][8] ),
    .Q(\delay_line[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51136_ (.CLK(clk),
    .D(\delay_line[11][9] ),
    .Q(\delay_line[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51137_ (.CLK(clk),
    .D(\delay_line[11][10] ),
    .Q(\delay_line[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51138_ (.CLK(clk),
    .D(net410),
    .Q(\delay_line[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51139_ (.CLK(clk),
    .D(\delay_line[11][12] ),
    .Q(\delay_line[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51140_ (.CLK(clk),
    .D(\delay_line[11][13] ),
    .Q(\delay_line[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51141_ (.CLK(clk),
    .D(net409),
    .Q(\delay_line[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51142_ (.CLK(clk),
    .D(net408),
    .Q(\delay_line[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51143_ (.CLK(clk),
    .D(\delay_line[12][0] ),
    .Q(\delay_line[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _51144_ (.CLK(clk),
    .D(\delay_line[12][1] ),
    .Q(\delay_line[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51145_ (.CLK(clk),
    .D(\delay_line[12][2] ),
    .Q(\delay_line[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51146_ (.CLK(clk),
    .D(net407),
    .Q(\delay_line[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51147_ (.CLK(clk),
    .D(\delay_line[12][4] ),
    .Q(\delay_line[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51148_ (.CLK(clk),
    .D(net406),
    .Q(\delay_line[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51149_ (.CLK(clk),
    .D(\delay_line[12][6] ),
    .Q(\delay_line[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51150_ (.CLK(clk),
    .D(net405),
    .Q(\delay_line[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51151_ (.CLK(clk),
    .D(\delay_line[12][8] ),
    .Q(\delay_line[13][8] ));
 sky130_fd_sc_hd__dfxtp_4 _51152_ (.CLK(clk),
    .D(net403),
    .Q(\delay_line[13][9] ));
 sky130_fd_sc_hd__dfxtp_4 _51153_ (.CLK(clk),
    .D(\delay_line[12][10] ),
    .Q(\delay_line[13][10] ));
 sky130_fd_sc_hd__dfxtp_4 _51154_ (.CLK(clk),
    .D(\delay_line[12][11] ),
    .Q(\delay_line[13][11] ));
 sky130_fd_sc_hd__dfxtp_4 _51155_ (.CLK(clk),
    .D(net402),
    .Q(\delay_line[13][12] ));
 sky130_fd_sc_hd__dfxtp_4 _51156_ (.CLK(clk),
    .D(net401),
    .Q(\delay_line[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51157_ (.CLK(clk),
    .D(net400),
    .Q(\delay_line[13][14] ));
 sky130_fd_sc_hd__dfxtp_4 _51158_ (.CLK(clk),
    .D(net399),
    .Q(\delay_line[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51159_ (.CLK(clk),
    .D(net398),
    .Q(\delay_line[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51160_ (.CLK(clk),
    .D(\delay_line[13][1] ),
    .Q(\delay_line[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _51161_ (.CLK(clk),
    .D(\delay_line[13][2] ),
    .Q(\delay_line[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51162_ (.CLK(clk),
    .D(\delay_line[13][3] ),
    .Q(\delay_line[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _51163_ (.CLK(clk),
    .D(\delay_line[13][4] ),
    .Q(\delay_line[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51164_ (.CLK(clk),
    .D(net397),
    .Q(\delay_line[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51165_ (.CLK(clk),
    .D(\delay_line[13][6] ),
    .Q(\delay_line[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _51166_ (.CLK(clk),
    .D(\delay_line[13][7] ),
    .Q(\delay_line[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51167_ (.CLK(clk),
    .D(net396),
    .Q(\delay_line[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _51168_ (.CLK(clk),
    .D(\delay_line[13][9] ),
    .Q(\delay_line[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51169_ (.CLK(clk),
    .D(\delay_line[13][10] ),
    .Q(\delay_line[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _51170_ (.CLK(clk),
    .D(\delay_line[13][11] ),
    .Q(\delay_line[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51171_ (.CLK(clk),
    .D(\delay_line[13][12] ),
    .Q(\delay_line[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _51172_ (.CLK(clk),
    .D(\delay_line[13][13] ),
    .Q(\delay_line[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51173_ (.CLK(clk),
    .D(net395),
    .Q(\delay_line[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51174_ (.CLK(clk),
    .D(\delay_line[13][15] ),
    .Q(\delay_line[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51175_ (.CLK(clk),
    .D(net394),
    .Q(\delay_line[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _51176_ (.CLK(clk),
    .D(net393),
    .Q(\delay_line[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51177_ (.CLK(clk),
    .D(\delay_line[14][2] ),
    .Q(\delay_line[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51178_ (.CLK(clk),
    .D(net392),
    .Q(\delay_line[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51179_ (.CLK(clk),
    .D(\delay_line[14][4] ),
    .Q(\delay_line[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51180_ (.CLK(clk),
    .D(net391),
    .Q(\delay_line[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51181_ (.CLK(clk),
    .D(\delay_line[14][6] ),
    .Q(\delay_line[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51182_ (.CLK(clk),
    .D(\delay_line[14][7] ),
    .Q(\delay_line[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51183_ (.CLK(clk),
    .D(net390),
    .Q(\delay_line[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51184_ (.CLK(clk),
    .D(\delay_line[14][9] ),
    .Q(\delay_line[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51185_ (.CLK(clk),
    .D(\delay_line[14][10] ),
    .Q(\delay_line[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51186_ (.CLK(clk),
    .D(\delay_line[14][11] ),
    .Q(\delay_line[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51187_ (.CLK(clk),
    .D(\delay_line[14][12] ),
    .Q(\delay_line[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51188_ (.CLK(clk),
    .D(\delay_line[14][13] ),
    .Q(\delay_line[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51189_ (.CLK(clk),
    .D(net389),
    .Q(\delay_line[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51190_ (.CLK(clk),
    .D(net388),
    .Q(\delay_line[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51191_ (.CLK(clk),
    .D(\delay_line[15][0] ),
    .Q(\delay_line[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51192_ (.CLK(clk),
    .D(\delay_line[15][1] ),
    .Q(\delay_line[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51193_ (.CLK(clk),
    .D(\delay_line[15][2] ),
    .Q(\delay_line[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51194_ (.CLK(clk),
    .D(\delay_line[15][3] ),
    .Q(\delay_line[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51195_ (.CLK(clk),
    .D(net387),
    .Q(\delay_line[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51196_ (.CLK(clk),
    .D(\delay_line[15][5] ),
    .Q(\delay_line[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51197_ (.CLK(clk),
    .D(\delay_line[15][6] ),
    .Q(\delay_line[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51198_ (.CLK(clk),
    .D(\delay_line[15][7] ),
    .Q(\delay_line[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51199_ (.CLK(clk),
    .D(\delay_line[15][8] ),
    .Q(\delay_line[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51200_ (.CLK(clk),
    .D(net386),
    .Q(\delay_line[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51201_ (.CLK(clk),
    .D(\delay_line[15][10] ),
    .Q(\delay_line[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51202_ (.CLK(clk),
    .D(\delay_line[15][11] ),
    .Q(\delay_line[16][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51203_ (.CLK(clk),
    .D(\delay_line[15][12] ),
    .Q(\delay_line[16][12] ));
 sky130_fd_sc_hd__dfxtp_2 _51204_ (.CLK(clk),
    .D(\delay_line[15][13] ),
    .Q(\delay_line[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51205_ (.CLK(clk),
    .D(\delay_line[15][14] ),
    .Q(\delay_line[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51206_ (.CLK(clk),
    .D(\delay_line[15][15] ),
    .Q(\delay_line[16][15] ));
 sky130_fd_sc_hd__dfxtp_2 _51207_ (.CLK(clk),
    .D(\delay_line[16][0] ),
    .Q(\delay_line[17][0] ));
 sky130_fd_sc_hd__dfxtp_4 _51208_ (.CLK(clk),
    .D(\delay_line[16][1] ),
    .Q(\delay_line[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _51209_ (.CLK(clk),
    .D(\delay_line[16][2] ),
    .Q(\delay_line[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51210_ (.CLK(clk),
    .D(\delay_line[16][3] ),
    .Q(\delay_line[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _51211_ (.CLK(clk),
    .D(\delay_line[16][4] ),
    .Q(\delay_line[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51212_ (.CLK(clk),
    .D(\delay_line[16][5] ),
    .Q(\delay_line[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51213_ (.CLK(clk),
    .D(net385),
    .Q(\delay_line[17][6] ));
 sky130_fd_sc_hd__dfxtp_4 _51214_ (.CLK(clk),
    .D(net384),
    .Q(\delay_line[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 _51215_ (.CLK(clk),
    .D(net383),
    .Q(\delay_line[17][8] ));
 sky130_fd_sc_hd__dfxtp_2 _51216_ (.CLK(clk),
    .D(\delay_line[16][9] ),
    .Q(\delay_line[17][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51217_ (.CLK(clk),
    .D(net382),
    .Q(\delay_line[17][10] ));
 sky130_fd_sc_hd__dfxtp_2 _51218_ (.CLK(clk),
    .D(net381),
    .Q(\delay_line[17][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51219_ (.CLK(clk),
    .D(\delay_line[16][12] ),
    .Q(\delay_line[17][12] ));
 sky130_fd_sc_hd__dfxtp_2 _51220_ (.CLK(clk),
    .D(\delay_line[16][13] ),
    .Q(\delay_line[17][13] ));
 sky130_fd_sc_hd__dfxtp_2 _51221_ (.CLK(clk),
    .D(net380),
    .Q(\delay_line[17][14] ));
 sky130_fd_sc_hd__dfxtp_2 _51222_ (.CLK(clk),
    .D(net379),
    .Q(\delay_line[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51223_ (.CLK(clk),
    .D(net378),
    .Q(\delay_line[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51224_ (.CLK(clk),
    .D(\delay_line[17][1] ),
    .Q(\delay_line[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51225_ (.CLK(clk),
    .D(\delay_line[17][2] ),
    .Q(\delay_line[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51226_ (.CLK(clk),
    .D(\delay_line[17][3] ),
    .Q(\delay_line[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51227_ (.CLK(clk),
    .D(\delay_line[17][4] ),
    .Q(\delay_line[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51228_ (.CLK(clk),
    .D(\delay_line[17][5] ),
    .Q(\delay_line[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51229_ (.CLK(clk),
    .D(\delay_line[17][6] ),
    .Q(\delay_line[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51230_ (.CLK(clk),
    .D(\delay_line[17][7] ),
    .Q(\delay_line[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51231_ (.CLK(clk),
    .D(net377),
    .Q(\delay_line[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51232_ (.CLK(clk),
    .D(net376),
    .Q(\delay_line[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51233_ (.CLK(clk),
    .D(\delay_line[17][10] ),
    .Q(\delay_line[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51234_ (.CLK(clk),
    .D(\delay_line[17][11] ),
    .Q(\delay_line[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51235_ (.CLK(clk),
    .D(\delay_line[17][12] ),
    .Q(\delay_line[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51236_ (.CLK(clk),
    .D(\delay_line[17][13] ),
    .Q(\delay_line[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51237_ (.CLK(clk),
    .D(\delay_line[17][14] ),
    .Q(\delay_line[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51238_ (.CLK(clk),
    .D(\delay_line[17][15] ),
    .Q(\delay_line[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51239_ (.CLK(clk),
    .D(\delay_line[18][0] ),
    .Q(\delay_line[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51240_ (.CLK(clk),
    .D(net375),
    .Q(\delay_line[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51241_ (.CLK(clk),
    .D(\delay_line[18][2] ),
    .Q(\delay_line[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51242_ (.CLK(clk),
    .D(\delay_line[18][3] ),
    .Q(\delay_line[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51243_ (.CLK(clk),
    .D(\delay_line[18][4] ),
    .Q(\delay_line[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51244_ (.CLK(clk),
    .D(\delay_line[18][5] ),
    .Q(\delay_line[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51245_ (.CLK(clk),
    .D(\delay_line[18][6] ),
    .Q(\delay_line[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51246_ (.CLK(clk),
    .D(\delay_line[18][7] ),
    .Q(\delay_line[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51247_ (.CLK(clk),
    .D(\delay_line[18][8] ),
    .Q(\delay_line[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51248_ (.CLK(clk),
    .D(\delay_line[18][9] ),
    .Q(\delay_line[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51249_ (.CLK(clk),
    .D(net373),
    .Q(\delay_line[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51250_ (.CLK(clk),
    .D(\delay_line[18][11] ),
    .Q(\delay_line[19][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51251_ (.CLK(clk),
    .D(\delay_line[18][12] ),
    .Q(\delay_line[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51252_ (.CLK(clk),
    .D(\delay_line[18][13] ),
    .Q(\delay_line[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51253_ (.CLK(clk),
    .D(\delay_line[18][14] ),
    .Q(\delay_line[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51254_ (.CLK(clk),
    .D(net372),
    .Q(\delay_line[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51255_ (.CLK(clk),
    .D(\delay_line[19][0] ),
    .Q(\delay_line[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51256_ (.CLK(clk),
    .D(\delay_line[19][1] ),
    .Q(\delay_line[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51257_ (.CLK(clk),
    .D(\delay_line[19][2] ),
    .Q(\delay_line[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51258_ (.CLK(clk),
    .D(\delay_line[19][3] ),
    .Q(\delay_line[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51259_ (.CLK(clk),
    .D(net371),
    .Q(\delay_line[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51260_ (.CLK(clk),
    .D(\delay_line[19][5] ),
    .Q(\delay_line[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51261_ (.CLK(clk),
    .D(\delay_line[19][6] ),
    .Q(\delay_line[20][6] ));
 sky130_fd_sc_hd__dfxtp_2 _51262_ (.CLK(clk),
    .D(net370),
    .Q(\delay_line[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51263_ (.CLK(clk),
    .D(\delay_line[19][8] ),
    .Q(\delay_line[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51264_ (.CLK(clk),
    .D(\delay_line[19][9] ),
    .Q(\delay_line[20][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51265_ (.CLK(clk),
    .D(\delay_line[19][10] ),
    .Q(\delay_line[20][10] ));
 sky130_fd_sc_hd__dfxtp_2 _51266_ (.CLK(clk),
    .D(\delay_line[19][11] ),
    .Q(\delay_line[20][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51267_ (.CLK(clk),
    .D(\delay_line[19][12] ),
    .Q(\delay_line[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51268_ (.CLK(clk),
    .D(\delay_line[19][13] ),
    .Q(\delay_line[20][13] ));
 sky130_fd_sc_hd__dfxtp_2 _51269_ (.CLK(clk),
    .D(\delay_line[19][14] ),
    .Q(\delay_line[20][14] ));
 sky130_fd_sc_hd__dfxtp_2 _51270_ (.CLK(clk),
    .D(\delay_line[19][15] ),
    .Q(\delay_line[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51271_ (.CLK(clk),
    .D(\delay_line[20][0] ),
    .Q(\delay_line[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51272_ (.CLK(clk),
    .D(net368),
    .Q(\delay_line[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51273_ (.CLK(clk),
    .D(net367),
    .Q(\delay_line[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51274_ (.CLK(clk),
    .D(\delay_line[20][3] ),
    .Q(\delay_line[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51275_ (.CLK(clk),
    .D(\delay_line[20][4] ),
    .Q(\delay_line[21][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51276_ (.CLK(clk),
    .D(net366),
    .Q(\delay_line[21][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51277_ (.CLK(clk),
    .D(\delay_line[20][6] ),
    .Q(\delay_line[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51278_ (.CLK(clk),
    .D(\delay_line[20][7] ),
    .Q(\delay_line[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51279_ (.CLK(clk),
    .D(\delay_line[20][8] ),
    .Q(\delay_line[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51280_ (.CLK(clk),
    .D(\delay_line[20][9] ),
    .Q(\delay_line[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51281_ (.CLK(clk),
    .D(\delay_line[20][10] ),
    .Q(\delay_line[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51282_ (.CLK(clk),
    .D(\delay_line[20][11] ),
    .Q(\delay_line[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51283_ (.CLK(clk),
    .D(\delay_line[20][12] ),
    .Q(\delay_line[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51284_ (.CLK(clk),
    .D(net364),
    .Q(\delay_line[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51285_ (.CLK(clk),
    .D(net363),
    .Q(\delay_line[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51286_ (.CLK(clk),
    .D(net362),
    .Q(\delay_line[21][15] ));
 sky130_fd_sc_hd__dfxtp_2 _51287_ (.CLK(clk),
    .D(\delay_line[21][0] ),
    .Q(\delay_line[22][0] ));
 sky130_fd_sc_hd__dfxtp_2 _51288_ (.CLK(clk),
    .D(\delay_line[21][1] ),
    .Q(\delay_line[22][1] ));
 sky130_fd_sc_hd__dfxtp_2 _51289_ (.CLK(clk),
    .D(\delay_line[21][2] ),
    .Q(\delay_line[22][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51290_ (.CLK(clk),
    .D(\delay_line[21][3] ),
    .Q(\delay_line[22][3] ));
 sky130_fd_sc_hd__dfxtp_2 _51291_ (.CLK(clk),
    .D(\delay_line[21][4] ),
    .Q(\delay_line[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51292_ (.CLK(clk),
    .D(\delay_line[21][5] ),
    .Q(\delay_line[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51293_ (.CLK(clk),
    .D(\delay_line[21][6] ),
    .Q(\delay_line[22][6] ));
 sky130_fd_sc_hd__dfxtp_2 _51294_ (.CLK(clk),
    .D(\delay_line[21][7] ),
    .Q(\delay_line[22][7] ));
 sky130_fd_sc_hd__dfxtp_2 _51295_ (.CLK(clk),
    .D(net359),
    .Q(\delay_line[22][8] ));
 sky130_fd_sc_hd__dfxtp_2 _51296_ (.CLK(clk),
    .D(\delay_line[21][9] ),
    .Q(\delay_line[22][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51297_ (.CLK(clk),
    .D(\delay_line[21][10] ),
    .Q(\delay_line[22][10] ));
 sky130_fd_sc_hd__dfxtp_2 _51298_ (.CLK(clk),
    .D(\delay_line[21][11] ),
    .Q(\delay_line[22][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51299_ (.CLK(clk),
    .D(net357),
    .Q(\delay_line[22][12] ));
 sky130_fd_sc_hd__dfxtp_2 _51300_ (.CLK(clk),
    .D(\delay_line[21][13] ),
    .Q(\delay_line[22][13] ));
 sky130_fd_sc_hd__dfxtp_2 _51301_ (.CLK(clk),
    .D(\delay_line[21][14] ),
    .Q(\delay_line[22][14] ));
 sky130_fd_sc_hd__dfxtp_2 _51302_ (.CLK(clk),
    .D(\delay_line[21][15] ),
    .Q(\delay_line[22][15] ));
 sky130_fd_sc_hd__dfxtp_2 _51303_ (.CLK(clk),
    .D(\delay_line[22][0] ),
    .Q(\delay_line[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51304_ (.CLK(clk),
    .D(net356),
    .Q(\delay_line[23][1] ));
 sky130_fd_sc_hd__dfxtp_2 _51305_ (.CLK(clk),
    .D(net355),
    .Q(\delay_line[23][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51306_ (.CLK(clk),
    .D(net354),
    .Q(\delay_line[23][3] ));
 sky130_fd_sc_hd__dfxtp_2 _51307_ (.CLK(clk),
    .D(\delay_line[22][4] ),
    .Q(\delay_line[23][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51308_ (.CLK(clk),
    .D(net353),
    .Q(\delay_line[23][5] ));
 sky130_fd_sc_hd__dfxtp_4 _51309_ (.CLK(clk),
    .D(\delay_line[22][6] ),
    .Q(\delay_line[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51310_ (.CLK(clk),
    .D(net352),
    .Q(\delay_line[23][7] ));
 sky130_fd_sc_hd__dfxtp_2 _51311_ (.CLK(clk),
    .D(\delay_line[22][8] ),
    .Q(\delay_line[23][8] ));
 sky130_fd_sc_hd__dfxtp_2 _51312_ (.CLK(clk),
    .D(\delay_line[22][9] ),
    .Q(\delay_line[23][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51313_ (.CLK(clk),
    .D(\delay_line[22][10] ),
    .Q(\delay_line[23][10] ));
 sky130_fd_sc_hd__dfxtp_4 _51314_ (.CLK(clk),
    .D(\delay_line[22][11] ),
    .Q(\delay_line[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51315_ (.CLK(clk),
    .D(\delay_line[22][12] ),
    .Q(\delay_line[23][12] ));
 sky130_fd_sc_hd__dfxtp_2 _51316_ (.CLK(clk),
    .D(\delay_line[22][13] ),
    .Q(\delay_line[23][13] ));
 sky130_fd_sc_hd__dfxtp_4 _51317_ (.CLK(clk),
    .D(net351),
    .Q(\delay_line[23][14] ));
 sky130_fd_sc_hd__dfxtp_2 _51318_ (.CLK(clk),
    .D(net350),
    .Q(\delay_line[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51319_ (.CLK(clk),
    .D(\delay_line[23][0] ),
    .Q(\delay_line[24][0] ));
 sky130_fd_sc_hd__dfxtp_2 _51320_ (.CLK(clk),
    .D(\delay_line[23][1] ),
    .Q(\delay_line[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51321_ (.CLK(clk),
    .D(\delay_line[23][2] ),
    .Q(\delay_line[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51322_ (.CLK(clk),
    .D(\delay_line[23][3] ),
    .Q(\delay_line[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51323_ (.CLK(clk),
    .D(\delay_line[23][4] ),
    .Q(\delay_line[24][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51324_ (.CLK(clk),
    .D(\delay_line[23][5] ),
    .Q(\delay_line[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51325_ (.CLK(clk),
    .D(\delay_line[23][6] ),
    .Q(\delay_line[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51326_ (.CLK(clk),
    .D(net349),
    .Q(\delay_line[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51327_ (.CLK(clk),
    .D(\delay_line[23][8] ),
    .Q(\delay_line[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51328_ (.CLK(clk),
    .D(\delay_line[23][9] ),
    .Q(\delay_line[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51329_ (.CLK(clk),
    .D(\delay_line[23][10] ),
    .Q(\delay_line[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51330_ (.CLK(clk),
    .D(\delay_line[23][11] ),
    .Q(\delay_line[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51331_ (.CLK(clk),
    .D(net347),
    .Q(\delay_line[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51332_ (.CLK(clk),
    .D(\delay_line[23][13] ),
    .Q(\delay_line[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51333_ (.CLK(clk),
    .D(\delay_line[23][14] ),
    .Q(\delay_line[24][14] ));
 sky130_fd_sc_hd__dfxtp_2 _51334_ (.CLK(clk),
    .D(\delay_line[23][15] ),
    .Q(\delay_line[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51335_ (.CLK(clk),
    .D(\delay_line[24][0] ),
    .Q(\delay_line[25][0] ));
 sky130_fd_sc_hd__dfxtp_2 _51336_ (.CLK(clk),
    .D(net345),
    .Q(\delay_line[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51337_ (.CLK(clk),
    .D(net344),
    .Q(\delay_line[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51338_ (.CLK(clk),
    .D(\delay_line[24][3] ),
    .Q(\delay_line[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51339_ (.CLK(clk),
    .D(net343),
    .Q(\delay_line[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51340_ (.CLK(clk),
    .D(\delay_line[24][5] ),
    .Q(\delay_line[25][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51341_ (.CLK(clk),
    .D(\delay_line[24][6] ),
    .Q(\delay_line[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51342_ (.CLK(clk),
    .D(\delay_line[24][7] ),
    .Q(\delay_line[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51343_ (.CLK(clk),
    .D(net342),
    .Q(\delay_line[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51344_ (.CLK(clk),
    .D(\delay_line[24][9] ),
    .Q(\delay_line[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51345_ (.CLK(clk),
    .D(\delay_line[24][10] ),
    .Q(\delay_line[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51346_ (.CLK(clk),
    .D(\delay_line[24][11] ),
    .Q(\delay_line[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51347_ (.CLK(clk),
    .D(\delay_line[24][12] ),
    .Q(\delay_line[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51348_ (.CLK(clk),
    .D(\delay_line[24][13] ),
    .Q(\delay_line[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51349_ (.CLK(clk),
    .D(\delay_line[24][14] ),
    .Q(\delay_line[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51350_ (.CLK(clk),
    .D(\delay_line[24][15] ),
    .Q(\delay_line[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51351_ (.CLK(clk),
    .D(\delay_line[25][0] ),
    .Q(\delay_line[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51352_ (.CLK(clk),
    .D(\delay_line[25][1] ),
    .Q(\delay_line[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51353_ (.CLK(clk),
    .D(\delay_line[25][2] ),
    .Q(\delay_line[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51354_ (.CLK(clk),
    .D(\delay_line[25][3] ),
    .Q(\delay_line[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51355_ (.CLK(clk),
    .D(\delay_line[25][4] ),
    .Q(\delay_line[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51356_ (.CLK(clk),
    .D(\delay_line[25][5] ),
    .Q(\delay_line[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51357_ (.CLK(clk),
    .D(\delay_line[25][6] ),
    .Q(\delay_line[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51358_ (.CLK(clk),
    .D(\delay_line[25][7] ),
    .Q(\delay_line[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51359_ (.CLK(clk),
    .D(\delay_line[25][8] ),
    .Q(\delay_line[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51360_ (.CLK(clk),
    .D(\delay_line[25][9] ),
    .Q(\delay_line[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51361_ (.CLK(clk),
    .D(\delay_line[25][10] ),
    .Q(\delay_line[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51362_ (.CLK(clk),
    .D(\delay_line[25][11] ),
    .Q(\delay_line[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51363_ (.CLK(clk),
    .D(\delay_line[25][12] ),
    .Q(\delay_line[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51364_ (.CLK(clk),
    .D(\delay_line[25][13] ),
    .Q(\delay_line[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51365_ (.CLK(clk),
    .D(\delay_line[25][14] ),
    .Q(\delay_line[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51366_ (.CLK(clk),
    .D(\delay_line[25][15] ),
    .Q(\delay_line[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51367_ (.CLK(clk),
    .D(\delay_line[26][0] ),
    .Q(\delay_line[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51368_ (.CLK(clk),
    .D(\delay_line[26][1] ),
    .Q(\delay_line[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51369_ (.CLK(clk),
    .D(\delay_line[26][2] ),
    .Q(\delay_line[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51370_ (.CLK(clk),
    .D(\delay_line[26][3] ),
    .Q(\delay_line[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51371_ (.CLK(clk),
    .D(\delay_line[26][4] ),
    .Q(\delay_line[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51372_ (.CLK(clk),
    .D(\delay_line[26][5] ),
    .Q(\delay_line[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51373_ (.CLK(clk),
    .D(\delay_line[26][6] ),
    .Q(\delay_line[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51374_ (.CLK(clk),
    .D(\delay_line[26][7] ),
    .Q(\delay_line[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51375_ (.CLK(clk),
    .D(\delay_line[26][8] ),
    .Q(\delay_line[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51376_ (.CLK(clk),
    .D(\delay_line[26][9] ),
    .Q(\delay_line[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51377_ (.CLK(clk),
    .D(\delay_line[26][10] ),
    .Q(\delay_line[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51378_ (.CLK(clk),
    .D(\delay_line[26][11] ),
    .Q(\delay_line[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51379_ (.CLK(clk),
    .D(\delay_line[26][12] ),
    .Q(\delay_line[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51380_ (.CLK(clk),
    .D(\delay_line[26][13] ),
    .Q(\delay_line[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51381_ (.CLK(clk),
    .D(\delay_line[26][14] ),
    .Q(\delay_line[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51382_ (.CLK(clk),
    .D(\delay_line[26][15] ),
    .Q(\delay_line[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51383_ (.CLK(clk),
    .D(\delay_line[27][0] ),
    .Q(\delay_line[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51384_ (.CLK(clk),
    .D(\delay_line[27][1] ),
    .Q(\delay_line[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51385_ (.CLK(clk),
    .D(\delay_line[27][2] ),
    .Q(\delay_line[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51386_ (.CLK(clk),
    .D(\delay_line[27][3] ),
    .Q(\delay_line[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51387_ (.CLK(clk),
    .D(\delay_line[27][4] ),
    .Q(\delay_line[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51388_ (.CLK(clk),
    .D(net333),
    .Q(\delay_line[28][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51389_ (.CLK(clk),
    .D(net332),
    .Q(\delay_line[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51390_ (.CLK(clk),
    .D(\delay_line[27][7] ),
    .Q(\delay_line[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51391_ (.CLK(clk),
    .D(\delay_line[27][8] ),
    .Q(\delay_line[28][8] ));
 sky130_fd_sc_hd__dfxtp_2 _51392_ (.CLK(clk),
    .D(net331),
    .Q(\delay_line[28][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51393_ (.CLK(clk),
    .D(\delay_line[27][10] ),
    .Q(\delay_line[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51394_ (.CLK(clk),
    .D(net330),
    .Q(\delay_line[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51395_ (.CLK(clk),
    .D(\delay_line[27][12] ),
    .Q(\delay_line[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51396_ (.CLK(clk),
    .D(\delay_line[27][13] ),
    .Q(\delay_line[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51397_ (.CLK(clk),
    .D(\delay_line[27][14] ),
    .Q(\delay_line[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51398_ (.CLK(clk),
    .D(\delay_line[27][15] ),
    .Q(\delay_line[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51399_ (.CLK(clk),
    .D(\delay_line[28][0] ),
    .Q(\delay_line[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51400_ (.CLK(clk),
    .D(\delay_line[28][1] ),
    .Q(\delay_line[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51401_ (.CLK(clk),
    .D(\delay_line[28][2] ),
    .Q(\delay_line[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51402_ (.CLK(clk),
    .D(net328),
    .Q(\delay_line[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51403_ (.CLK(clk),
    .D(net327),
    .Q(\delay_line[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51404_ (.CLK(clk),
    .D(\delay_line[28][5] ),
    .Q(\delay_line[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51405_ (.CLK(clk),
    .D(\delay_line[28][6] ),
    .Q(\delay_line[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51406_ (.CLK(clk),
    .D(\delay_line[28][7] ),
    .Q(\delay_line[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51407_ (.CLK(clk),
    .D(\delay_line[28][8] ),
    .Q(\delay_line[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51408_ (.CLK(clk),
    .D(\delay_line[28][9] ),
    .Q(\delay_line[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51409_ (.CLK(clk),
    .D(\delay_line[28][10] ),
    .Q(\delay_line[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51410_ (.CLK(clk),
    .D(net326),
    .Q(\delay_line[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51411_ (.CLK(clk),
    .D(net325),
    .Q(\delay_line[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51412_ (.CLK(clk),
    .D(net324),
    .Q(\delay_line[29][13] ));
 sky130_fd_sc_hd__dfxtp_2 _51413_ (.CLK(clk),
    .D(\delay_line[28][14] ),
    .Q(\delay_line[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51414_ (.CLK(clk),
    .D(\delay_line[28][15] ),
    .Q(\delay_line[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51415_ (.CLK(clk),
    .D(\delay_line[29][0] ),
    .Q(\delay_line[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51416_ (.CLK(clk),
    .D(\delay_line[29][1] ),
    .Q(\delay_line[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51417_ (.CLK(clk),
    .D(\delay_line[29][2] ),
    .Q(\delay_line[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51418_ (.CLK(clk),
    .D(\delay_line[29][3] ),
    .Q(\delay_line[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51419_ (.CLK(clk),
    .D(\delay_line[29][4] ),
    .Q(\delay_line[30][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51420_ (.CLK(clk),
    .D(\delay_line[29][5] ),
    .Q(\delay_line[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51421_ (.CLK(clk),
    .D(\delay_line[29][6] ),
    .Q(\delay_line[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51422_ (.CLK(clk),
    .D(\delay_line[29][7] ),
    .Q(\delay_line[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51423_ (.CLK(clk),
    .D(net322),
    .Q(\delay_line[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51424_ (.CLK(clk),
    .D(net321),
    .Q(\delay_line[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51425_ (.CLK(clk),
    .D(\delay_line[29][10] ),
    .Q(\delay_line[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51426_ (.CLK(clk),
    .D(\delay_line[29][11] ),
    .Q(\delay_line[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51427_ (.CLK(clk),
    .D(\delay_line[29][12] ),
    .Q(\delay_line[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51428_ (.CLK(clk),
    .D(\delay_line[29][13] ),
    .Q(\delay_line[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51429_ (.CLK(clk),
    .D(\delay_line[29][14] ),
    .Q(\delay_line[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51430_ (.CLK(clk),
    .D(\delay_line[29][15] ),
    .Q(\delay_line[30][15] ));
 sky130_fd_sc_hd__dfxtp_4 _51431_ (.CLK(clk),
    .D(\delay_line[30][0] ),
    .Q(\delay_line[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51432_ (.CLK(clk),
    .D(net320),
    .Q(\delay_line[31][1] ));
 sky130_fd_sc_hd__dfxtp_4 _51433_ (.CLK(clk),
    .D(\delay_line[30][2] ),
    .Q(\delay_line[31][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51434_ (.CLK(clk),
    .D(\delay_line[30][3] ),
    .Q(\delay_line[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51435_ (.CLK(clk),
    .D(\delay_line[30][4] ),
    .Q(\delay_line[31][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51436_ (.CLK(clk),
    .D(\delay_line[30][5] ),
    .Q(\delay_line[31][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51437_ (.CLK(clk),
    .D(\delay_line[30][6] ),
    .Q(\delay_line[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51438_ (.CLK(clk),
    .D(\delay_line[30][7] ),
    .Q(\delay_line[31][7] ));
 sky130_fd_sc_hd__dfxtp_2 _51439_ (.CLK(clk),
    .D(\delay_line[30][8] ),
    .Q(\delay_line[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51440_ (.CLK(clk),
    .D(\delay_line[30][9] ),
    .Q(\delay_line[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51441_ (.CLK(clk),
    .D(\delay_line[30][10] ),
    .Q(\delay_line[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51442_ (.CLK(clk),
    .D(\delay_line[30][11] ),
    .Q(\delay_line[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51443_ (.CLK(clk),
    .D(\delay_line[30][12] ),
    .Q(\delay_line[31][12] ));
 sky130_fd_sc_hd__dfxtp_2 _51444_ (.CLK(clk),
    .D(\delay_line[30][13] ),
    .Q(\delay_line[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51445_ (.CLK(clk),
    .D(\delay_line[30][14] ),
    .Q(\delay_line[31][14] ));
 sky130_fd_sc_hd__dfxtp_2 _51446_ (.CLK(clk),
    .D(net319),
    .Q(\delay_line[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51447_ (.CLK(clk),
    .D(\delay_line[31][0] ),
    .Q(\delay_line[32][0] ));
 sky130_fd_sc_hd__dfxtp_2 _51448_ (.CLK(clk),
    .D(\delay_line[31][1] ),
    .Q(\delay_line[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51449_ (.CLK(clk),
    .D(\delay_line[31][2] ),
    .Q(\delay_line[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51450_ (.CLK(clk),
    .D(\delay_line[31][3] ),
    .Q(\delay_line[32][3] ));
 sky130_fd_sc_hd__dfxtp_2 _51451_ (.CLK(clk),
    .D(net318),
    .Q(\delay_line[32][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51452_ (.CLK(clk),
    .D(\delay_line[31][5] ),
    .Q(\delay_line[32][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51453_ (.CLK(clk),
    .D(\delay_line[31][6] ),
    .Q(\delay_line[32][6] ));
 sky130_fd_sc_hd__dfxtp_2 _51454_ (.CLK(clk),
    .D(net317),
    .Q(\delay_line[32][7] ));
 sky130_fd_sc_hd__dfxtp_2 _51455_ (.CLK(clk),
    .D(\delay_line[31][8] ),
    .Q(\delay_line[32][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51456_ (.CLK(clk),
    .D(\delay_line[31][9] ),
    .Q(\delay_line[32][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51457_ (.CLK(clk),
    .D(\delay_line[31][10] ),
    .Q(\delay_line[32][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51458_ (.CLK(clk),
    .D(net316),
    .Q(\delay_line[32][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51459_ (.CLK(clk),
    .D(\delay_line[31][12] ),
    .Q(\delay_line[32][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51460_ (.CLK(clk),
    .D(\delay_line[31][13] ),
    .Q(\delay_line[32][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51461_ (.CLK(clk),
    .D(\delay_line[31][14] ),
    .Q(\delay_line[32][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51462_ (.CLK(clk),
    .D(\delay_line[31][15] ),
    .Q(\delay_line[32][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51463_ (.CLK(clk),
    .D(\delay_line[32][0] ),
    .Q(\delay_line[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51464_ (.CLK(clk),
    .D(\delay_line[32][1] ),
    .Q(\delay_line[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51465_ (.CLK(clk),
    .D(\delay_line[32][2] ),
    .Q(\delay_line[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51466_ (.CLK(clk),
    .D(\delay_line[32][3] ),
    .Q(\delay_line[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51467_ (.CLK(clk),
    .D(\delay_line[32][4] ),
    .Q(\delay_line[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51468_ (.CLK(clk),
    .D(\delay_line[32][5] ),
    .Q(\delay_line[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51469_ (.CLK(clk),
    .D(\delay_line[32][6] ),
    .Q(\delay_line[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51470_ (.CLK(clk),
    .D(\delay_line[32][7] ),
    .Q(\delay_line[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51471_ (.CLK(clk),
    .D(\delay_line[32][8] ),
    .Q(\delay_line[33][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51472_ (.CLK(clk),
    .D(\delay_line[32][9] ),
    .Q(\delay_line[33][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51473_ (.CLK(clk),
    .D(\delay_line[32][10] ),
    .Q(\delay_line[33][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51474_ (.CLK(clk),
    .D(\delay_line[32][11] ),
    .Q(\delay_line[33][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51475_ (.CLK(clk),
    .D(\delay_line[32][12] ),
    .Q(\delay_line[33][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51476_ (.CLK(clk),
    .D(\delay_line[32][13] ),
    .Q(\delay_line[33][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51477_ (.CLK(clk),
    .D(\delay_line[32][14] ),
    .Q(\delay_line[33][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51478_ (.CLK(clk),
    .D(\delay_line[32][15] ),
    .Q(\delay_line[33][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51479_ (.CLK(clk),
    .D(net315),
    .Q(\delay_line[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51480_ (.CLK(clk),
    .D(\delay_line[33][1] ),
    .Q(\delay_line[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51481_ (.CLK(clk),
    .D(net314),
    .Q(\delay_line[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51482_ (.CLK(clk),
    .D(net313),
    .Q(\delay_line[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51483_ (.CLK(clk),
    .D(\delay_line[33][4] ),
    .Q(\delay_line[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51484_ (.CLK(clk),
    .D(net312),
    .Q(\delay_line[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51485_ (.CLK(clk),
    .D(\delay_line[33][6] ),
    .Q(\delay_line[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51486_ (.CLK(clk),
    .D(\delay_line[33][7] ),
    .Q(\delay_line[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51487_ (.CLK(clk),
    .D(\delay_line[33][8] ),
    .Q(\delay_line[34][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51488_ (.CLK(clk),
    .D(\delay_line[33][9] ),
    .Q(\delay_line[34][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51489_ (.CLK(clk),
    .D(\delay_line[33][10] ),
    .Q(\delay_line[34][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51490_ (.CLK(clk),
    .D(\delay_line[33][11] ),
    .Q(\delay_line[34][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51491_ (.CLK(clk),
    .D(\delay_line[33][12] ),
    .Q(\delay_line[34][12] ));
 sky130_fd_sc_hd__dfxtp_4 _51492_ (.CLK(clk),
    .D(net311),
    .Q(\delay_line[34][13] ));
 sky130_fd_sc_hd__dfxtp_2 _51493_ (.CLK(clk),
    .D(net310),
    .Q(\delay_line[34][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51494_ (.CLK(clk),
    .D(\delay_line[33][15] ),
    .Q(\delay_line[34][15] ));
 sky130_fd_sc_hd__dfxtp_2 _51495_ (.CLK(clk),
    .D(\delay_line[34][0] ),
    .Q(\delay_line[35][0] ));
 sky130_fd_sc_hd__dfxtp_4 _51496_ (.CLK(clk),
    .D(\delay_line[34][1] ),
    .Q(\delay_line[35][1] ));
 sky130_fd_sc_hd__dfxtp_2 _51497_ (.CLK(clk),
    .D(net307),
    .Q(\delay_line[35][2] ));
 sky130_fd_sc_hd__dfxtp_2 _51498_ (.CLK(clk),
    .D(\delay_line[34][3] ),
    .Q(\delay_line[35][3] ));
 sky130_fd_sc_hd__dfxtp_2 _51499_ (.CLK(clk),
    .D(\delay_line[34][4] ),
    .Q(\delay_line[35][4] ));
 sky130_fd_sc_hd__dfxtp_2 _51500_ (.CLK(clk),
    .D(\delay_line[34][5] ),
    .Q(\delay_line[35][5] ));
 sky130_fd_sc_hd__dfxtp_2 _51501_ (.CLK(clk),
    .D(\delay_line[34][6] ),
    .Q(\delay_line[35][6] ));
 sky130_fd_sc_hd__dfxtp_2 _51502_ (.CLK(clk),
    .D(\delay_line[34][7] ),
    .Q(\delay_line[35][7] ));
 sky130_fd_sc_hd__dfxtp_2 _51503_ (.CLK(clk),
    .D(\delay_line[34][8] ),
    .Q(\delay_line[35][8] ));
 sky130_fd_sc_hd__dfxtp_2 _51504_ (.CLK(clk),
    .D(\delay_line[34][9] ),
    .Q(\delay_line[35][9] ));
 sky130_fd_sc_hd__dfxtp_2 _51505_ (.CLK(clk),
    .D(\delay_line[34][10] ),
    .Q(\delay_line[35][10] ));
 sky130_fd_sc_hd__dfxtp_2 _51506_ (.CLK(clk),
    .D(\delay_line[34][11] ),
    .Q(\delay_line[35][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51507_ (.CLK(clk),
    .D(\delay_line[34][12] ),
    .Q(\delay_line[35][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51508_ (.CLK(clk),
    .D(\delay_line[34][13] ),
    .Q(\delay_line[35][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51509_ (.CLK(clk),
    .D(\delay_line[34][14] ),
    .Q(\delay_line[35][14] ));
 sky130_fd_sc_hd__dfxtp_2 _51510_ (.CLK(clk),
    .D(\delay_line[34][15] ),
    .Q(\delay_line[35][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51511_ (.CLK(clk),
    .D(\delay_line[35][0] ),
    .Q(\delay_line[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51512_ (.CLK(clk),
    .D(\delay_line[35][1] ),
    .Q(\delay_line[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51513_ (.CLK(clk),
    .D(\delay_line[35][2] ),
    .Q(\delay_line[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51514_ (.CLK(clk),
    .D(\delay_line[35][3] ),
    .Q(\delay_line[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51515_ (.CLK(clk),
    .D(\delay_line[35][4] ),
    .Q(\delay_line[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51516_ (.CLK(clk),
    .D(\delay_line[35][5] ),
    .Q(\delay_line[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51517_ (.CLK(clk),
    .D(\delay_line[35][6] ),
    .Q(\delay_line[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51518_ (.CLK(clk),
    .D(\delay_line[35][7] ),
    .Q(\delay_line[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51519_ (.CLK(clk),
    .D(\delay_line[35][8] ),
    .Q(\delay_line[36][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51520_ (.CLK(clk),
    .D(\delay_line[35][9] ),
    .Q(\delay_line[36][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51521_ (.CLK(clk),
    .D(\delay_line[35][10] ),
    .Q(\delay_line[36][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51522_ (.CLK(clk),
    .D(\delay_line[35][11] ),
    .Q(\delay_line[36][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51523_ (.CLK(clk),
    .D(net301),
    .Q(\delay_line[36][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51524_ (.CLK(clk),
    .D(net300),
    .Q(\delay_line[36][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51525_ (.CLK(clk),
    .D(\delay_line[35][14] ),
    .Q(\delay_line[36][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51526_ (.CLK(clk),
    .D(\delay_line[35][15] ),
    .Q(\delay_line[36][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51527_ (.CLK(clk),
    .D(\delay_line[36][0] ),
    .Q(\delay_line[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51528_ (.CLK(clk),
    .D(net298),
    .Q(\delay_line[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51529_ (.CLK(clk),
    .D(\delay_line[36][2] ),
    .Q(\delay_line[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51530_ (.CLK(clk),
    .D(\delay_line[36][3] ),
    .Q(\delay_line[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51531_ (.CLK(clk),
    .D(\delay_line[36][4] ),
    .Q(\delay_line[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51532_ (.CLK(clk),
    .D(\delay_line[36][5] ),
    .Q(\delay_line[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51533_ (.CLK(clk),
    .D(\delay_line[36][6] ),
    .Q(\delay_line[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51534_ (.CLK(clk),
    .D(net297),
    .Q(\delay_line[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51535_ (.CLK(clk),
    .D(\delay_line[36][8] ),
    .Q(\delay_line[37][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51536_ (.CLK(clk),
    .D(net296),
    .Q(\delay_line[37][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51537_ (.CLK(clk),
    .D(\delay_line[36][10] ),
    .Q(\delay_line[37][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51538_ (.CLK(clk),
    .D(\delay_line[36][11] ),
    .Q(\delay_line[37][11] ));
 sky130_fd_sc_hd__dfxtp_2 _51539_ (.CLK(clk),
    .D(\delay_line[36][12] ),
    .Q(\delay_line[37][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51540_ (.CLK(clk),
    .D(\delay_line[36][13] ),
    .Q(\delay_line[37][13] ));
 sky130_fd_sc_hd__dfxtp_2 _51541_ (.CLK(clk),
    .D(net295),
    .Q(\delay_line[37][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51542_ (.CLK(clk),
    .D(net294),
    .Q(\delay_line[37][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51543_ (.CLK(clk),
    .D(\delay_line[37][0] ),
    .Q(\delay_line[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51544_ (.CLK(clk),
    .D(net293),
    .Q(\delay_line[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51545_ (.CLK(clk),
    .D(\delay_line[37][2] ),
    .Q(\delay_line[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51546_ (.CLK(clk),
    .D(\delay_line[37][3] ),
    .Q(\delay_line[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51547_ (.CLK(clk),
    .D(\delay_line[37][4] ),
    .Q(\delay_line[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51548_ (.CLK(clk),
    .D(\delay_line[37][5] ),
    .Q(\delay_line[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51549_ (.CLK(clk),
    .D(\delay_line[37][6] ),
    .Q(\delay_line[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51550_ (.CLK(clk),
    .D(net292),
    .Q(\delay_line[38][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51551_ (.CLK(clk),
    .D(\delay_line[37][8] ),
    .Q(\delay_line[38][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51552_ (.CLK(clk),
    .D(\delay_line[37][9] ),
    .Q(\delay_line[38][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51553_ (.CLK(clk),
    .D(\delay_line[37][10] ),
    .Q(\delay_line[38][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51554_ (.CLK(clk),
    .D(\delay_line[37][11] ),
    .Q(\delay_line[38][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51555_ (.CLK(clk),
    .D(\delay_line[37][12] ),
    .Q(\delay_line[38][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51556_ (.CLK(clk),
    .D(\delay_line[37][13] ),
    .Q(\delay_line[38][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51557_ (.CLK(clk),
    .D(\delay_line[37][14] ),
    .Q(\delay_line[38][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51558_ (.CLK(clk),
    .D(net291),
    .Q(\delay_line[38][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51559_ (.CLK(clk),
    .D(\delay_line[38][0] ),
    .Q(\delay_line[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51560_ (.CLK(clk),
    .D(\delay_line[38][1] ),
    .Q(\delay_line[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51561_ (.CLK(clk),
    .D(\delay_line[38][2] ),
    .Q(\delay_line[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51562_ (.CLK(clk),
    .D(net289),
    .Q(\delay_line[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51563_ (.CLK(clk),
    .D(net288),
    .Q(\delay_line[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51564_ (.CLK(clk),
    .D(\delay_line[38][5] ),
    .Q(\delay_line[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51565_ (.CLK(clk),
    .D(\delay_line[38][6] ),
    .Q(\delay_line[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51566_ (.CLK(clk),
    .D(\delay_line[38][7] ),
    .Q(\delay_line[39][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51567_ (.CLK(clk),
    .D(net287),
    .Q(\delay_line[39][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51568_ (.CLK(clk),
    .D(net286),
    .Q(\delay_line[39][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51569_ (.CLK(clk),
    .D(\delay_line[38][10] ),
    .Q(\delay_line[39][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51570_ (.CLK(clk),
    .D(\delay_line[38][11] ),
    .Q(\delay_line[39][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51571_ (.CLK(clk),
    .D(net285),
    .Q(\delay_line[39][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51572_ (.CLK(clk),
    .D(\delay_line[38][13] ),
    .Q(\delay_line[39][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51573_ (.CLK(clk),
    .D(\delay_line[38][14] ),
    .Q(\delay_line[39][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51574_ (.CLK(clk),
    .D(net284),
    .Q(\delay_line[39][15] ));
 sky130_fd_sc_hd__dfxtp_1 _51575_ (.CLK(clk),
    .D(\delay_line[39][0] ),
    .Q(\delay_line[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _51576_ (.CLK(clk),
    .D(\delay_line[39][1] ),
    .Q(\delay_line[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _51577_ (.CLK(clk),
    .D(\delay_line[39][2] ),
    .Q(\delay_line[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _51578_ (.CLK(clk),
    .D(\delay_line[39][3] ),
    .Q(\delay_line[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _51579_ (.CLK(clk),
    .D(\delay_line[39][4] ),
    .Q(\delay_line[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 _51580_ (.CLK(clk),
    .D(\delay_line[39][5] ),
    .Q(\delay_line[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 _51581_ (.CLK(clk),
    .D(net283),
    .Q(\delay_line[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 _51582_ (.CLK(clk),
    .D(\delay_line[39][7] ),
    .Q(\delay_line[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 _51583_ (.CLK(clk),
    .D(net281),
    .Q(\delay_line[40][8] ));
 sky130_fd_sc_hd__dfxtp_1 _51584_ (.CLK(clk),
    .D(\delay_line[39][9] ),
    .Q(\delay_line[40][9] ));
 sky130_fd_sc_hd__dfxtp_1 _51585_ (.CLK(clk),
    .D(\delay_line[39][10] ),
    .Q(\delay_line[40][10] ));
 sky130_fd_sc_hd__dfxtp_1 _51586_ (.CLK(clk),
    .D(\delay_line[39][11] ),
    .Q(\delay_line[40][11] ));
 sky130_fd_sc_hd__dfxtp_1 _51587_ (.CLK(clk),
    .D(\delay_line[39][12] ),
    .Q(\delay_line[40][12] ));
 sky130_fd_sc_hd__dfxtp_1 _51588_ (.CLK(clk),
    .D(\delay_line[39][13] ),
    .Q(\delay_line[40][13] ));
 sky130_fd_sc_hd__dfxtp_1 _51589_ (.CLK(clk),
    .D(\delay_line[39][14] ),
    .Q(\delay_line[40][14] ));
 sky130_fd_sc_hd__dfxtp_1 _51590_ (.CLK(clk),
    .D(\delay_line[39][15] ),
    .Q(\delay_line[40][15] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12040 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(data_in[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(data_in[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(data_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(data_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(data_in[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(data_in[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(data_in[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(data_in[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(data_in[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(data_in[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(data_in[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(data_in[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(data_in[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(data_in[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(data_in[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(data_out[0]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(data_out[10]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(data_out[11]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(data_out[12]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(data_out[13]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(data_out[14]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(data_out[15]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(data_out[16]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(data_out[17]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(data_out[18]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(data_out[19]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(data_out[1]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(data_out[20]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(data_out[21]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(data_out[22]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(data_out[23]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(data_out[24]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(data_out[25]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(data_out[26]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(data_out[27]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(data_out[28]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(data_out[29]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(data_out[2]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(data_out[30]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(data_out[31]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(data_out[32]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(data_out[33]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(data_out[34]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(data_out[35]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(data_out[36]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(data_out[37]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(data_out[38]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(data_out[39]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(data_out[3]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(data_out[40]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(data_out[4]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(data_out[5]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(data_out[6]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(data_out[7]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(data_out[8]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(data_out[9]));
 sky130_fd_sc_hd__buf_4 wire58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_2 wire59 (.A(_17754_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 wire60 (.A(_19232_),
    .X(net60));
 sky130_fd_sc_hd__buf_1 wire61 (.A(_16000_),
    .X(net61));
 sky130_fd_sc_hd__buf_1 wire62 (.A(_14871_),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 wire63 (.A(_16976_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 wire64 (.A(_16420_),
    .X(net64));
 sky130_fd_sc_hd__buf_4 wire65 (.A(_15719_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 wire66 (.A(_16778_),
    .X(net66));
 sky130_fd_sc_hd__buf_4 wire67 (.A(_15068_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 wire68 (.A(_15066_),
    .X(net68));
 sky130_fd_sc_hd__buf_1 wire69 (.A(_03527_),
    .X(net69));
 sky130_fd_sc_hd__buf_2 wire70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap71 (.A(_16813_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 wire72 (.A(_14499_),
    .X(net72));
 sky130_fd_sc_hd__buf_1 max_cap73 (.A(_13704_),
    .X(net73));
 sky130_fd_sc_hd__buf_4 wire74 (.A(_16341_),
    .X(net74));
 sky130_fd_sc_hd__buf_1 max_cap75 (.A(_00799_),
    .X(net75));
 sky130_fd_sc_hd__buf_4 wire76 (.A(_16751_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 wire77 (.A(_16402_),
    .X(net77));
 sky130_fd_sc_hd__buf_4 wire78 (.A(_15721_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 wire79 (.A(_15643_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 max_cap80 (.A(_12555_),
    .X(net80));
 sky130_fd_sc_hd__buf_4 wire81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 wire82 (.A(_10972_),
    .X(net82));
 sky130_fd_sc_hd__buf_1 wire83 (.A(_05281_),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 wire84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 max_cap85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 wire86 (.A(_16017_),
    .X(net86));
 sky130_fd_sc_hd__buf_4 wire87 (.A(_12294_),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire88 (.A(_14858_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 max_cap89 (.A(_09482_),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 wire90 (.A(_04422_),
    .X(net90));
 sky130_fd_sc_hd__buf_1 max_cap91 (.A(_04437_),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 max_cap92 (.A(_00598_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 max_cap93 (.A(_00348_),
    .X(net93));
 sky130_fd_sc_hd__buf_1 wire94 (.A(_18217_),
    .X(net94));
 sky130_fd_sc_hd__buf_1 max_cap95 (.A(_06046_),
    .X(net95));
 sky130_fd_sc_hd__buf_1 max_cap96 (.A(_19537_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 max_cap97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__buf_1 wire98 (.A(_18209_),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 max_cap99 (.A(_10130_),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 max_cap100 (.A(_07726_),
    .X(net100));
 sky130_fd_sc_hd__buf_1 max_cap101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__buf_1 wire102 (.A(_00817_),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 max_cap103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_1 wire104 (.A(_20860_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 max_cap105 (.A(_19484_),
    .X(net105));
 sky130_fd_sc_hd__buf_1 wire106 (.A(_07924_),
    .X(net106));
 sky130_fd_sc_hd__buf_1 max_cap107 (.A(_00992_),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 wire108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 max_cap109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 wire110 (.A(_24724_),
    .X(net110));
 sky130_fd_sc_hd__buf_1 wire111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 wire112 (.A(_22913_),
    .X(net112));
 sky130_fd_sc_hd__buf_1 max_cap113 (.A(_21651_),
    .X(net113));
 sky130_fd_sc_hd__buf_2 wire114 (.A(_19380_),
    .X(net114));
 sky130_fd_sc_hd__buf_1 max_cap115 (.A(_24721_),
    .X(net115));
 sky130_fd_sc_hd__buf_1 max_cap116 (.A(_23516_),
    .X(net116));
 sky130_fd_sc_hd__buf_2 max_cap117 (.A(_22981_),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 wire118 (.A(_18691_),
    .X(net118));
 sky130_fd_sc_hd__buf_2 wire119 (.A(_18536_),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 max_cap120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 max_cap121 (.A(_18530_),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 max_cap122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 wire123 (.A(_17854_),
    .X(net123));
 sky130_fd_sc_hd__buf_1 max_cap124 (.A(_16581_),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 max_cap125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 wire126 (.A(_12675_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 max_cap127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 wire128 (.A(_07056_),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 wire129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 max_cap130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 wire131 (.A(_06677_),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 wire132 (.A(_04072_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 max_cap133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 wire134 (.A(_02690_),
    .X(net134));
 sky130_fd_sc_hd__buf_1 max_cap135 (.A(_00988_),
    .X(net135));
 sky130_fd_sc_hd__buf_1 max_cap136 (.A(_00285_),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 wire137 (.A(_22911_),
    .X(net137));
 sky130_fd_sc_hd__buf_1 max_cap138 (.A(_18688_),
    .X(net138));
 sky130_fd_sc_hd__buf_2 max_cap139 (.A(_17807_),
    .X(net139));
 sky130_fd_sc_hd__buf_1 max_cap140 (.A(_02622_),
    .X(net140));
 sky130_fd_sc_hd__buf_2 wire141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 max_cap142 (.A(_19379_),
    .X(net142));
 sky130_fd_sc_hd__buf_1 wire143 (.A(_17132_),
    .X(net143));
 sky130_fd_sc_hd__buf_1 max_cap144 (.A(_15589_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 max_cap145 (.A(_13327_),
    .X(net145));
 sky130_fd_sc_hd__buf_1 wire146 (.A(_10318_),
    .X(net146));
 sky130_fd_sc_hd__buf_1 wire147 (.A(_19941_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 wire148 (.A(_07283_),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 wire149 (.A(_15587_),
    .X(net149));
 sky130_fd_sc_hd__buf_1 max_cap150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_1 wire151 (.A(_13729_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 max_cap152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 wire153 (.A(_11203_),
    .X(net153));
 sky130_fd_sc_hd__buf_1 max_cap154 (.A(_10094_),
    .X(net154));
 sky130_fd_sc_hd__buf_1 wire155 (.A(_09598_),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 max_cap156 (.A(_06073_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 max_cap157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 wire158 (.A(_15962_),
    .X(net158));
 sky130_fd_sc_hd__buf_1 max_cap159 (.A(_15935_),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 wire160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 max_cap161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 wire162 (.A(_15882_),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 max_cap163 (.A(_12772_),
    .X(net163));
 sky130_fd_sc_hd__buf_1 max_cap164 (.A(_12524_),
    .X(net164));
 sky130_fd_sc_hd__buf_1 max_cap165 (.A(_11143_),
    .X(net165));
 sky130_fd_sc_hd__buf_1 max_cap166 (.A(_08989_),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 max_cap167 (.A(_07007_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 max_cap168 (.A(_06522_),
    .X(net168));
 sky130_fd_sc_hd__buf_1 max_cap169 (.A(_05221_),
    .X(net169));
 sky130_fd_sc_hd__buf_1 max_cap170 (.A(_21788_),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 max_cap171 (.A(_21213_),
    .X(net171));
 sky130_fd_sc_hd__buf_1 max_cap172 (.A(_19821_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 max_cap173 (.A(_16579_),
    .X(net173));
 sky130_fd_sc_hd__buf_1 wire174 (.A(_15872_),
    .X(net174));
 sky130_fd_sc_hd__buf_1 max_cap175 (.A(_13529_),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 max_cap176 (.A(_12521_),
    .X(net176));
 sky130_fd_sc_hd__buf_1 max_cap177 (.A(_11483_),
    .X(net177));
 sky130_fd_sc_hd__buf_1 wire178 (.A(_10563_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 max_cap179 (.A(_08424_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 max_cap180 (.A(_01753_),
    .X(net180));
 sky130_fd_sc_hd__buf_1 max_cap181 (.A(_19818_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 max_cap182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 wire183 (.A(_18427_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 max_cap184 (.A(_24699_),
    .X(net184));
 sky130_fd_sc_hd__buf_1 max_cap185 (.A(_23304_),
    .X(net185));
 sky130_fd_sc_hd__buf_1 max_cap186 (.A(_13158_),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 max_cap187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_1 wire188 (.A(_12518_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 max_cap189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 wire190 (.A(_11746_),
    .X(net190));
 sky130_fd_sc_hd__buf_1 max_cap191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_1 wire192 (.A(_11360_),
    .X(net192));
 sky130_fd_sc_hd__buf_1 max_cap193 (.A(_10456_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 max_cap194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 wire195 (.A(_10430_),
    .X(net195));
 sky130_fd_sc_hd__buf_1 max_cap196 (.A(_10309_),
    .X(net196));
 sky130_fd_sc_hd__buf_1 wire197 (.A(_08996_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 max_cap198 (.A(_08465_),
    .X(net198));
 sky130_fd_sc_hd__buf_1 max_cap199 (.A(_08058_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 max_cap200 (.A(_07392_),
    .X(net200));
 sky130_fd_sc_hd__buf_1 max_cap201 (.A(_05325_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 max_cap202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 max_cap203 (.A(_04392_),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 max_cap204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 max_cap205 (.A(_01421_),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 max_cap206 (.A(_01043_),
    .X(net206));
 sky130_fd_sc_hd__buf_1 max_cap207 (.A(_21854_),
    .X(net207));
 sky130_fd_sc_hd__buf_1 max_cap208 (.A(_20950_),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 max_cap209 (.A(_19291_),
    .X(net209));
 sky130_fd_sc_hd__buf_1 max_cap210 (.A(_18735_),
    .X(net210));
 sky130_fd_sc_hd__buf_1 max_cap211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_1 wire212 (.A(_18113_),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 wire213 (.A(_24974_),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 wire214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 wire215 (.A(_17256_),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 max_cap216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 wire217 (.A(_12593_),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 max_cap218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_1 wire219 (.A(_12332_),
    .X(net219));
 sky130_fd_sc_hd__buf_1 max_cap220 (.A(_12194_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 wire221 (.A(_11424_),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 max_cap222 (.A(_11066_),
    .X(net222));
 sky130_fd_sc_hd__buf_1 wire223 (.A(_10799_),
    .X(net223));
 sky130_fd_sc_hd__buf_1 max_cap224 (.A(_08870_),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 max_cap225 (.A(_06791_),
    .X(net225));
 sky130_fd_sc_hd__buf_1 max_cap226 (.A(_06692_),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 max_cap227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 max_cap228 (.A(_04523_),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 max_cap229 (.A(_03937_),
    .X(net229));
 sky130_fd_sc_hd__buf_1 max_cap230 (.A(_02178_),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 max_cap231 (.A(_01801_),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 max_cap232 (.A(_01177_),
    .X(net232));
 sky130_fd_sc_hd__buf_1 max_cap233 (.A(_24466_),
    .X(net233));
 sky130_fd_sc_hd__buf_1 max_cap234 (.A(_23586_),
    .X(net234));
 sky130_fd_sc_hd__buf_1 max_cap235 (.A(_21304_),
    .X(net235));
 sky130_fd_sc_hd__buf_1 max_cap236 (.A(_20832_),
    .X(net236));
 sky130_fd_sc_hd__buf_1 max_cap237 (.A(_19075_),
    .X(net237));
 sky130_fd_sc_hd__buf_1 wire238 (.A(_17917_),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 max_cap239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_1 wire240 (.A(_09536_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 max_cap241 (.A(_05656_),
    .X(net241));
 sky130_fd_sc_hd__buf_4 wire242 (.A(_24424_),
    .X(net242));
 sky130_fd_sc_hd__buf_1 wire243 (.A(_13882_),
    .X(net243));
 sky130_fd_sc_hd__buf_1 wire244 (.A(_12594_),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 wire245 (.A(_12017_),
    .X(net245));
 sky130_fd_sc_hd__buf_1 max_cap246 (.A(_11978_),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 max_cap247 (.A(_11417_),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 max_cap248 (.A(_10320_),
    .X(net248));
 sky130_fd_sc_hd__buf_1 wire249 (.A(_08326_),
    .X(net249));
 sky130_fd_sc_hd__buf_1 wire250 (.A(_07993_),
    .X(net250));
 sky130_fd_sc_hd__buf_1 wire251 (.A(_06435_),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 max_cap252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__buf_1 wire253 (.A(_04391_),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 max_cap254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 wire255 (.A(_02685_),
    .X(net255));
 sky130_fd_sc_hd__buf_1 max_cap256 (.A(_01657_),
    .X(net256));
 sky130_fd_sc_hd__buf_1 wire257 (.A(_01651_),
    .X(net257));
 sky130_fd_sc_hd__buf_1 max_cap258 (.A(_00753_),
    .X(net258));
 sky130_fd_sc_hd__buf_1 wire259 (.A(_23640_),
    .X(net259));
 sky130_fd_sc_hd__buf_1 max_cap260 (.A(_20541_),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 wire261 (.A(_19082_),
    .X(net261));
 sky130_fd_sc_hd__buf_1 wire262 (.A(_11448_),
    .X(net262));
 sky130_fd_sc_hd__buf_1 max_cap263 (.A(_11239_),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 max_cap264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 wire265 (.A(_10774_),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 max_cap266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 wire267 (.A(_07000_),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 max_cap268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 wire269 (.A(_05384_),
    .X(net269));
 sky130_fd_sc_hd__buf_1 max_cap270 (.A(_04758_),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 max_cap271 (.A(_01498_),
    .X(net271));
 sky130_fd_sc_hd__buf_1 max_cap272 (.A(_23468_),
    .X(net272));
 sky130_fd_sc_hd__buf_1 max_cap273 (.A(_21919_),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 wire274 (.A(_19285_),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 max_cap275 (.A(_19068_),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 max_cap276 (.A(_11562_),
    .X(net276));
 sky130_fd_sc_hd__buf_1 wire277 (.A(_05649_),
    .X(net277));
 sky130_fd_sc_hd__buf_1 max_cap278 (.A(_01296_),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 max_cap279 (.A(_25069_),
    .X(net279));
 sky130_fd_sc_hd__buf_1 wire280 (.A(_03216_),
    .X(net280));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout281 (.A(\delay_line[39][8] ),
    .X(net281));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout282 (.A(\delay_line[39][7] ),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_2 fanout283 (.A(\delay_line[39][6] ),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 fanout284 (.A(\delay_line[38][15] ),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 fanout285 (.A(\delay_line[38][12] ),
    .X(net285));
 sky130_fd_sc_hd__buf_1 fanout286 (.A(\delay_line[38][9] ),
    .X(net286));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout287 (.A(\delay_line[38][8] ),
    .X(net287));
 sky130_fd_sc_hd__buf_1 fanout288 (.A(\delay_line[38][4] ),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 fanout289 (.A(\delay_line[38][3] ),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 fanout290 (.A(\delay_line[38][2] ),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 fanout291 (.A(\delay_line[37][15] ),
    .X(net291));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout292 (.A(\delay_line[37][7] ),
    .X(net292));
 sky130_fd_sc_hd__buf_2 fanout293 (.A(\delay_line[37][1] ),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 fanout294 (.A(\delay_line[36][15] ),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 fanout295 (.A(\delay_line[36][14] ),
    .X(net295));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout296 (.A(\delay_line[36][9] ),
    .X(net296));
 sky130_fd_sc_hd__buf_1 fanout297 (.A(\delay_line[36][7] ),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 fanout298 (.A(\delay_line[36][1] ),
    .X(net298));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout299 (.A(\delay_line[35][14] ),
    .X(net299));
 sky130_fd_sc_hd__buf_1 fanout300 (.A(\delay_line[35][13] ),
    .X(net300));
 sky130_fd_sc_hd__buf_1 fanout301 (.A(\delay_line[35][12] ),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 fanout302 (.A(\delay_line[35][0] ),
    .X(net302));
 sky130_fd_sc_hd__buf_1 fanout303 (.A(\delay_line[34][15] ),
    .X(net303));
 sky130_fd_sc_hd__buf_1 fanout304 (.A(\delay_line[34][14] ),
    .X(net304));
 sky130_fd_sc_hd__buf_1 fanout305 (.A(\delay_line[34][12] ),
    .X(net305));
 sky130_fd_sc_hd__buf_1 fanout306 (.A(\delay_line[34][11] ),
    .X(net306));
 sky130_fd_sc_hd__buf_1 fanout307 (.A(\delay_line[34][2] ),
    .X(net307));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout308 (.A(\delay_line[34][1] ),
    .X(net308));
 sky130_fd_sc_hd__buf_1 fanout309 (.A(\delay_line[33][15] ),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 fanout310 (.A(\delay_line[33][14] ),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 fanout311 (.A(\delay_line[33][13] ),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_2 fanout312 (.A(\delay_line[33][5] ),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 fanout313 (.A(\delay_line[33][3] ),
    .X(net313));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout314 (.A(\delay_line[33][2] ),
    .X(net314));
 sky130_fd_sc_hd__buf_1 fanout315 (.A(\delay_line[33][0] ),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_2 fanout316 (.A(\delay_line[31][11] ),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 fanout317 (.A(\delay_line[31][7] ),
    .X(net317));
 sky130_fd_sc_hd__buf_1 fanout318 (.A(\delay_line[31][4] ),
    .X(net318));
 sky130_fd_sc_hd__buf_1 fanout319 (.A(\delay_line[30][15] ),
    .X(net319));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout320 (.A(\delay_line[30][1] ),
    .X(net320));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout321 (.A(\delay_line[29][9] ),
    .X(net321));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout322 (.A(\delay_line[29][8] ),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 fanout323 (.A(\delay_line[29][1] ),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 fanout324 (.A(\delay_line[28][13] ),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 fanout325 (.A(\delay_line[28][12] ),
    .X(net325));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout326 (.A(\delay_line[28][11] ),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 fanout327 (.A(\delay_line[28][4] ),
    .X(net327));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout328 (.A(\delay_line[28][3] ),
    .X(net328));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout329 (.A(\delay_line[27][15] ),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 fanout330 (.A(\delay_line[27][11] ),
    .X(net330));
 sky130_fd_sc_hd__buf_1 fanout331 (.A(\delay_line[27][9] ),
    .X(net331));
 sky130_fd_sc_hd__buf_1 fanout332 (.A(\delay_line[27][6] ),
    .X(net332));
 sky130_fd_sc_hd__buf_1 fanout333 (.A(\delay_line[27][5] ),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_2 fanout334 (.A(\delay_line[26][14] ),
    .X(net334));
 sky130_fd_sc_hd__buf_1 fanout335 (.A(\delay_line[26][13] ),
    .X(net335));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout336 (.A(\delay_line[26][12] ),
    .X(net336));
 sky130_fd_sc_hd__buf_1 fanout337 (.A(\delay_line[26][9] ),
    .X(net337));
 sky130_fd_sc_hd__buf_1 fanout338 (.A(\delay_line[26][5] ),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 fanout339 (.A(\delay_line[26][2] ),
    .X(net339));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout340 (.A(\delay_line[25][14] ),
    .X(net340));
 sky130_fd_sc_hd__buf_1 fanout341 (.A(\delay_line[24][12] ),
    .X(net341));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout342 (.A(\delay_line[24][8] ),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(\delay_line[24][4] ),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 fanout344 (.A(\delay_line[24][2] ),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 fanout345 (.A(\delay_line[24][1] ),
    .X(net345));
 sky130_fd_sc_hd__buf_2 fanout346 (.A(\delay_line[24][0] ),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 fanout347 (.A(\delay_line[23][12] ),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_2 fanout348 (.A(\delay_line[23][10] ),
    .X(net348));
 sky130_fd_sc_hd__buf_2 fanout349 (.A(\delay_line[23][7] ),
    .X(net349));
 sky130_fd_sc_hd__buf_1 fanout350 (.A(\delay_line[22][15] ),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 fanout351 (.A(\delay_line[22][14] ),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 fanout352 (.A(\delay_line[22][7] ),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 fanout353 (.A(\delay_line[22][5] ),
    .X(net353));
 sky130_fd_sc_hd__buf_2 fanout354 (.A(\delay_line[22][3] ),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 fanout355 (.A(\delay_line[22][2] ),
    .X(net355));
 sky130_fd_sc_hd__buf_2 fanout356 (.A(\delay_line[22][1] ),
    .X(net356));
 sky130_fd_sc_hd__buf_1 fanout357 (.A(\delay_line[21][12] ),
    .X(net357));
 sky130_fd_sc_hd__buf_1 fanout358 (.A(\delay_line[21][10] ),
    .X(net358));
 sky130_fd_sc_hd__buf_1 fanout359 (.A(\delay_line[21][8] ),
    .X(net359));
 sky130_fd_sc_hd__buf_1 fanout360 (.A(\delay_line[21][4] ),
    .X(net360));
 sky130_fd_sc_hd__buf_1 fanout361 (.A(\delay_line[21][2] ),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 fanout362 (.A(\delay_line[20][15] ),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 fanout363 (.A(\delay_line[20][14] ),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 fanout364 (.A(\delay_line[20][13] ),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 fanout365 (.A(\delay_line[20][6] ),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 fanout366 (.A(\delay_line[20][5] ),
    .X(net366));
 sky130_fd_sc_hd__buf_1 fanout367 (.A(\delay_line[20][2] ),
    .X(net367));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout368 (.A(\delay_line[20][1] ),
    .X(net368));
 sky130_fd_sc_hd__buf_1 fanout369 (.A(\delay_line[19][13] ),
    .X(net369));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout370 (.A(\delay_line[19][7] ),
    .X(net370));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout371 (.A(\delay_line[19][4] ),
    .X(net371));
 sky130_fd_sc_hd__buf_1 fanout372 (.A(\delay_line[18][15] ),
    .X(net372));
 sky130_fd_sc_hd__buf_1 fanout373 (.A(\delay_line[18][10] ),
    .X(net373));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout374 (.A(\delay_line[18][2] ),
    .X(net374));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout375 (.A(\delay_line[18][1] ),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_2 fanout376 (.A(\delay_line[17][9] ),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_2 fanout377 (.A(\delay_line[17][8] ),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 fanout378 (.A(\delay_line[17][0] ),
    .X(net378));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout379 (.A(\delay_line[16][15] ),
    .X(net379));
 sky130_fd_sc_hd__buf_1 fanout380 (.A(\delay_line[16][14] ),
    .X(net380));
 sky130_fd_sc_hd__buf_1 fanout381 (.A(\delay_line[16][11] ),
    .X(net381));
 sky130_fd_sc_hd__buf_1 fanout382 (.A(\delay_line[16][10] ),
    .X(net382));
 sky130_fd_sc_hd__buf_1 fanout383 (.A(\delay_line[16][8] ),
    .X(net383));
 sky130_fd_sc_hd__buf_1 fanout384 (.A(\delay_line[16][7] ),
    .X(net384));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout385 (.A(\delay_line[16][6] ),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 fanout386 (.A(\delay_line[15][9] ),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 fanout387 (.A(\delay_line[15][4] ),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_2 fanout388 (.A(\delay_line[14][15] ),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 fanout389 (.A(\delay_line[14][14] ),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 fanout390 (.A(\delay_line[14][8] ),
    .X(net390));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout391 (.A(\delay_line[14][5] ),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_2 fanout392 (.A(\delay_line[14][3] ),
    .X(net392));
 sky130_fd_sc_hd__buf_1 fanout393 (.A(\delay_line[14][1] ),
    .X(net393));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout394 (.A(\delay_line[14][0] ),
    .X(net394));
 sky130_fd_sc_hd__buf_4 fanout395 (.A(\delay_line[13][14] ),
    .X(net395));
 sky130_fd_sc_hd__buf_2 fanout396 (.A(\delay_line[13][8] ),
    .X(net396));
 sky130_fd_sc_hd__buf_2 fanout397 (.A(\delay_line[13][5] ),
    .X(net397));
 sky130_fd_sc_hd__buf_2 fanout398 (.A(\delay_line[13][0] ),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 fanout399 (.A(\delay_line[12][15] ),
    .X(net399));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout400 (.A(\delay_line[12][14] ),
    .X(net400));
 sky130_fd_sc_hd__buf_1 fanout401 (.A(\delay_line[12][13] ),
    .X(net401));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout402 (.A(\delay_line[12][12] ),
    .X(net402));
 sky130_fd_sc_hd__buf_1 fanout403 (.A(\delay_line[12][9] ),
    .X(net403));
 sky130_fd_sc_hd__buf_1 fanout404 (.A(\delay_line[12][8] ),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 fanout405 (.A(\delay_line[12][7] ),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_2 fanout406 (.A(\delay_line[12][5] ),
    .X(net406));
 sky130_fd_sc_hd__buf_2 fanout407 (.A(\delay_line[12][3] ),
    .X(net407));
 sky130_fd_sc_hd__buf_2 fanout408 (.A(\delay_line[11][15] ),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 fanout409 (.A(\delay_line[11][14] ),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_4 fanout410 (.A(\delay_line[11][11] ),
    .X(net410));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout411 (.A(\delay_line[10][13] ),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 fanout412 (.A(\delay_line[10][7] ),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_2 fanout413 (.A(\delay_line[10][4] ),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_2 fanout414 (.A(\delay_line[10][2] ),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_2 fanout415 (.A(\delay_line[10][0] ),
    .X(net415));
 sky130_fd_sc_hd__buf_1 fanout416 (.A(\delay_line[9][13] ),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 fanout417 (.A(\delay_line[9][12] ),
    .X(net417));
 sky130_fd_sc_hd__buf_2 fanout418 (.A(\delay_line[9][11] ),
    .X(net418));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout419 (.A(\delay_line[9][8] ),
    .X(net419));
 sky130_fd_sc_hd__buf_1 fanout420 (.A(\delay_line[9][7] ),
    .X(net420));
 sky130_fd_sc_hd__buf_1 fanout421 (.A(\delay_line[9][6] ),
    .X(net421));
 sky130_fd_sc_hd__buf_1 fanout422 (.A(\delay_line[9][3] ),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_2 fanout423 (.A(\delay_line[8][14] ),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 fanout424 (.A(\delay_line[8][8] ),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_2 fanout425 (.A(\delay_line[7][9] ),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_2 fanout426 (.A(\delay_line[6][13] ),
    .X(net426));
 sky130_fd_sc_hd__buf_1 fanout427 (.A(\delay_line[6][11] ),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 fanout428 (.A(\delay_line[6][6] ),
    .X(net428));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout429 (.A(\delay_line[6][5] ),
    .X(net429));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout430 (.A(\delay_line[5][10] ),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 fanout431 (.A(\delay_line[5][2] ),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_4 fanout432 (.A(\delay_line[4][14] ),
    .X(net432));
 sky130_fd_sc_hd__buf_4 fanout433 (.A(\delay_line[4][12] ),
    .X(net433));
 sky130_fd_sc_hd__buf_1 fanout434 (.A(\delay_line[4][4] ),
    .X(net434));
 sky130_fd_sc_hd__buf_1 fanout435 (.A(\delay_line[3][14] ),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 fanout436 (.A(\delay_line[3][3] ),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_2 fanout437 (.A(\delay_line[3][1] ),
    .X(net437));
 sky130_fd_sc_hd__buf_1 fanout438 (.A(\delay_line[2][15] ),
    .X(net438));
 sky130_fd_sc_hd__buf_1 fanout439 (.A(\delay_line[2][13] ),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_2 fanout440 (.A(\delay_line[2][10] ),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_2 fanout441 (.A(\delay_line[2][9] ),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 fanout442 (.A(\delay_line[2][8] ),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 fanout443 (.A(\delay_line[2][5] ),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_2 fanout444 (.A(\delay_line[2][4] ),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_2 fanout445 (.A(\delay_line[1][15] ),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_2 fanout446 (.A(\delay_line[1][14] ),
    .X(net446));
 sky130_fd_sc_hd__buf_1 fanout447 (.A(\delay_line[1][13] ),
    .X(net447));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout448 (.A(\delay_line[1][11] ),
    .X(net448));
 sky130_fd_sc_hd__buf_1 fanout449 (.A(\delay_line[1][10] ),
    .X(net449));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout450 (.A(\delay_line[1][8] ),
    .X(net450));
 sky130_fd_sc_hd__buf_1 fanout451 (.A(\delay_line[1][4] ),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_2 fanout452 (.A(\delay_line[0][14] ),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 fanout453 (.A(\delay_line[0][13] ),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 fanout454 (.A(\delay_line[0][12] ),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_2 fanout455 (.A(\delay_line[0][8] ),
    .X(net455));
endmodule
