VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO FIR_Lowpass_Filter
  CLASS BLOCK ;
  FOREIGN FIR_Lowpass_Filter ;
  ORIGIN 0.000 0.000 ;
  SIZE 905.110 BY 915.830 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 903.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 899.540 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 899.540 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 899.540 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 899.540 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 899.540 644.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 795.930 899.540 797.530 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 903.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 903.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 899.540 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 899.540 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 899.540 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 899.540 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 899.540 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 792.630 899.540 794.230 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 28.600 905.110 29.200 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 599.800 905.110 600.400 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 656.920 905.110 657.520 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 714.040 905.110 714.640 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 771.160 905.110 771.760 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 828.280 905.110 828.880 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 885.400 905.110 886.000 ;
    END
  END data_in[15]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 85.720 905.110 86.320 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 142.840 905.110 143.440 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 199.960 905.110 200.560 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 257.080 905.110 257.680 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 314.200 905.110 314.800 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 371.320 905.110 371.920 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 428.440 905.110 429.040 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 485.560 905.110 486.160 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.110 542.680 905.110 543.280 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END data_out[31]
  PIN data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END data_out[32]
  PIN data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END data_out[33]
  PIN data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END data_out[34]
  PIN data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 4.000 784.000 ;
    END
  END data_out[35]
  PIN data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END data_out[36]
  PIN data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.920 4.000 827.520 ;
    END
  END data_out[37]
  PIN data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END data_out[38]
  PIN data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END data_out[39]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END data_out[3]
  PIN data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END data_out[40]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END data_out[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 899.300 903.125 ;
      LAYER met1 ;
        RECT 5.520 10.640 899.300 903.280 ;
      LAYER met2 ;
        RECT 558.600 72.345 681.560 72.660 ;
      LAYER met3 ;
        RECT 13.640 72.195 898.080 72.495 ;
      LAYER met4 ;
        RECT 36.880 71.725 174.240 72.345 ;
        RECT 176.640 71.725 177.540 72.345 ;
        RECT 179.940 71.725 327.840 72.345 ;
        RECT 330.240 71.725 331.140 72.345 ;
        RECT 333.540 71.725 481.440 72.345 ;
        RECT 483.840 71.725 484.740 72.345 ;
        RECT 487.140 71.725 635.040 72.345 ;
        RECT 637.440 71.725 638.340 72.345 ;
        RECT 640.740 71.725 788.640 72.345 ;
        RECT 791.040 71.725 791.940 72.345 ;
        RECT 794.340 71.725 814.580 72.345 ;
  END
END FIR_Lowpass_Filter
END LIBRARY

